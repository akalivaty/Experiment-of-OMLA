//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT89), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(KEYINPUT89), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n212), .A2(G43gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT15), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n218), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT14), .B(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n210), .A2(new_n211), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n221), .ZN(new_n224));
  INV_X1    g023(.A(new_n219), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n208), .A2(KEYINPUT89), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT15), .A4(new_n209), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT91), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n223), .A2(new_n228), .A3(KEYINPUT91), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G15gat), .B(G22gat), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT16), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G1gat), .B2(new_n235), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G8gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n228), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(KEYINPUT17), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n239), .B(G8gat), .Z(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n241), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n207), .B1(new_n250), .B2(KEYINPUT93), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n246), .B1(new_n234), .B2(new_n242), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n244), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT18), .A3(new_n244), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n255));
  INV_X1    g054(.A(new_n241), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(new_n240), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n244), .B(KEYINPUT13), .Z(new_n258));
  AOI22_X1  g057(.A1(new_n254), .A2(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT93), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n248), .A2(new_n260), .A3(new_n249), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n251), .A2(new_n253), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n255), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n258), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n263), .A2(new_n250), .A3(new_n253), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n207), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G169gat), .ZN(new_n272));
  INV_X1    g071(.A(G176gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT26), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n274), .B(new_n275), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT64), .B(G190gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n280), .B1(KEYINPUT28), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT28), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(G183gat), .C1(new_n291), .C2(new_n292), .ZN(new_n295));
  INV_X1    g094(.A(G183gat), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT65), .B(KEYINPUT27), .C1(new_n296), .C2(KEYINPUT66), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n290), .A2(new_n293), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n284), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(new_n288), .A3(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n275), .A2(KEYINPUT24), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT24), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n306), .A2(new_n308), .A3(new_n278), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n301), .A2(new_n303), .B1(new_n296), .B2(new_n285), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n306), .A2(new_n308), .A3(new_n278), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G113gat), .ZN(new_n318));
  INV_X1    g117(.A(G113gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G127gat), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G134gat), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n321), .A2(new_n322), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n326), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(KEYINPUT1), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n316), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n331), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n299), .B2(new_n315), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n271), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT32), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G15gat), .B(G43gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT67), .Z(new_n340));
  INV_X1    g139(.A(G71gat), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G99gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(G99gat), .A3(new_n343), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n336), .A2(new_n338), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  OAI211_X1 g149(.A(KEYINPUT32), .B(new_n335), .C1(new_n350), .C2(new_n337), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n334), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n298), .A2(new_n284), .B1(new_n310), .B2(new_n314), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n333), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n353), .B(new_n355), .C1(new_n269), .C2(new_n270), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT34), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(KEYINPUT68), .A3(KEYINPUT34), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n349), .A2(new_n359), .A3(new_n351), .A4(new_n360), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n352), .A2(KEYINPUT69), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(new_n370), .A3(new_n364), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n361), .A3(KEYINPUT69), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT70), .B1(new_n373), .B2(KEYINPUT36), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT36), .ZN(new_n376));
  AOI211_X1 g175(.A(new_n375), .B(new_n376), .C1(new_n371), .C2(new_n372), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n369), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT40), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  XOR2_X1   g179(.A(G155gat), .B(G162gat), .Z(new_n381));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT2), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(G141gat), .ZN(new_n385));
  INV_X1    g184(.A(G141gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(G148gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n383), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n381), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(G148gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n384), .A2(G141gat), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n391), .A2(new_n392), .B1(KEYINPUT2), .B2(new_n382), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT78), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT78), .B(new_n381), .C1(new_n393), .C2(new_n394), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n380), .B(new_n331), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n389), .B1(new_n388), .B2(KEYINPUT77), .ZN(new_n399));
  XNOR2_X1  g198(.A(G155gat), .B(G162gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n393), .B2(KEYINPUT78), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT4), .B1(new_n402), .B2(new_n333), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(KEYINPUT3), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n331), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n402), .A2(new_n333), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n331), .B(new_n397), .C1(new_n399), .C2(new_n401), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n412), .A2(KEYINPUT39), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(G57gat), .B(G85gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n412), .B2(KEYINPUT39), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n379), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n429), .B(KEYINPUT74), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n316), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n430), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n354), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(G211gat), .A2(G218gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(G211gat), .A2(G218gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G197gat), .ZN(new_n438));
  INV_X1    g237(.A(G204gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G197gat), .A2(G204gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT22), .ZN(new_n442));
  NAND2_X1  g241(.A1(G211gat), .A2(G218gat), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n440), .A2(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n437), .B1(new_n444), .B2(KEYINPUT72), .ZN(new_n445));
  NOR2_X1   g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446));
  AND2_X1   g245(.A1(G197gat), .A2(G204gat), .ZN(new_n447));
  OAI22_X1  g246(.A1(new_n446), .A2(new_n447), .B1(new_n435), .B2(KEYINPUT22), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n449));
  XNOR2_X1  g248(.A(G211gat), .B(G218gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n445), .A2(KEYINPUT73), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT73), .B1(new_n445), .B2(new_n451), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n432), .A2(new_n434), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n444), .A2(KEYINPUT72), .A3(new_n437), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n445), .A2(new_n451), .A3(KEYINPUT73), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n433), .B1(new_n354), .B2(KEYINPUT29), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n316), .A2(new_n430), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n428), .B1(new_n455), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT76), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n454), .B1(new_n432), .B2(new_n434), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n461), .A3(new_n463), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(KEYINPUT76), .A3(new_n428), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT30), .B(new_n428), .C1(new_n455), .C2(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT75), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n471), .A2(new_n476), .A3(KEYINPUT30), .A4(new_n428), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n471), .A2(new_n428), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n413), .A2(new_n380), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n331), .B1(new_n396), .B2(new_n397), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n408), .A2(new_n481), .A3(new_n483), .A4(new_n410), .ZN(new_n484));
  INV_X1    g283(.A(new_n414), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n411), .B1(new_n485), .B2(new_n482), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n404), .A2(KEYINPUT5), .A3(new_n410), .A4(new_n408), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n420), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n416), .A2(new_n422), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(KEYINPUT40), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n425), .A2(new_n480), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT37), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n428), .B1(new_n471), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n496), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n467), .A2(new_n472), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n499), .B2(new_n495), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n420), .B1(new_n488), .B2(new_n489), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT85), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n508), .A2(KEYINPUT85), .A3(new_n509), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n490), .A2(new_n507), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT29), .B1(new_n402), .B2(new_n405), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT80), .B1(new_n515), .B2(new_n454), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT80), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT3), .B1(new_n396), .B2(new_n397), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n461), .B(new_n517), .C1(new_n518), .C2(KEYINPUT29), .ZN(new_n519));
  INV_X1    g318(.A(new_n402), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n448), .A2(new_n450), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n444), .A2(new_n437), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n431), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n520), .B(new_n521), .C1(KEYINPUT3), .C2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n407), .B(KEYINPUT79), .C1(new_n402), .C2(new_n524), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n516), .A2(new_n519), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G228gat), .A2(G233gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n461), .B1(new_n518), .B2(KEYINPUT29), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n445), .A2(new_n451), .A3(new_n431), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n405), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G22gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G78gat), .B(G106gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G50gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT81), .B(G22gat), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n537), .B(new_n540), .C1(new_n542), .C2(new_n536), .ZN(new_n543));
  INV_X1    g342(.A(new_n535), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n542), .B(new_n544), .C1(new_n528), .C2(new_n529), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n546), .A3(new_n542), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n544), .B1(new_n528), .B2(new_n529), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT82), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n543), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n494), .A2(new_n514), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(KEYINPUT83), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT83), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(new_n543), .C1(new_n550), .C2(new_n540), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n490), .A2(new_n507), .ZN(new_n556));
  INV_X1    g355(.A(new_n509), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n512), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n553), .B(new_n555), .C1(new_n558), .C2(new_n480), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n378), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n480), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n551), .A2(new_n561), .A3(new_n373), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT35), .ZN(new_n563));
  NOR4_X1   g362(.A1(new_n480), .A2(new_n363), .A3(KEYINPUT35), .A4(new_n365), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n513), .A2(new_n510), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n551), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n268), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT100), .ZN(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT97), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  INV_X1    g376(.A(G92gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT8), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G106gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n345), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n580), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(KEYINPUT98), .A3(new_n580), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n575), .A2(new_n576), .ZN(new_n590));
  OAI211_X1 g389(.A(G85gat), .B(G92gat), .C1(KEYINPUT97), .C2(KEYINPUT7), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n583), .A2(new_n588), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n587), .B(new_n586), .C1(new_n595), .C2(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n241), .B2(KEYINPUT17), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n234), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n256), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n574), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n573), .A3(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  INV_X1    g409(.A(KEYINPUT9), .ZN(new_n611));
  INV_X1    g410(.A(G78gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n341), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G57gat), .B(G64gat), .Z(new_n614));
  XOR2_X1   g413(.A(G71gat), .B(G78gat), .Z(new_n615));
  OAI211_X1 g414(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(KEYINPUT94), .ZN(new_n616));
  OR2_X1    g415(.A1(G57gat), .A2(G64gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(G57gat), .A2(G64gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G78gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(KEYINPUT94), .A3(new_n618), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n616), .A2(new_n622), .A3(KEYINPUT95), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT95), .B1(new_n616), .B2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n610), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n616), .A2(new_n622), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n616), .A2(new_n622), .A3(KEYINPUT95), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n626), .ZN(new_n633));
  INV_X1    g432(.A(new_n610), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G183gat), .B(G211gat), .Z(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT21), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n245), .B1(new_n632), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n636), .A2(new_n637), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n639), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n638), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n609), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n628), .B1(new_n596), .B2(new_n594), .ZN(new_n661));
  INV_X1    g460(.A(new_n597), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n625), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n663), .B2(KEYINPUT10), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n630), .A2(new_n631), .A3(new_n596), .A4(new_n594), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n597), .A2(new_n616), .A3(new_n622), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT99), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n632), .A2(new_n662), .A3(new_n668), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n659), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n667), .A2(new_n658), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n657), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT99), .B1(new_n667), .B2(new_n668), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n660), .B(KEYINPUT10), .C1(new_n665), .C2(new_n666), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n658), .ZN(new_n679));
  INV_X1    g478(.A(new_n674), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n656), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n569), .B1(new_n653), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n675), .A2(new_n681), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n652), .A4(new_n609), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n568), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n558), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n236), .ZN(G1324gat));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  INV_X1    g489(.A(new_n480), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n693), .B2(G8gat), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n698));
  MUX2_X1   g497(.A(KEYINPUT102), .B(new_n698), .S(new_n696), .Z(new_n699));
  AOI22_X1  g498(.A1(new_n694), .A2(new_n697), .B1(new_n692), .B2(new_n699), .ZN(G1325gat));
  OAI21_X1  g499(.A(G15gat), .B1(new_n686), .B2(new_n378), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n367), .A2(G15gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n686), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n553), .A2(new_n555), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n686), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n563), .A2(new_n708), .A3(new_n566), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(new_n563), .B2(new_n566), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n560), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n609), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n560), .A2(new_n567), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(KEYINPUT44), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n682), .A2(new_n652), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n267), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT103), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n687), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n568), .A2(new_n712), .A3(new_n719), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n218), .A3(new_n558), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(G1328gat));
  OAI21_X1  g527(.A(G36gat), .B1(new_n723), .B2(new_n691), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n725), .A2(new_n221), .A3(new_n480), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1329gat));
  INV_X1    g531(.A(new_n378), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n213), .A2(new_n214), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n722), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n725), .B2(new_n366), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1330gat));
  OAI21_X1  g538(.A(G50gat), .B1(new_n723), .B2(new_n551), .ZN(new_n740));
  INV_X1    g539(.A(new_n704), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n212), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(KEYINPUT48), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n212), .B1(new_n722), .B2(new_n741), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n744), .B2(KEYINPUT105), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n747), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g547(.A1(new_n267), .A2(new_n684), .A3(new_n653), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n711), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n558), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n750), .A2(new_n691), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NOR3_X1   g557(.A1(new_n750), .A2(G71gat), .A3(new_n367), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n751), .A2(new_n733), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(G71gat), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n750), .A2(new_n704), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n612), .ZN(G1335gat));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n267), .A2(new_n652), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n712), .A4(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n768), .A2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(KEYINPUT110), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n567), .A2(KEYINPUT104), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n563), .A2(new_n708), .A3(new_n566), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n609), .B1(new_n779), .B2(new_n560), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n780), .B2(new_n767), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(new_n577), .A3(new_n558), .A4(new_n682), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n682), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT107), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n717), .B(new_n786), .C1(new_n780), .C2(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT108), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n715), .A2(new_n790), .A3(new_n717), .A4(new_n786), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n789), .A2(new_n792), .A3(new_n687), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n784), .B1(new_n577), .B2(new_n793), .ZN(G1336gat));
  NOR2_X1   g593(.A1(new_n691), .A2(G92gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n682), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n797));
  INV_X1    g596(.A(new_n787), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n480), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(G92gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n788), .A2(new_n480), .A3(new_n791), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n782), .B1(new_n770), .B2(new_n771), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n691), .A2(new_n684), .A3(G92gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT111), .B1(new_n807), .B2(KEYINPUT52), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n802), .A2(G92gat), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n801), .B1(new_n808), .B2(new_n812), .ZN(G1337gat));
  NAND4_X1  g612(.A1(new_n783), .A2(new_n345), .A3(new_n366), .A4(new_n682), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n789), .A2(new_n792), .A3(new_n378), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n345), .B2(new_n815), .ZN(G1338gat));
  INV_X1    g615(.A(new_n551), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n584), .A3(new_n682), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n789), .A2(new_n792), .A3(new_n704), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n584), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n781), .B1(new_n772), .B2(new_n775), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT113), .B1(new_n824), .B2(new_n818), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n798), .A2(new_n817), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT53), .B1(new_n826), .B2(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n824), .A2(KEYINPUT113), .A3(new_n818), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(G1339gat));
  OR3_X1    g629(.A1(new_n267), .A2(new_n653), .A3(new_n682), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n671), .B1(new_n664), .B2(new_n669), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT54), .B1(new_n833), .B2(new_n659), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n678), .A2(new_n658), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n678), .A2(new_n837), .A3(new_n658), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n657), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n832), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n712), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n656), .B1(new_n673), .B2(new_n837), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n670), .A2(new_n659), .A3(new_n672), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n679), .A2(KEYINPUT54), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n844), .A3(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n681), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n252), .A2(new_n244), .B1(new_n257), .B2(new_n258), .ZN(new_n847));
  INV_X1    g646(.A(new_n205), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n262), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n841), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n267), .A2(new_n840), .A3(new_n681), .A4(new_n845), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n682), .A2(new_n262), .A3(new_n849), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n682), .A2(new_n262), .A3(KEYINPUT114), .A4(new_n849), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n851), .B1(new_n857), .B2(new_n609), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n831), .B1(new_n858), .B2(new_n652), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n558), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n551), .A2(new_n691), .A3(new_n373), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n267), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n859), .A2(new_n704), .A3(new_n366), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n687), .A2(new_n480), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT115), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n268), .A2(new_n319), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  INV_X1    g668(.A(new_n867), .ZN(new_n870));
  OAI21_X1  g669(.A(G120gat), .B1(new_n870), .B2(new_n684), .ZN(new_n871));
  INV_X1    g670(.A(new_n862), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n682), .A2(new_n317), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT116), .Z(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(G1341gat));
  INV_X1    g674(.A(new_n652), .ZN(new_n876));
  OAI21_X1  g675(.A(G127gat), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n325), .A3(new_n652), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1342gat));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n323), .A3(new_n712), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(KEYINPUT117), .B2(KEYINPUT56), .ZN(new_n881));
  NAND2_X1  g680(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n881), .B(new_n882), .Z(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n870), .B2(new_n609), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1343gat));
  AND2_X1   g684(.A1(new_n378), .A2(new_n865), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n836), .B2(new_n839), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n842), .A2(new_n844), .A3(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n832), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n845), .A2(new_n681), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n267), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n712), .B1(new_n893), .B2(new_n853), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n876), .B1(new_n894), .B2(new_n851), .ZN(new_n895));
  AOI211_X1 g694(.A(new_n887), .B(new_n704), .C1(new_n895), .C2(new_n831), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT57), .B1(new_n859), .B2(new_n817), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n886), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n898), .B2(new_n268), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n733), .A2(new_n551), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n480), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n860), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n267), .A2(new_n386), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT58), .ZN(G1344gat));
  OR2_X1    g705(.A1(new_n898), .A2(new_n684), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(KEYINPUT59), .A3(new_n384), .ZN(new_n909));
  XOR2_X1   g708(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n910));
  NAND2_X1  g709(.A1(new_n859), .A2(new_n817), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT57), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n741), .A2(new_n887), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n685), .A2(new_n683), .A3(new_n268), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n895), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n912), .A2(new_n918), .A3(new_n682), .A4(new_n886), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n910), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n682), .A2(new_n384), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n909), .A2(new_n920), .B1(new_n903), .B2(new_n921), .ZN(G1345gat));
  NAND3_X1  g721(.A1(new_n860), .A2(new_n902), .A3(new_n652), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT121), .ZN(new_n924));
  INV_X1    g723(.A(G155gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n923), .B2(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n652), .A2(G155gat), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n924), .A2(new_n926), .B1(new_n898), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(G1346gat));
  NOR2_X1   g728(.A1(new_n609), .A2(G162gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n860), .A2(new_n902), .A3(new_n930), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT122), .Z(new_n932));
  OAI21_X1  g731(.A(G162gat), .B1(new_n898), .B2(new_n609), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT123), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n691), .A2(new_n558), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n864), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n272), .A3(new_n268), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n859), .A2(new_n687), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n551), .A2(new_n480), .A3(new_n373), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n267), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n938), .A2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n937), .B2(new_n684), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(new_n273), .A3(new_n682), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n937), .B2(new_n876), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n282), .A3(new_n652), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n937), .B2(new_n609), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n942), .A2(new_n281), .A3(new_n712), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n691), .A3(new_n901), .ZN(new_n956));
  AOI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n267), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n887), .B1(new_n859), .B2(new_n817), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n378), .A2(new_n936), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n958), .A2(new_n917), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n268), .A2(new_n438), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  AOI21_X1  g761(.A(G204gat), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n956), .A2(new_n682), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n960), .ZN(new_n967));
  OAI21_X1  g766(.A(G204gat), .B1(new_n967), .B2(new_n684), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1353gat));
  INV_X1    g768(.A(G211gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n956), .A2(new_n970), .A3(new_n652), .ZN(new_n971));
  NOR4_X1   g770(.A1(new_n958), .A2(new_n917), .A3(new_n876), .A4(new_n959), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n959), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n912), .A2(new_n918), .A3(new_n652), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  AND4_X1   g776(.A1(KEYINPUT63), .A2(new_n974), .A3(new_n977), .A4(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n979), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n971), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(KEYINPUT127), .B(new_n971), .C1(new_n978), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(G218gat), .B1(new_n967), .B2(new_n609), .ZN(new_n986));
  INV_X1    g785(.A(G218gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n956), .A2(new_n987), .A3(new_n712), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(G1355gat));
endmodule


