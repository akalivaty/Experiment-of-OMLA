//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n204), .B(new_n205), .ZN(G355));
  INV_X1    g0006(.A(KEYINPUT65), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n207), .B1(new_n208), .B2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G13), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n210), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n214), .B(new_n228), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n223), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n222), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT66), .B(G50), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(new_n230), .A2(G33), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G77), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n229), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT12), .B1(new_n261), .B2(G68), .ZN(new_n262));
  OR3_X1    g0062(.A1(new_n261), .A2(KEYINPUT12), .A3(G68), .ZN(new_n263));
  INV_X1    g0063(.A(new_n261), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n258), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n216), .B1(new_n260), .B2(G20), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n262), .A2(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT11), .B1(new_n256), .B2(new_n258), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(G232), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  OAI211_X1 g0075(.A(G226), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n274), .B(new_n276), .C1(new_n277), .C2(new_n224), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n280), .A3(G274), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT76), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  INV_X1    g0088(.A(new_n229), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(new_n279), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT76), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(new_n285), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n280), .A2(G238), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n287), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT77), .B1(new_n282), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n295), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT77), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n278), .A2(new_n281), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n296), .A2(new_n300), .A3(KEYINPUT13), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT13), .B1(new_n282), .B2(new_n295), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n301), .A2(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n308), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n271), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n303), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n270), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n282), .A2(new_n295), .A3(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n296), .A2(new_n300), .A3(KEYINPUT13), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n265), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT8), .B(G58), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n260), .A2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n323), .A2(new_n327), .B1(new_n325), .B2(new_n261), .ZN(new_n328));
  INV_X1    g0128(.A(new_n258), .ZN(new_n329));
  AND3_X1   g0129(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT79), .B1(G58), .B2(G68), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G159), .ZN(new_n334));
  INV_X1    g0134(.A(new_n254), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n333), .A2(new_n230), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n272), .A2(new_n273), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n342), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n230), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n230), .A3(new_n338), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n336), .B1(new_n347), .B2(G68), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n329), .B1(new_n348), .B2(KEYINPUT16), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n216), .B1(new_n346), .B2(new_n339), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n336), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n328), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G226), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G1698), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n355), .B1(G223), .B2(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G87), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n280), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n280), .A2(new_n293), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n286), .B1(new_n223), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n358), .A2(new_n360), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(G169), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT18), .B1(new_n353), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n347), .A2(G68), .ZN(new_n366));
  INV_X1    g0166(.A(new_n336), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(new_n258), .A3(new_n352), .ZN(new_n369));
  INV_X1    g0169(.A(new_n328), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n364), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n358), .A2(new_n360), .A3(new_n317), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G200), .B2(new_n363), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n353), .A2(KEYINPUT17), .A3(new_n376), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n365), .A2(new_n374), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n326), .A2(G77), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n323), .A2(new_n382), .B1(G77), .B2(new_n261), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n325), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(KEYINPUT72), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(KEYINPUT72), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n384), .B1(new_n388), .B2(new_n251), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n383), .B1(new_n389), .B2(new_n258), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI211_X1 g0191(.A(G232), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n392));
  OAI211_X1 g0192(.A(G238), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n393));
  INV_X1    g0193(.A(G107), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n337), .A2(new_n338), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n281), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n280), .A2(G244), .A3(new_n293), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n286), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT71), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n286), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n305), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(G200), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n390), .A2(new_n407), .A3(KEYINPUT73), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n403), .A2(new_n317), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT73), .B1(new_n390), .B2(new_n407), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OR3_X1    g0212(.A1(new_n322), .A2(new_n381), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(G1698), .B1(new_n337), .B2(new_n338), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G222), .B1(new_n342), .B2(G77), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n395), .A2(G1698), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT67), .B(G223), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n280), .B1(new_n418), .B2(KEYINPUT68), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT68), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n415), .B(new_n420), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n286), .B1(new_n354), .B2(new_n359), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G200), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n419), .B2(new_n421), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G190), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT9), .ZN(new_n429));
  INV_X1    g0229(.A(G150), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n335), .B1(new_n201), .B2(new_n230), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n252), .B2(new_n325), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n329), .ZN(new_n433));
  INV_X1    g0233(.A(G50), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n260), .B2(G20), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n265), .A2(new_n435), .B1(new_n434), .B2(new_n264), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n429), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT9), .B(new_n436), .C1(new_n432), .C2(new_n329), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n426), .A2(new_n428), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT75), .ZN(new_n444));
  INV_X1    g0244(.A(G200), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n441), .B1(new_n445), .B2(new_n427), .ZN(new_n446));
  INV_X1    g0246(.A(new_n428), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT10), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n440), .B1(new_n425), .B2(G200), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT75), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n428), .A4(new_n442), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT70), .B1(new_n427), .B2(G169), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(G179), .B2(new_n425), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n427), .A2(KEYINPUT70), .A3(new_n361), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(new_n433), .C2(new_n437), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n413), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n219), .A2(new_n275), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n225), .A2(G1698), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(new_n272), .C2(new_n273), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT87), .A2(G294), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT87), .A2(G294), .ZN(new_n464));
  OAI21_X1  g0264(.A(G33), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n462), .A2(KEYINPUT88), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT88), .B1(new_n462), .B2(new_n465), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n466), .A2(new_n467), .A3(new_n280), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n284), .A2(G1), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n469), .A2(new_n470), .B1(new_n289), .B2(new_n279), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G264), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT89), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n467), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n462), .A2(KEYINPUT88), .A3(new_n465), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n281), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT89), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n472), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n290), .A2(new_n470), .A3(new_n469), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n361), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n474), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(new_n472), .ZN(new_n484));
  OAI21_X1  g0284(.A(G169), .B1(new_n484), .B2(new_n481), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n395), .A2(new_n230), .A3(G87), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(new_n337), .B2(new_n338), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT81), .B(G116), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n277), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n230), .A2(G107), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n495), .A2(KEYINPUT23), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(KEYINPUT23), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n494), .A2(new_n230), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n491), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n491), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n258), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n210), .A2(G1), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n502), .A2(new_n495), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n260), .A2(G33), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n261), .A2(new_n506), .A3(new_n229), .A4(new_n257), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n502), .A2(new_n495), .ZN(new_n508));
  OAI221_X1 g0308(.A(new_n505), .B1(new_n507), .B2(new_n394), .C1(new_n504), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n483), .A2(new_n485), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n474), .A2(new_n480), .A3(new_n479), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n445), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n477), .A2(new_n317), .A3(new_n480), .A4(new_n472), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n501), .A2(new_n510), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n511), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n488), .A2(G68), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n251), .A2(new_n224), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(KEYINPUT19), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n522), .A2(KEYINPUT82), .A3(new_n230), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT82), .B1(new_n522), .B2(new_n230), .ZN(new_n524));
  NOR3_X1   g0324(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n258), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n507), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G87), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n388), .A2(new_n264), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n470), .A2(new_n219), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n290), .A2(new_n470), .B1(new_n532), .B2(new_n280), .ZN(new_n533));
  INV_X1    g0333(.A(G116), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT81), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT81), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G33), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n217), .A2(new_n275), .ZN(new_n540));
  INV_X1    g0340(.A(G244), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G1698), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n542), .C1(new_n272), .C2(new_n273), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n533), .B(G190), .C1(new_n544), .C2(new_n280), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n280), .B1(new_n539), .B2(new_n543), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n532), .A2(new_n280), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n280), .A2(G274), .A3(new_n470), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(G200), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n531), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n386), .A2(new_n387), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n528), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n527), .A2(new_n554), .A3(new_n530), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n555), .A2(KEYINPUT83), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n533), .B(G179), .C1(new_n544), .C2(new_n280), .ZN(new_n557));
  OAI21_X1  g0357(.A(G169), .B1(new_n546), .B2(new_n549), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n555), .A2(KEYINPUT83), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n552), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n471), .B2(G270), .ZN(new_n562));
  AND2_X1   g0362(.A1(KEYINPUT5), .A2(G41), .ZN(new_n563));
  NOR2_X1   g0363(.A1(KEYINPUT5), .A2(G41), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n470), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n565), .A2(new_n561), .A3(G270), .A4(new_n280), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n480), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT85), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT85), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n395), .A2(new_n571), .A3(G257), .A4(new_n275), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n337), .A2(G303), .A3(new_n338), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n280), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n568), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n281), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n565), .A2(G270), .A3(new_n280), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT84), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n481), .B1(new_n583), .B2(new_n566), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(G190), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(G20), .B1(G33), .B2(G283), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n277), .A2(G97), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n257), .B2(new_n229), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n535), .A2(new_n537), .A3(G20), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(KEYINPUT20), .A3(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n507), .A2(new_n534), .B1(new_n261), .B2(new_n538), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n579), .A2(new_n585), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n568), .A2(new_n578), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(G179), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n583), .A2(new_n566), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n576), .B1(new_n572), .B2(new_n570), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n480), .C1(new_n280), .C2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n305), .B1(new_n594), .B2(new_n596), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n604), .B2(new_n605), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n599), .B(new_n601), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT6), .ZN(new_n610));
  AND2_X1   g0410(.A1(G97), .A2(G107), .ZN(new_n611));
  NOR2_X1   g0411(.A1(G97), .A2(G107), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n394), .A2(KEYINPUT6), .A3(G97), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n394), .B1(new_n346), .B2(new_n339), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT80), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(KEYINPUT80), .B(new_n394), .C1(new_n346), .C2(new_n339), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n258), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n264), .A2(new_n224), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n507), .B2(new_n224), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(G250), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G283), .ZN(new_n626));
  OAI211_X1 g0426(.A(G244), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT4), .B1(new_n414), .B2(G244), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n281), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n565), .A2(G257), .A3(new_n280), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n480), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n631), .A2(new_n317), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(G200), .B1(new_n631), .B2(new_n634), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n621), .B(new_n624), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n617), .A2(new_n618), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n617), .A2(new_n618), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(new_n616), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n623), .B1(new_n640), .B2(new_n258), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n631), .A2(new_n634), .A3(new_n361), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n414), .A2(KEYINPUT4), .A3(G244), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n627), .A2(new_n628), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n625), .A4(new_n626), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n633), .B1(new_n645), .B2(new_n281), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(G169), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n637), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n609), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n459), .A2(new_n518), .A3(new_n560), .A4(new_n649), .ZN(G372));
  NOR2_X1   g0450(.A1(new_n315), .A2(new_n320), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n312), .B1(new_n651), .B2(new_n406), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n652), .A2(new_n379), .A3(new_n380), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n365), .A2(new_n374), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n452), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n456), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n511), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n483), .A2(new_n485), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n516), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n597), .A2(G179), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n604), .ZN(new_n664));
  INV_X1    g0464(.A(new_n593), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT20), .B1(new_n588), .B2(new_n589), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(G169), .B1(new_n667), .B2(new_n595), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT21), .B1(new_n600), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n604), .A2(new_n606), .A3(new_n605), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n662), .A2(new_n671), .A3(KEYINPUT90), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n515), .A2(new_n517), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n545), .A2(new_n550), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n557), .A2(new_n558), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n674), .A2(new_n675), .B1(new_n555), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n648), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n660), .A2(new_n672), .A3(new_n673), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n641), .A2(new_n647), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n560), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n621), .A2(new_n624), .ZN(new_n684));
  INV_X1    g0484(.A(new_n647), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n677), .A2(new_n681), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n555), .A2(new_n676), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n680), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n657), .B1(new_n458), .B2(new_n691), .ZN(G369));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n502), .A2(new_n230), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n662), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT91), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n518), .B1(new_n517), .B2(new_n700), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n693), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n693), .A3(new_n703), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n671), .A2(new_n699), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n662), .A2(new_n699), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n705), .A2(new_n706), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n598), .A2(new_n700), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n659), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n609), .B2(new_n714), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n712), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n212), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n233), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n525), .A2(new_n534), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G1), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n699), .B1(new_n680), .B2(new_n689), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n560), .A2(new_n682), .A3(new_n681), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n685), .A2(new_n684), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT26), .B1(new_n678), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n732), .A3(new_n687), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n516), .B1(new_n513), .B2(new_n514), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n637), .A3(new_n677), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n659), .A2(new_n511), .A3(KEYINPUT94), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT94), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n662), .B2(new_n671), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT95), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n733), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n736), .B(KEYINPUT95), .C1(new_n737), .C2(new_n739), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n699), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n729), .B1(new_n744), .B2(new_n728), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G330), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n546), .A2(new_n549), .A3(new_n361), .ZN(new_n748));
  AND4_X1   g0548(.A1(new_n748), .A2(new_n646), .A3(new_n581), .A4(new_n584), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT93), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n749), .A2(new_n474), .A3(new_n479), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n546), .A2(new_n549), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n646), .A2(G179), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n512), .A2(new_n604), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n474), .A2(new_n479), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n646), .A2(new_n581), .A3(new_n748), .A4(new_n584), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n753), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n760), .B2(new_n699), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n518), .A2(new_n649), .A3(new_n560), .A4(new_n700), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n747), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n746), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n726), .B1(new_n768), .B2(G1), .ZN(G364));
  INV_X1    g0569(.A(new_n717), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n210), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n260), .B1(new_n771), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n721), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n716), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n229), .B1(G20), .B2(new_n305), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n230), .A2(new_n361), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n445), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n230), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n317), .A3(G200), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n434), .B1(new_n785), .B2(new_n394), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n781), .A2(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n361), .A2(new_n445), .A3(G190), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n788), .A2(new_n222), .B1(new_n224), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n780), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n780), .A2(new_n317), .A3(G200), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n395), .B1(new_n794), .B2(new_n202), .C1(new_n216), .C2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n786), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n798));
  NAND2_X1  g0598(.A1(new_n784), .A2(new_n793), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n334), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n798), .A2(new_n799), .A3(new_n334), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(G87), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n797), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n795), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  INV_X1    g0607(.A(new_n794), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(G311), .ZN(new_n809));
  INV_X1    g0609(.A(new_n799), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n395), .B1(new_n810), .B2(G329), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n463), .A2(new_n464), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n803), .A2(G303), .B1(new_n813), .B2(new_n790), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n809), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G322), .A2(new_n787), .B1(new_n782), .B2(G326), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n785), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n779), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n778), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n720), .A2(new_n395), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n284), .B2(new_n233), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n246), .B2(new_n284), .ZN(new_n827));
  NAND3_X1  g0627(.A1(G355), .A2(new_n212), .A3(new_n395), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G116), .C2(new_n212), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n777), .B(new_n819), .C1(new_n823), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n822), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n716), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n776), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n391), .A2(new_n699), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n406), .B(new_n835), .C1(new_n410), .C2(new_n411), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n690), .A2(new_n700), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n406), .A2(new_n700), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(KEYINPUT99), .C1(new_n727), .C2(new_n842), .ZN(new_n843));
  OR3_X1    g0643(.A1(new_n727), .A2(KEYINPUT99), .A3(new_n842), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n766), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n845), .A2(new_n766), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n847), .A2(new_n777), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n778), .A2(new_n820), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n774), .B1(G77), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n806), .A2(KEYINPUT97), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n806), .A2(KEYINPUT97), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(G283), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n785), .A2(new_n218), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n802), .A2(new_n394), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n859), .B(new_n860), .C1(G303), .C2(new_n782), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n395), .B1(new_n810), .B2(G311), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n493), .B2(new_n794), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n787), .A2(G294), .B1(G97), .B2(new_n790), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n858), .A2(new_n861), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n806), .A2(G150), .B1(new_n808), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  INV_X1    g0668(.A(G143), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n783), .B2(new_n868), .C1(new_n869), .C2(new_n788), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT34), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n395), .B1(new_n799), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G50), .B2(new_n803), .ZN(new_n875));
  INV_X1    g0675(.A(new_n785), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(G68), .B1(new_n790), .B2(G58), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n872), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n870), .A2(new_n871), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n866), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n853), .B1(new_n880), .B2(new_n778), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n842), .B2(new_n821), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n850), .A2(new_n882), .ZN(G384));
  OR2_X1    g0683(.A1(new_n615), .A2(KEYINPUT35), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n615), .A2(KEYINPUT35), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(G116), .A3(new_n231), .A4(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  NOR4_X1   g0687(.A1(new_n330), .A2(new_n331), .A3(new_n232), .A4(new_n202), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(KEYINPUT101), .B1(new_n434), .B2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n260), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n371), .A2(new_n372), .ZN(new_n894));
  INV_X1    g0694(.A(new_n697), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n371), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n894), .A2(new_n896), .A3(new_n897), .A4(new_n377), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n366), .A2(new_n367), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n350), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n328), .B1(new_n901), .B2(new_n349), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT102), .B1(new_n902), .B2(new_n697), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n368), .A2(new_n258), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n348), .A2(KEYINPUT16), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n370), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n895), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n372), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n903), .A2(new_n908), .A3(new_n377), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n899), .B1(KEYINPUT37), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n381), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n893), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n898), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n760), .A2(new_n699), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT31), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n764), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n313), .A2(G169), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT14), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n310), .C1(new_n301), .C2(new_n304), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n271), .B(new_n699), .C1(new_n927), .C2(new_n651), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n271), .A2(new_n699), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n312), .A2(new_n321), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n924), .A2(new_n842), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n377), .B1(new_n353), .B2(new_n364), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n353), .A2(new_n697), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n898), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n381), .A2(new_n937), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n916), .A2(new_n898), .B1(new_n381), .B2(new_n912), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(KEYINPUT38), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n924), .A2(KEYINPUT40), .A3(new_n842), .A4(new_n931), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n459), .A2(new_n924), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n931), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n406), .A2(new_n699), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n840), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n953), .A2(new_n919), .B1(new_n654), .B2(new_n697), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n939), .A2(new_n940), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n893), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n918), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT39), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n312), .A2(new_n699), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT39), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n656), .B1(new_n745), .B2(new_n459), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n949), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n260), .B2(new_n771), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n949), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n892), .B1(new_n967), .B2(new_n968), .ZN(G367));
  INV_X1    g0769(.A(new_n718), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n731), .B(new_n637), .C1(new_n641), .C2(new_n700), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n682), .A2(new_n699), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n970), .A2(KEYINPUT104), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n531), .A2(new_n699), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT103), .Z(new_n977));
  MUX2_X1   g0777(.A(new_n687), .B(new_n678), .S(new_n977), .Z(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT104), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n718), .B2(new_n973), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n975), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n980), .B1(new_n975), .B2(new_n982), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n978), .A2(new_n979), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n707), .A2(new_n708), .A3(new_n973), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n731), .B1(new_n971), .B2(new_n662), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n987), .A2(KEYINPUT42), .B1(new_n700), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n985), .B(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n721), .B(KEYINPUT41), .Z(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT44), .B1(new_n712), .B2(new_n974), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n995), .B(new_n973), .C1(new_n709), .C2(new_n711), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n709), .A2(new_n711), .A3(new_n973), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1000), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n970), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n705), .B(new_n706), .C1(new_n671), .C2(new_n699), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n709), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n717), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n709), .A2(new_n770), .A3(new_n1004), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1008), .A2(new_n767), .A3(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1001), .B(new_n1002), .C1(new_n994), .C2(new_n996), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n718), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT106), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1003), .B(new_n1010), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n993), .B1(new_n1014), .B2(new_n768), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n992), .B1(new_n1015), .B2(new_n773), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n978), .A2(new_n822), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n857), .A2(G159), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n783), .A2(new_n869), .B1(new_n802), .B2(new_n222), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G150), .B2(new_n787), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n395), .B1(new_n799), .B2(new_n868), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n808), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n785), .A2(new_n202), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G68), .B2(new_n790), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n803), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n224), .B2(new_n785), .C1(new_n394), .C2(new_n791), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT108), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT107), .B(G311), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G303), .A2(new_n787), .B1(new_n782), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1027), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n342), .B1(new_n794), .B2(new_n817), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G317), .B2(new_n810), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n802), .A2(new_n493), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1035), .B1(KEYINPUT46), .B2(new_n1036), .C1(new_n856), .C2(new_n812), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1025), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n778), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n823), .B1(new_n212), .B2(new_n388), .C1(new_n825), .C2(new_n241), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1017), .A2(new_n774), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1016), .A2(new_n1042), .ZN(G387));
  INV_X1    g0843(.A(new_n1008), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n768), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n721), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(KEYINPUT111), .B1(new_n767), .B2(new_n1008), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT111), .B2(new_n1046), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n238), .A2(new_n284), .A3(new_n395), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n324), .B2(G50), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n284), .C1(new_n216), .C2(new_n202), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n324), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n342), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n723), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n720), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n823), .B1(new_n394), .B2(new_n212), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n774), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n794), .A2(new_n216), .B1(new_n799), .B2(new_n430), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n342), .B(new_n1058), .C1(new_n325), .C2(new_n806), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n787), .A2(G50), .B1(new_n876), .B2(G97), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n802), .A2(new_n202), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G159), .B2(new_n782), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n553), .A2(new_n790), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n787), .A2(G317), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n782), .A2(G322), .B1(new_n808), .B2(G303), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n856), .C2(new_n1029), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n803), .A2(new_n813), .B1(new_n790), .B2(G283), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT109), .Z(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n395), .B1(new_n810), .B2(G326), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n493), .C2(new_n785), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1064), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1057), .B1(new_n1078), .B2(new_n778), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n707), .B2(new_n831), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT110), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1044), .B2(new_n773), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1048), .A2(new_n1082), .ZN(G393));
  NAND2_X1  g0883(.A1(new_n1003), .A2(new_n1012), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n1045), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n1014), .A3(new_n721), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1003), .A2(new_n1012), .A3(new_n773), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n823), .B1(new_n224), .B2(new_n212), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n249), .B2(new_n824), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n777), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT112), .Z(new_n1091));
  AOI22_X1  g0891(.A1(G150), .A2(new_n782), .B1(new_n787), .B2(G159), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  NOR2_X1   g0893(.A1(new_n791), .A2(new_n202), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n395), .B1(new_n794), .B2(new_n324), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n859), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n802), .A2(new_n216), .B1(new_n799), .B2(new_n869), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT113), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n857), .A2(G50), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1093), .A2(new_n1096), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G311), .A2(new_n787), .B1(new_n782), .B2(G317), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT52), .Z(new_n1102));
  AOI21_X1  g0902(.A(new_n395), .B1(new_n810), .B2(G322), .ZN(new_n1103));
  INV_X1    g0903(.A(G294), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n794), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n857), .B2(G303), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n394), .A2(new_n785), .B1(new_n802), .B2(new_n817), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n538), .B2(new_n790), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1102), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1100), .A2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1091), .B1(new_n779), .B2(new_n1110), .C1(new_n973), .C2(new_n831), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1087), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1086), .A2(new_n1112), .ZN(G390));
  NAND2_X1  g0913(.A1(new_n959), .A2(new_n961), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n820), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n802), .A2(new_n430), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n342), .B1(new_n810), .B2(G125), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n794), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n857), .B2(G137), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n787), .A2(G132), .B1(G159), .B2(new_n790), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n782), .A2(G128), .B1(new_n876), .B2(G50), .ZN(new_n1123));
  AND4_X1   g0923(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1094), .B1(G116), .B2(new_n787), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n817), .B2(new_n783), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n856), .A2(new_n394), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n342), .B1(new_n799), .B2(new_n1104), .C1(new_n794), .C2(new_n224), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n216), .A2(new_n785), .B1(new_n802), .B2(new_n218), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n778), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n777), .B1(new_n324), .B2(new_n851), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1115), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n721), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n918), .B2(new_n956), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1136), .A2(new_n1137), .B1(new_n953), .B2(new_n960), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n740), .A2(new_n741), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n733), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n743), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n700), .A3(new_n839), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n950), .B1(new_n1142), .B2(new_n952), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n960), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n957), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1138), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n765), .A2(KEYINPUT114), .A3(new_n842), .A4(new_n931), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n924), .A2(G330), .A3(new_n842), .A4(new_n931), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT114), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1138), .B(new_n1148), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n458), .A2(new_n766), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n951), .B1(new_n727), .B2(new_n839), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n924), .A2(G330), .A3(new_n842), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n950), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n1151), .B2(new_n1160), .ZN(new_n1161));
  AND4_X1   g0961(.A1(new_n952), .A2(new_n1142), .A3(new_n1160), .A4(new_n1148), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n964), .B(new_n1157), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1135), .B1(new_n1155), .B2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n656), .B(new_n1156), .C1(new_n745), .C2(new_n459), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n951), .B1(new_n744), .B2(new_n839), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1148), .A3(new_n1160), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1147), .A2(new_n1150), .B1(new_n950), .B2(new_n1159), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n1158), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1153), .A2(new_n1154), .A3(new_n1165), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1134), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n837), .A2(new_n838), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n699), .B(new_n1172), .C1(new_n742), .C2(new_n743), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n931), .B1(new_n1173), .B2(new_n951), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1145), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1144), .B1(new_n1158), .B2(new_n950), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1174), .A2(new_n1175), .B1(new_n1114), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1154), .B(new_n773), .C1(new_n1177), .C2(new_n1151), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT115), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT115), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1153), .A2(new_n1180), .A3(new_n773), .A4(new_n1154), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT116), .B1(new_n1171), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1154), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1175), .B1(new_n1166), .B2(new_n950), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1151), .B1(new_n1185), .B2(new_n1138), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1163), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n1170), .A3(new_n721), .ZN(new_n1188));
  AND4_X1   g0988(.A1(KEYINPUT116), .A2(new_n1182), .A3(new_n1188), .A4(new_n1133), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1183), .A2(new_n1189), .ZN(G378));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n433), .A2(new_n437), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n697), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n452), .A2(new_n456), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n452), .B2(new_n456), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n457), .A2(new_n1194), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1196), .A3(new_n1191), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n944), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n747), .B1(new_n1203), .B2(new_n957), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n935), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT40), .B1(new_n919), .B2(new_n932), .ZN(new_n1206));
  OAI21_X1  g1006(.A(G330), .B1(new_n943), .B2(new_n944), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n963), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT119), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n935), .A2(new_n1204), .A3(new_n1202), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n954), .A2(new_n962), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1208), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1210), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(KEYINPUT119), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n773), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n777), .B1(new_n434), .B2(new_n851), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n395), .A2(G41), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n817), .B2(new_n799), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1061), .B(new_n1221), .C1(G58), .C2(new_n876), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT117), .Z(new_n1223));
  OAI22_X1  g1023(.A1(new_n791), .A2(new_n216), .B1(new_n795), .B2(new_n224), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n394), .A2(new_n788), .B1(new_n783), .B2(new_n534), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n553), .C2(new_n808), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT118), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT58), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT58), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G33), .A2(G41), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1220), .A2(G50), .A3(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n795), .A2(new_n873), .B1(new_n794), .B2(new_n868), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1119), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n803), .B2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n782), .A2(G125), .B1(G150), .B2(new_n790), .ZN(new_n1236));
  INV_X1    g1036(.A(G128), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1235), .B(new_n1236), .C1(new_n1237), .C2(new_n788), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1239));
  INV_X1    g1039(.A(G124), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1231), .B1(new_n799), .B2(new_n1240), .C1(new_n785), .C2(new_n334), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1238), .B2(KEYINPUT59), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1232), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1229), .A2(new_n1230), .A3(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1219), .B1(new_n1244), .B2(new_n779), .C1(new_n821), .C2(new_n1208), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1218), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1170), .A2(new_n1165), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT57), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n964), .A2(new_n1157), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1148), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1138), .A2(new_n1256), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1257), .B2(new_n1169), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n721), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1247), .B1(new_n1250), .B2(new_n1259), .ZN(G375));
  NAND2_X1  g1060(.A1(new_n950), .A2(new_n820), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n774), .B1(G68), .B2(new_n852), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n817), .A2(new_n788), .B1(new_n783), .B2(new_n1104), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1023), .B(new_n1263), .C1(G97), .C2(new_n803), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n857), .A2(new_n538), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n794), .A2(new_n394), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n395), .B(new_n1266), .C1(G303), .C2(new_n810), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1063), .A3(new_n1265), .A4(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G132), .A2(new_n782), .B1(new_n787), .B2(G137), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n856), .B2(new_n1119), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(KEYINPUT121), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(KEYINPUT121), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n222), .A2(new_n785), .B1(new_n802), .B2(new_n334), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n395), .B1(new_n799), .B2(new_n1237), .C1(new_n794), .C2(new_n430), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(G50), .C2(new_n790), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1268), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1262), .B1(new_n1277), .B2(new_n778), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1169), .A2(new_n773), .B1(new_n1261), .B2(new_n1278), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n993), .B(KEYINPUT120), .Z(new_n1280));
  NAND2_X1  g1080(.A1(new_n1163), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(new_n1281), .B2(new_n1282), .ZN(G381));
  NAND3_X1  g1083(.A1(new_n1048), .A2(new_n833), .A3(new_n1082), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G390), .A2(new_n1284), .A3(G384), .A4(G381), .ZN(new_n1285));
  INV_X1    g1085(.A(G387), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1182), .A2(new_n1188), .A3(new_n1133), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1251), .B1(new_n1289), .B2(new_n1258), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1135), .B1(new_n1249), .B2(new_n1252), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1246), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1285), .A2(new_n1286), .A3(new_n1288), .A4(new_n1292), .ZN(G407));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1288), .A3(new_n698), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G407), .A2(G213), .A3(new_n1294), .ZN(G409));
  AND2_X1   g1095(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1245), .B1(new_n1296), .B2(new_n772), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1280), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1289), .A2(new_n1258), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1299), .B2(KEYINPUT123), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1248), .A2(new_n1249), .A3(new_n1280), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT123), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1287), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT122), .B1(G378), .B2(new_n1292), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT116), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1287), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1182), .A2(new_n1188), .A3(KEYINPUT116), .A4(new_n1133), .ZN(new_n1309));
  AND4_X1   g1109(.A1(KEYINPUT122), .A2(new_n1292), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1305), .B1(new_n1306), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  INV_X1    g1112(.A(G213), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(G343), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n1312), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT122), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(G375), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1292), .A2(KEYINPUT122), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1304), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT125), .B1(new_n1321), .B2(new_n1314), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1314), .A2(G2897), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1163), .A2(KEYINPUT60), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1282), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n721), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1325), .A2(new_n1282), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1279), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n850), .A3(new_n882), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G384), .B(new_n1279), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT124), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1324), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1332), .B(new_n1333), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1334), .B1(new_n1335), .B2(new_n1324), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1332), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1316), .A2(new_n1322), .A3(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1332), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1311), .A2(new_n1315), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1337), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G393), .A2(G396), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1284), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1016), .A2(new_n1042), .A3(G390), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(G390), .B1(new_n1016), .B2(new_n1042), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1347), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1350), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1347), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1352), .A2(new_n1353), .A3(new_n1348), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1351), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1345), .A2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(KEYINPUT61), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1316), .A2(new_n1322), .A3(KEYINPUT63), .A4(new_n1341), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT63), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1342), .A2(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1336), .B1(new_n1314), .B2(new_n1321), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1357), .A2(new_n1358), .A3(new_n1360), .A4(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1356), .A2(new_n1362), .ZN(G405));
  OR2_X1    g1163(.A1(new_n1355), .A2(KEYINPUT127), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1355), .A2(KEYINPUT127), .ZN(new_n1365));
  OR2_X1    g1165(.A1(new_n1341), .A2(KEYINPUT126), .ZN(new_n1366));
  OAI22_X1  g1166(.A1(new_n1306), .A2(new_n1310), .B1(new_n1287), .B2(new_n1292), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1332), .B(KEYINPUT126), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1369), .A2(new_n1367), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  NAND4_X1  g1171(.A1(new_n1364), .A2(new_n1365), .A3(new_n1368), .A4(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1368), .ZN(new_n1373));
  OAI211_X1 g1173(.A(new_n1355), .B(KEYINPUT127), .C1(new_n1373), .C2(new_n1370), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1372), .A2(new_n1374), .ZN(G402));
endmodule


