//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G113), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n470), .B2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n465), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AOI21_X1  g057(.A(new_n464), .B1(new_n475), .B2(new_n477), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n478), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND3_X1   g064(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT3), .B1(new_n476), .B2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n470), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n495), .A2(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n475), .A2(new_n477), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n501), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n494), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G50), .A3(G543), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n507), .A2(new_n509), .A3(new_n515), .A4(new_n517), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n514), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n518), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n521), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(G51), .B1(G89), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n507), .A2(new_n509), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n526), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(G64), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n539), .B1(new_n542), .B2(G651), .ZN(new_n543));
  AOI211_X1 g118(.A(KEYINPUT70), .B(new_n513), .C1(new_n540), .C2(new_n541), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n537), .B(new_n538), .C1(new_n543), .C2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND3_X1  g121(.A1(new_n511), .A2(new_n518), .A3(G81), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n518), .A2(G43), .A3(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT71), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n530), .B2(new_n532), .ZN(new_n555));
  INV_X1    g130(.A(G68), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n506), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND3_X1  g141(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n518), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n510), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n526), .A2(G91), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(G299));
  OAI221_X1 g152(.A(new_n519), .B1(new_n520), .B2(new_n521), .C1(new_n512), .C2(new_n513), .ZN(G303));
  NAND4_X1  g153(.A1(new_n511), .A2(new_n518), .A3(KEYINPUT72), .A4(G87), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n521), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n525), .A2(G49), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n530), .A2(new_n585), .A3(new_n532), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(G288));
  NAND3_X1  g163(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n513), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n511), .A2(new_n518), .A3(G86), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n515), .A2(new_n517), .A3(G48), .A4(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n533), .A2(G60), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n513), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n524), .A2(new_n600), .B1(new_n601), .B2(new_n521), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n521), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n510), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n606), .A2(new_n609), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n518), .A2(new_n615), .A3(G543), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(G54), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(KEYINPUT74), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(KEYINPUT74), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n605), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n605), .B1(new_n621), .B2(G868), .ZN(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(G299), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G168), .B2(new_n624), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(G168), .B2(new_n624), .ZN(G280));
  INV_X1    g202(.A(new_n621), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G559), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G860), .B2(new_n621), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT75), .ZN(G148));
  NAND2_X1  g207(.A1(new_n559), .A2(new_n624), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n630), .B2(new_n624), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n462), .A2(new_n479), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2100), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n478), .A2(G135), .ZN(new_n640));
  NOR2_X1   g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(G123), .B2(new_n483), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2435), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2438), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n652), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT76), .Z(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT77), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n665), .B(KEYINPUT17), .Z(new_n668));
  OAI21_X1  g243(.A(new_n667), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n663), .A3(new_n661), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n665), .A3(new_n661), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n682), .A2(KEYINPUT20), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n678), .A3(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(KEYINPUT20), .C2(new_n682), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT78), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G21), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G286), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1966), .ZN(new_n700));
  INV_X1    g275(.A(G28), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n701), .B2(KEYINPUT30), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n644), .A2(G29), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT27), .B(G1996), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT89), .B1(G29), .B2(G32), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n478), .A2(G141), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n483), .A2(G129), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n479), .A2(G105), .ZN(new_n713));
  AND4_X1   g288(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  MUX2_X1   g290(.A(KEYINPUT89), .B(new_n708), .S(new_n715), .Z(new_n716));
  AOI21_X1  g291(.A(new_n705), .B1(new_n707), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G19), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G16), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n559), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1341), .Z(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2078), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n727), .A2(new_n728), .A3(G29), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n481), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT88), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2084), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n717), .A2(new_n726), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G20), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT23), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT23), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n738), .B2(new_n735), .ZN(new_n739));
  INV_X1    g314(.A(G1956), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n722), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n722), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT92), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT92), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n744), .A2(KEYINPUT29), .A3(new_n745), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n748), .A2(G2090), .A3(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n741), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n733), .B1(KEYINPUT94), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  NOR2_X1   g329(.A1(G5), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G171), .B2(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G1961), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT90), .Z(new_n758));
  NAND4_X1  g333(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n483), .A2(G128), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n478), .A2(G140), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT83), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(KEYINPUT83), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n722), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n722), .A2(G26), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT28), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT28), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G2067), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n748), .A2(new_n749), .ZN(new_n774));
  INV_X1    g349(.A(G2090), .ZN(new_n775));
  AOI21_X1  g350(.A(KEYINPUT93), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n774), .A2(KEYINPUT93), .A3(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n478), .A2(G139), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n479), .A2(G103), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT85), .Z(new_n783));
  OAI211_X1 g358(.A(new_n778), .B(new_n781), .C1(new_n783), .C2(new_n464), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT86), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT86), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT87), .ZN(new_n787));
  AOI21_X1  g362(.A(KEYINPUT87), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g363(.A(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2072), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G33), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AND3_X1   g367(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(new_n789), .B2(new_n792), .ZN(new_n794));
  OAI221_X1 g369(.A(new_n773), .B1(new_n776), .B2(new_n777), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n756), .A2(G1961), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n716), .A2(new_n707), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n731), .A2(G2084), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n759), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G23), .B(G288), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT33), .ZN(new_n803));
  INV_X1    g378(.A(G1976), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  INV_X1    g382(.A(G1981), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  MUX2_X1   g386(.A(G22), .B(G303), .S(G16), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT81), .B(G1971), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n803), .A2(new_n804), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n810), .A2(new_n811), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G24), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G290), .B2(G16), .ZN(new_n819));
  MUX2_X1   g394(.A(new_n818), .B(new_n819), .S(KEYINPUT80), .Z(new_n820));
  INV_X1    g395(.A(G1986), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n805), .A2(new_n809), .A3(new_n814), .A4(new_n815), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n820), .A2(new_n821), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n722), .A2(G25), .ZN(new_n826));
  OR2_X1    g401(.A1(G95), .A2(G2105), .ZN(new_n827));
  INV_X1    g402(.A(G107), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n470), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n478), .A2(G131), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n483), .A2(G119), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n826), .B1(new_n833), .B2(new_n722), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G1991), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT79), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n825), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n816), .A2(new_n822), .A3(new_n824), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  AOI211_X1 g417(.A(new_n825), .B(new_n839), .C1(new_n823), .C2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n822), .A4(new_n816), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(G4), .A2(G16), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n621), .B2(G16), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT82), .B(G1348), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n801), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT95), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n801), .A2(new_n846), .A3(new_n853), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G311));
  NAND2_X1  g430(.A1(new_n851), .A2(KEYINPUT96), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n801), .A2(new_n846), .A3(new_n857), .A4(new_n850), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(G150));
  NAND2_X1  g434(.A1(new_n533), .A2(G67), .ZN(new_n860));
  INV_X1    g435(.A(G80), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n506), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G651), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n525), .A2(G55), .B1(G93), .B2(new_n526), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n621), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n871));
  INV_X1    g446(.A(new_n552), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n551), .B1(new_n547), .B2(new_n548), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n558), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n553), .A2(KEYINPUT97), .A3(new_n558), .ZN(new_n877));
  INV_X1    g452(.A(new_n864), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n862), .B2(G651), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n865), .A2(new_n871), .A3(new_n559), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n870), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n867), .B1(new_n884), .B2(G860), .ZN(G145));
  XNOR2_X1  g460(.A(new_n481), .B(new_n488), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n644), .ZN(new_n887));
  INV_X1    g462(.A(new_n714), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n765), .A2(new_n766), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G164), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(G164), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n714), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n787), .B2(new_n788), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n785), .A2(new_n786), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n833), .B(new_n637), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n483), .A2(G130), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n478), .A2(G142), .ZN(new_n902));
  NOR2_X1   g477(.A1(G106), .A2(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n900), .B(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n897), .A2(new_n899), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n897), .B2(new_n899), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n887), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n907), .A2(new_n908), .A3(new_n887), .ZN(new_n912));
  OAI211_X1 g487(.A(KEYINPUT98), .B(new_n887), .C1(new_n907), .C2(new_n908), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g490(.A1(new_n865), .A2(new_n624), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n629), .B(new_n883), .ZN(new_n917));
  INV_X1    g492(.A(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n618), .ZN(new_n919));
  NAND3_X1  g494(.A1(G299), .A2(new_n617), .A3(new_n613), .ZN(new_n920));
  AOI211_X1 g495(.A(KEYINPUT99), .B(KEYINPUT41), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n924), .B2(KEYINPUT99), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n920), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n917), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n599), .A2(G303), .A3(new_n603), .ZN(new_n930));
  OAI21_X1  g505(.A(G166), .B1(new_n598), .B2(new_n602), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(G305), .ZN(new_n932));
  AOI21_X1  g507(.A(G305), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(G288), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(G305), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G288), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n930), .A2(new_n931), .A3(G305), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n934), .A2(new_n940), .A3(KEYINPUT100), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  MUX2_X1   g520(.A(new_n941), .B(new_n945), .S(KEYINPUT42), .Z(new_n946));
  XNOR2_X1  g521(.A(new_n929), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n916), .B1(new_n947), .B2(new_n624), .ZN(G295));
  OAI21_X1  g523(.A(new_n916), .B1(new_n947), .B2(new_n624), .ZN(G331));
  XOR2_X1   g524(.A(G286), .B(KEYINPUT101), .Z(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n880), .A2(G301), .A3(new_n881), .ZN(new_n952));
  AOI21_X1  g527(.A(G301), .B1(new_n880), .B2(new_n881), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n882), .A2(G171), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n880), .A2(G301), .A3(new_n881), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n950), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n958));
  INV_X1    g533(.A(new_n924), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n960), .A2(new_n945), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n952), .A2(new_n953), .A3(new_n951), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n928), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n957), .A3(new_n959), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(KEYINPUT104), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n934), .A2(new_n940), .A3(KEYINPUT100), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT100), .B1(new_n934), .B2(new_n940), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n954), .A2(new_n925), .A3(new_n957), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT105), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n961), .A2(new_n966), .A3(KEYINPUT105), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT102), .B1(new_n943), .B2(new_n944), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n954), .A2(new_n925), .A3(new_n957), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n954), .A2(new_n957), .B1(new_n919), .B2(new_n920), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n968), .B2(new_n969), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n964), .A2(new_n984), .A3(new_n971), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n985), .A3(new_n976), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT103), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n989), .A3(KEYINPUT43), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n978), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND4_X1   g568(.A1(KEYINPUT43), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n986), .A2(new_n975), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT44), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(G397));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n504), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n465), .A2(new_n473), .A3(G40), .A4(new_n480), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n889), .B(new_n772), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n833), .A2(new_n837), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n714), .B(G1996), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n833), .A2(new_n837), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G290), .A2(G1986), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n1003), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT48), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1003), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(G1996), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT46), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1004), .B2(new_n714), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1005), .B1(new_n1020), .B2(new_n1003), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n772), .B2(new_n767), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT127), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1013), .B(new_n1019), .C1(new_n1003), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT63), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT108), .B(G8), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n503), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT68), .B1(new_n483), .B2(G126), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n495), .A2(new_n496), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n499), .A2(new_n497), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n502), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  AND4_X1   g609(.A1(G40), .A2(new_n465), .A3(new_n480), .A4(new_n473), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1027), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n592), .A2(new_n808), .A3(new_n593), .A4(new_n594), .ZN(new_n1037));
  INV_X1    g612(.A(G86), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n594), .B1(new_n521), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1039), .B2(new_n591), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1040), .A3(KEYINPUT110), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT49), .B1(new_n1041), .B2(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g617(.A1(KEYINPUT111), .A2(KEYINPUT49), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1037), .A2(new_n1040), .B1(KEYINPUT110), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1036), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n583), .A2(new_n584), .A3(new_n587), .A4(G1976), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1026), .C1(new_n999), .C2(new_n1002), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT52), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT109), .B(G1976), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1049), .A2(new_n1051), .A3(new_n1026), .A4(new_n1046), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1048), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT117), .ZN(new_n1054));
  INV_X1    g629(.A(G1971), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n504), .B2(new_n998), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT106), .ZN(new_n1059));
  NOR4_X1   g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1002), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1002), .B1(new_n999), .B2(new_n1000), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT106), .B1(new_n1061), .B2(new_n1056), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1002), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n504), .A2(new_n1065), .A3(new_n998), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT107), .B(G2090), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1063), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G166), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(new_n1073), .B(KEYINPUT55), .Z(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(G8), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(new_n1035), .C1(new_n1034), .C2(new_n1065), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1065), .B1(new_n504), .B2(new_n998), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT116), .B1(new_n1079), .B2(new_n1002), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1080), .A3(new_n1066), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(new_n1068), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1027), .B1(new_n1082), .B2(new_n1063), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1054), .B(new_n1076), .C1(new_n1075), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1064), .A2(new_n1085), .A3(new_n1066), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1035), .C1(new_n1034), .C2(KEYINPUT45), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n1058), .B2(new_n1002), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1057), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1090), .B2(G1966), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(G168), .A3(new_n1026), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1025), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1075), .B1(new_n1071), .B2(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1053), .A2(KEYINPUT112), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1045), .A2(new_n1097), .A3(new_n1048), .A4(new_n1052), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1095), .A2(new_n1099), .A3(new_n1092), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1076), .A2(KEYINPUT63), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1094), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1001), .A2(new_n1035), .A3(new_n1056), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1059), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1061), .A2(KEYINPUT106), .A3(new_n1056), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1971), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1107), .B2(new_n1069), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1074), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1086), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1087), .B1(new_n1001), .B2(new_n1035), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1058), .A2(KEYINPUT118), .A3(new_n1002), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1056), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1966), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1111), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1116), .A2(G286), .A3(new_n1027), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1109), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1118), .A2(KEYINPUT119), .A3(new_n1101), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1093), .B1(new_n1103), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1076), .A2(new_n1099), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1037), .B(KEYINPUT114), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n938), .A2(new_n804), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT115), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1045), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1036), .B(KEYINPUT113), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1120), .A2(new_n1121), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G286), .A2(new_n1026), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1091), .B2(new_n1026), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1116), .B2(new_n1072), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(KEYINPUT51), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1091), .A2(KEYINPUT124), .A3(new_n1131), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT124), .B1(new_n1091), .B2(new_n1131), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT126), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(KEYINPUT62), .C1(new_n1135), .C2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(G1961), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1144));
  INV_X1    g719(.A(G2078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1105), .A2(new_n1145), .A3(new_n1106), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1090), .A2(KEYINPUT53), .A3(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(G301), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(KEYINPUT62), .ZN(new_n1152));
  INV_X1    g727(.A(G1348), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1067), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  INV_X1    g730(.A(new_n618), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n999), .A2(new_n1002), .A3(G2067), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n618), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1156), .B(new_n1157), .C1(new_n1067), .C2(new_n1153), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT60), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT121), .B(G1996), .Z(new_n1163));
  NAND4_X1  g738(.A1(new_n1001), .A2(new_n1035), .A3(new_n1056), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT122), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT58), .B(G1341), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1049), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1061), .A2(new_n1168), .A3(new_n1056), .A4(new_n1163), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n560), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1170), .B2(new_n560), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1159), .B(new_n1162), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1081), .A2(new_n740), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1104), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT56), .B(G2072), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G299), .B(KEYINPUT57), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1175), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1180), .A2(KEYINPUT123), .A3(new_n1181), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1081), .A2(new_n740), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1181), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1184), .A2(new_n1185), .B1(new_n1186), .B2(KEYINPUT61), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(KEYINPUT120), .A3(new_n1185), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1182), .A2(new_n1183), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT61), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1174), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1191), .A2(new_n1160), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1194), .A2(new_n1182), .A3(new_n1188), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1151), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(G40), .B1(new_n463), .B2(new_n464), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1197), .A2(new_n1147), .A3(G2078), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1001), .A2(new_n480), .A3(new_n1056), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI211_X1 g775(.A(new_n1144), .B(new_n1200), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1201));
  OAI21_X1  g776(.A(KEYINPUT125), .B1(new_n1201), .B2(G301), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1148), .A2(new_n1199), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1203), .A2(new_n1204), .A3(G171), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1148), .A2(G301), .A3(new_n1149), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1201), .A2(G301), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1150), .A2(KEYINPUT54), .ZN(new_n1209));
  AOI22_X1  g784(.A1(new_n1207), .A2(KEYINPUT54), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI22_X1  g785(.A1(new_n1143), .A2(new_n1152), .B1(new_n1196), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1084), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1129), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g788(.A(new_n1008), .B(new_n1007), .C1(G1986), .C2(G290), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1010), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1014), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1024), .B1(new_n1213), .B2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g792(.A1(G401), .A2(new_n460), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n914), .A2(new_n675), .A3(new_n1219), .ZN(new_n1220));
  AND3_X1   g794(.A1(new_n1220), .A2(new_n991), .A3(new_n695), .ZN(G308));
  NAND3_X1  g795(.A1(new_n1220), .A2(new_n991), .A3(new_n695), .ZN(G225));
endmodule


