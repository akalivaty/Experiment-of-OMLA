//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n205), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT89), .B(G197gat), .Z(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n206), .B2(new_n207), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT12), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT12), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n210), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(G8gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT16), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n221), .A2(G1gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n219), .B(new_n220), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G15gat), .B(G22gat), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n222), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n223), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n228), .A2(new_n229), .A3(new_n218), .A4(G8gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT90), .ZN(new_n233));
  OR3_X1    g032(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(new_n234), .ZN(new_n237));
  AND2_X1   g036(.A1(G43gat), .A2(G50gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(G43gat), .A2(G50gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT15), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G43gat), .ZN(new_n241));
  INV_X1    g040(.A(G50gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT15), .ZN(new_n244));
  NAND2_X1  g043(.A1(G43gat), .A2(G50gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G29gat), .A2(G36gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n240), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n232), .ZN(new_n249));
  NOR3_X1   g048(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n237), .A2(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n252), .ZN(new_n255));
  NOR4_X1   g054(.A1(new_n236), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n234), .B2(new_n233), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n246), .A3(new_n247), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT17), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n259), .A2(KEYINPUT91), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT91), .B1(new_n259), .B2(new_n260), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n231), .B(new_n254), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n231), .A2(KEYINPUT93), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n226), .A2(new_n266), .A3(new_n230), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n263), .A2(KEYINPUT18), .A3(new_n264), .A4(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n264), .B(KEYINPUT13), .Z(new_n270));
  INV_X1    g069(.A(new_n267), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n226), .B2(new_n230), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n271), .A2(new_n272), .A3(new_n253), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n259), .B1(new_n265), .B2(new_n267), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n263), .A2(new_n264), .A3(new_n268), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT18), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n217), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  AND4_X1   g079(.A1(new_n279), .A2(new_n269), .A3(new_n275), .A4(new_n217), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G113gat), .B(G120gat), .Z(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT64), .B(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT23), .A3(new_n205), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  OR2_X1    g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n291), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT65), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT65), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(new_n291), .C1(new_n298), .C2(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(G169gat), .A3(G176gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(new_n311), .C1(new_n295), .C2(new_n296), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT67), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n297), .A2(KEYINPUT25), .ZN(new_n314));
  INV_X1    g113(.A(new_n301), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT68), .B(G190gat), .Z(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n306), .A3(new_n308), .A4(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n295), .B(KEYINPUT26), .Z(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n294), .ZN(new_n323));
  INV_X1    g122(.A(new_n316), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT27), .B(G183gat), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT28), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n324), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n299), .B(new_n323), .C1(new_n330), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n321), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n304), .A2(KEYINPUT65), .B1(new_n313), .B2(new_n319), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n306), .B1(new_n335), .B2(new_n308), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n290), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G227gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n305), .A2(new_n308), .A3(new_n320), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT69), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n288), .A2(new_n289), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n321), .A4(new_n333), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n337), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT32), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT33), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT71), .ZN(new_n350));
  XOR2_X1   g149(.A(G71gat), .B(G99gat), .Z(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n345), .B(KEYINPUT32), .C1(new_n347), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n344), .ZN(new_n357));
  INV_X1    g156(.A(new_n340), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT34), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT34), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n353), .A2(new_n355), .B1(new_n360), .B2(new_n362), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT72), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n340), .B1(new_n337), .B2(new_n344), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT34), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n353), .A3(new_n355), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n366), .A2(KEYINPUT36), .A3(new_n368), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT36), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n363), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(new_n367), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G197gat), .B(G204gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n378));
  INV_X1    g177(.A(G211gat), .ZN(new_n379));
  INV_X1    g178(.A(G218gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT74), .ZN(new_n385));
  INV_X1    g184(.A(G155gat), .ZN(new_n386));
  INV_X1    g185(.A(G162gat), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT2), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G141gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G148gat), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT77), .B(G148gat), .Z(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n391), .ZN(new_n394));
  XNOR2_X1  g193(.A(G155gat), .B(G162gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  INV_X1    g196(.A(G148gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G141gat), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT2), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(new_n395), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n396), .A2(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n403), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n397), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n385), .A2(new_n404), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G78gat), .B(G106gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT83), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT31), .B(G50gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n408), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n414), .B(G22gat), .Z(new_n415));
  OR2_X1    g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n415), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n385), .ZN(new_n419));
  INV_X1    g218(.A(G226gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n339), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n334), .A2(new_n336), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n341), .A2(new_n333), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n421), .A2(KEYINPUT29), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n419), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n334), .B2(new_n336), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n341), .A2(new_n333), .A3(new_n421), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n385), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n427), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT75), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n427), .A2(new_n430), .A3(new_n437), .A4(new_n434), .ZN(new_n438));
  XOR2_X1   g237(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n430), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n342), .A2(new_n321), .A3(new_n333), .A4(new_n421), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n425), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n385), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n433), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT30), .A4(new_n434), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT84), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n440), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n290), .A2(new_n396), .A3(new_n401), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n343), .A2(KEYINPUT79), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n288), .A2(new_n457), .A3(new_n289), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n459), .A3(new_n402), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n454), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464));
  OR3_X1    g263(.A1(new_n463), .A2(KEYINPUT39), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT0), .ZN(new_n467));
  XNOR2_X1  g266(.A(G57gat), .B(G85gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  NOR2_X1   g268(.A1(new_n405), .A2(new_n343), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n405), .B2(new_n459), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT39), .B(new_n472), .C1(new_n463), .C2(new_n464), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n474), .A2(new_n475), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n290), .A2(KEYINPUT4), .A3(new_n396), .A4(new_n401), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n453), .B1(new_n405), .B2(new_n343), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n478), .A3(new_n479), .A4(new_n464), .ZN(new_n480));
  INV_X1    g279(.A(new_n458), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n457), .B1(new_n288), .B2(new_n289), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n405), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n452), .ZN(new_n484));
  INV_X1    g283(.A(new_n464), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT5), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n485), .A2(KEYINPUT5), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n454), .A2(new_n460), .A3(new_n462), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n469), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n476), .A2(new_n477), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n449), .A2(new_n451), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT5), .B1(new_n471), .B2(new_n464), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n485), .B1(new_n452), .B2(new_n453), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n460), .A2(new_n494), .A3(new_n478), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n469), .B(new_n489), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT85), .B1(new_n498), .B2(new_n490), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n427), .A2(new_n430), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n434), .B1(new_n505), .B2(KEYINPUT37), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n436), .A2(new_n438), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n385), .B1(new_n423), .B2(new_n426), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n428), .A2(new_n429), .A3(new_n419), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT37), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n434), .A2(new_n509), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n514), .B(new_n515), .C1(new_n505), .C2(new_n507), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n504), .A2(new_n510), .A3(new_n511), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n418), .B1(new_n492), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n490), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g319(.A(new_n498), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT81), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n490), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .A4(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n502), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n498), .B1(new_n522), .B2(new_n490), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT82), .B1(new_n526), .B2(new_n520), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n440), .B(new_n447), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n418), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n376), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n366), .A2(new_n368), .A3(new_n371), .A4(new_n529), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT35), .B1(new_n532), .B2(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n449), .A2(new_n451), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT88), .B1(new_n374), .B2(new_n367), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n364), .A2(new_n536), .A3(new_n371), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT35), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n416), .A2(new_n538), .A3(new_n417), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n499), .A2(new_n500), .B1(KEYINPUT6), .B2(new_n490), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n503), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n534), .A2(new_n535), .A3(new_n537), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n282), .B1(new_n531), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G183gat), .B(G211gat), .Z(new_n545));
  XOR2_X1   g344(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n546));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(G57gat), .A2(G64gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G57gat), .A2(G64gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n548), .ZN(new_n554));
  NOR2_X1   g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n547), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(G57gat), .A2(G64gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT94), .A4(new_n550), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n550), .B2(new_n560), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n568), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n571), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n546), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n564), .B1(new_n557), .B2(new_n562), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n265), .A2(new_n267), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n570), .A2(new_n571), .ZN(new_n582));
  INV_X1    g381(.A(new_n546), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n577), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n577), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n545), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n577), .A2(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n579), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n577), .A2(new_n580), .A3(new_n584), .ZN(new_n590));
  INV_X1    g389(.A(new_n545), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT8), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n597), .A2(new_n600), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n606), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n237), .A2(new_n248), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n255), .ZN(new_n616));
  INV_X1    g415(.A(G232gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n339), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n595), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  OAI221_X1 g421(.A(KEYINPUT99), .B1(new_n620), .B2(new_n619), .C1(new_n253), .C2(new_n614), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n614), .B(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n626), .B(new_n254), .C1(new_n261), .C2(new_n262), .ZN(new_n627));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n624), .B2(new_n627), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT97), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT96), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n630), .B2(new_n631), .ZN(new_n639));
  OAI211_X1 g438(.A(KEYINPUT97), .B(new_n636), .C1(new_n630), .C2(new_n631), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n638), .B2(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n605), .A2(new_n607), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n578), .A2(new_n653), .A3(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT102), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n578), .A2(new_n653), .A3(new_n656), .A4(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n566), .A2(new_n614), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n578), .A2(new_n653), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n650), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n661), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n650), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT103), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n667), .A3(new_n650), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n663), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n648), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n648), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n666), .A2(new_n668), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT104), .B(new_n672), .C1(new_n673), .C2(new_n663), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n594), .A2(new_n645), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n544), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n524), .A2(new_n502), .ZN(new_n679));
  INV_X1    g478(.A(new_n527), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n222), .ZN(G1324gat));
  AND3_X1   g482(.A1(new_n440), .A2(new_n447), .A3(new_n450), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n450), .B1(new_n440), .B2(new_n447), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n544), .A2(new_n686), .A3(new_n677), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G8gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  MUX2_X1   g490(.A(new_n689), .B(KEYINPUT42), .S(new_n691), .Z(G1325gat));
  OAI21_X1  g491(.A(G15gat), .B1(new_n678), .B2(new_n376), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n535), .A2(new_n537), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n678), .B2(new_n695), .ZN(G1326gat));
  NOR2_X1   g495(.A1(new_n678), .A2(new_n529), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  NOR3_X1   g498(.A1(new_n593), .A2(new_n644), .A3(new_n676), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n544), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(G29gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n681), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n593), .B(KEYINPUT105), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(new_n282), .A3(new_n676), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n531), .A2(new_n543), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n645), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n371), .B1(new_n367), .B2(KEYINPUT72), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n356), .A2(KEYINPUT72), .A3(new_n363), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(new_n714), .A3(new_n418), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n448), .B1(new_n679), .B2(new_n680), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n538), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n535), .A2(new_n541), .A3(new_n537), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n686), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT106), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n533), .A2(new_n542), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n531), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n645), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n709), .B1(new_n712), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n681), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n705), .A2(new_n728), .ZN(G1328gat));
  INV_X1    g528(.A(G36gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n701), .A2(new_n730), .A3(new_n686), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT46), .Z(new_n732));
  OAI21_X1  g531(.A(G36gat), .B1(new_n727), .B2(new_n534), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1329gat));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n376), .B(new_n709), .C1(new_n712), .C2(new_n725), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n241), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n701), .A2(new_n241), .A3(new_n535), .A4(new_n537), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n736), .B2(new_n241), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI221_X1 g540(.A(new_n738), .B1(new_n735), .B2(KEYINPUT47), .C1(new_n736), .C2(new_n241), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1330gat));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  AND4_X1   g543(.A1(new_n242), .A2(new_n544), .A3(new_n418), .A4(new_n700), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n723), .A2(new_n645), .A3(new_n724), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n710), .B2(new_n645), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n418), .B(new_n708), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(G50gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n744), .B1(new_n750), .B2(KEYINPUT109), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n242), .B1(new_n726), .B2(new_n418), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n752), .B(KEYINPUT48), .C1(new_n753), .C2(new_n745), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n751), .A2(new_n754), .ZN(G1331gat));
  NAND3_X1  g554(.A1(new_n593), .A2(new_n644), .A3(new_n282), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n675), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n723), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n703), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n686), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n762), .B2(new_n761), .ZN(G1333gat));
  XOR2_X1   g564(.A(new_n694), .B(KEYINPUT110), .Z(new_n766));
  AND2_X1   g565(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n767), .A2(G71gat), .ZN(new_n768));
  INV_X1    g567(.A(new_n376), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n758), .A2(G71gat), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n768), .B2(new_n770), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n418), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT112), .B(G78gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1335gat));
  AND2_X1   g576(.A1(new_n277), .A2(new_n278), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n269), .A2(new_n275), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n213), .B(new_n216), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n276), .A2(new_n279), .A3(new_n217), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n593), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n723), .A2(new_n645), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n645), .A4(new_n783), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n675), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n601), .A3(new_n703), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n676), .B(new_n783), .C1(new_n746), .C2(new_n748), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT113), .B1(new_n790), .B2(new_n681), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G85gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n790), .A2(KEYINPUT113), .A3(new_n681), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  NAND2_X1  g593(.A1(new_n686), .A2(G92gat), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n534), .B(new_n675), .C1(new_n786), .C2(new_n787), .ZN(new_n796));
  OAI221_X1 g595(.A(KEYINPUT52), .B1(new_n790), .B2(new_n795), .C1(new_n796), .C2(G92gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  AOI21_X1  g597(.A(G92gat), .B1(new_n788), .B2(new_n686), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n790), .A2(new_n795), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1337gat));
  INV_X1    g601(.A(G99gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n790), .A2(new_n803), .A3(new_n376), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n535), .A3(new_n537), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n803), .ZN(G1338gat));
  NAND2_X1  g605(.A1(new_n418), .A2(G106gat), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n529), .B(new_n675), .C1(new_n786), .C2(new_n787), .ZN(new_n808));
  OAI221_X1 g607(.A(KEYINPUT53), .B1(new_n790), .B2(new_n807), .C1(new_n808), .C2(G106gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g609(.A(G106gat), .B1(new_n788), .B2(new_n418), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n790), .A2(new_n807), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(G1339gat));
  NOR2_X1   g613(.A1(new_n756), .A2(new_n676), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n658), .A2(new_n662), .A3(new_n650), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n818), .A2(new_n663), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n658), .A2(new_n662), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n819), .A3(new_n649), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n648), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n669), .A2(new_n672), .ZN(new_n825));
  INV_X1    g624(.A(new_n663), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n658), .A2(new_n662), .A3(new_n650), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n672), .B1(new_n663), .B2(new_n819), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n273), .A2(new_n274), .A3(new_n270), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n264), .B1(new_n263), .B2(new_n268), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n833), .A2(new_n834), .B1(new_n211), .B2(new_n212), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n781), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n832), .B(new_n836), .C1(new_n641), .C2(new_n643), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n671), .A2(new_n781), .A3(new_n674), .A4(new_n835), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n838), .B(new_n839), .C1(new_n831), .C2(new_n282), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n644), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n782), .A2(new_n825), .A3(new_n830), .A4(new_n824), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n839), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT115), .B(new_n837), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n706), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n839), .B1(new_n831), .B2(new_n282), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n644), .A3(new_n840), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT115), .B1(new_n848), .B2(new_n837), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n816), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n686), .A2(new_n681), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n715), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n782), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n529), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT116), .ZN(new_n857));
  AND4_X1   g656(.A1(new_n535), .A2(new_n857), .A3(new_n537), .A4(new_n851), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n782), .A2(G113gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  AOI21_X1  g659(.A(G120gat), .B1(new_n854), .B2(new_n676), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n676), .A2(G120gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(G1341gat));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n853), .A2(new_n864), .A3(new_n594), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT117), .B1(new_n854), .B2(new_n593), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n865), .A2(G127gat), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n707), .A2(G127gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n858), .B2(new_n868), .ZN(G1342gat));
  AND2_X1   g668(.A1(new_n850), .A2(new_n703), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n534), .A2(new_n645), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT118), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(G134gat), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n870), .A2(new_n873), .A3(new_n874), .A4(new_n715), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT56), .Z(new_n876));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n645), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n874), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n850), .A2(new_n881), .A3(new_n418), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n851), .A2(new_n376), .ZN(new_n883));
  XOR2_X1   g682(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n820), .B2(new_n823), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n825), .A3(new_n830), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n839), .B1(new_n886), .B2(new_n282), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n839), .C1(new_n886), .C2(new_n282), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n644), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n593), .B1(new_n891), .B2(new_n837), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n418), .B1(new_n892), .B2(new_n815), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n882), .A2(new_n894), .A3(new_n782), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n769), .A2(new_n529), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n282), .A2(G141gat), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n850), .A2(new_n897), .A3(new_n851), .A4(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT121), .B1(new_n901), .B2(KEYINPUT58), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n895), .B2(G141gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n896), .A2(new_n905), .A3(new_n900), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n903), .A2(KEYINPUT122), .A3(new_n905), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n880), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n901), .A2(KEYINPUT121), .A3(KEYINPUT58), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n916), .A2(KEYINPUT123), .A3(new_n910), .A4(new_n911), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1344gat));
  AND2_X1   g717(.A1(new_n870), .A2(new_n897), .ZN(new_n919));
  INV_X1    g718(.A(new_n393), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n534), .A4(new_n676), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n850), .A2(new_n418), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT57), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n893), .A2(new_n881), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n675), .B(new_n883), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n398), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n676), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT124), .B1(new_n930), .B2(new_n883), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n922), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n882), .A2(new_n894), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n675), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(KEYINPUT59), .A3(new_n920), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n921), .B1(new_n932), .B2(new_n935), .ZN(G1345gat));
  NOR3_X1   g735(.A1(new_n933), .A2(new_n386), .A3(new_n706), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n852), .A2(new_n593), .A3(new_n897), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n386), .B2(new_n938), .ZN(G1346gat));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n387), .A3(new_n873), .ZN(new_n940));
  OAI21_X1  g739(.A(G162gat), .B1(new_n933), .B2(new_n644), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n703), .A2(new_n534), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n850), .A2(new_n715), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G169gat), .B1(new_n944), .B2(new_n782), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n766), .A2(new_n943), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT125), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n857), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n282), .A2(new_n205), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1348gat));
  AOI21_X1  g749(.A(G176gat), .B1(new_n944), .B2(new_n676), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n675), .A2(new_n292), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n948), .B2(new_n952), .ZN(G1349gat));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n707), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G183gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n594), .A2(new_n328), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g756(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n317), .B1(new_n948), .B2(new_n707), .ZN(new_n961));
  INV_X1    g760(.A(new_n957), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(G1350gat));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n645), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G190gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n965), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n944), .A2(new_n316), .A3(new_n645), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT127), .Z(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(G1351gat));
  AND3_X1   g771(.A1(new_n923), .A2(new_n376), .A3(new_n943), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n782), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n943), .A2(new_n376), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n924), .B2(new_n925), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n782), .A2(G197gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  INV_X1    g777(.A(G204gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n979), .A3(new_n676), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT62), .Z(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n930), .B2(new_n975), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n973), .A2(new_n379), .A3(new_n593), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n379), .B1(new_n976), .B2(new_n593), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(KEYINPUT63), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n380), .A3(new_n645), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n976), .A2(new_n645), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n380), .ZN(G1355gat));
endmodule


