//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n462), .A2(new_n464), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  INV_X1    g050(.A(G113), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n468), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n467), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n465), .A2(new_n466), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n492), .A3(new_n466), .A4(new_n489), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n474), .A2(G138), .A3(new_n482), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(new_n482), .A3(new_n466), .A4(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n482), .B2(G114), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI211_X1 g082(.A(KEYINPUT70), .B(new_n500), .C1(new_n502), .C2(new_n504), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n497), .B(new_n499), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n494), .A2(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n511), .B1(new_n516), .B2(new_n515), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(KEYINPUT71), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(KEYINPUT71), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n514), .B1(new_n523), .B2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n518), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT5), .B(G543), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n517), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  INV_X1    g111(.A(G77), .ZN(new_n537));
  INV_X1    g112(.A(G543), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n531), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n541), .B1(new_n537), .B2(new_n538), .C1(new_n531), .C2(new_n536), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(G651), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n545));
  INV_X1    g120(.A(new_n518), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n515), .A2(new_n516), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n531), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT74), .B(G90), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n546), .A2(G52), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n544), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n545), .A2(new_n550), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(new_n554), .A3(new_n544), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  AND2_X1   g131(.A1(new_n511), .A2(G56), .ZN(new_n557));
  AND2_X1   g132(.A1(G68), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n546), .A2(G43), .B1(G81), .B2(new_n548), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n559), .A2(new_n560), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  AND3_X1   g145(.A1(new_n517), .A2(G91), .A3(new_n511), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(G65), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(G65), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n511), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G78), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n538), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n572), .B1(G651), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n546), .A2(G53), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  INV_X1    g158(.A(G168), .ZN(G286));
  AND2_X1   g159(.A1(new_n548), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n518), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n518), .A2(new_n591), .B1(new_n520), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n513), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n518), .A2(new_n598), .B1(new_n520), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n513), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(new_n548), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n531), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n546), .A2(G54), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g188(.A(new_n612), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n579), .A2(new_n581), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  OAI21_X1  g196(.A(G868), .B1(new_n611), .B2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g199(.A(new_n474), .ZN(new_n625));
  NOR3_X1   g200(.A1(new_n470), .A2(new_n625), .A3(G2105), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n626), .B(new_n627), .Z(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT13), .B(G2100), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n468), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n483), .A2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT80), .B(G2096), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(G14), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n651), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n671));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n668), .A2(new_n669), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT84), .ZN(new_n679));
  INV_X1    g254(.A(new_n670), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n673), .A2(new_n680), .A3(new_n677), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(G4), .A2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT89), .Z(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n611), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT91), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT90), .B(G1348), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(G20), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT23), .Z(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G299), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1956), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n483), .A2(G129), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT26), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n471), .A2(G105), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n468), .A2(G141), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n705), .B1(new_n715), .B2(new_n704), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT27), .B(G1996), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G19), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n565), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT92), .B(G1341), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n704), .B1(KEYINPUT24), .B2(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT24), .B2(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n479), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n720), .A2(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT94), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(KEYINPUT94), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n732), .A2(new_n733), .B1(new_n482), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n468), .A2(G139), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n704), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n704), .B2(G33), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n740), .A2(G2072), .B1(new_n720), .B2(new_n721), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n694), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n694), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n743), .A2(G1966), .B1(new_n704), .B2(new_n635), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G1966), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2072), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n744), .B(new_n752), .C1(new_n739), .C2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n727), .A2(new_n741), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n696), .A2(new_n697), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n468), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n483), .A2(G128), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n482), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n704), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2067), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n703), .A2(new_n755), .A3(new_n756), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n704), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n704), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT29), .Z(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n704), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n704), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n694), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n694), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n773), .B(new_n779), .C1(G1961), .C2(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n716), .A2(new_n717), .B1(new_n725), .B2(new_n724), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n781), .B2(G1961), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n768), .B(new_n782), .C1(KEYINPUT95), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(KEYINPUT95), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n694), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n694), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n788), .A2(KEYINPUT87), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(KEYINPUT87), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n789), .A2(new_n790), .A3(G1971), .ZN(new_n791));
  OAI21_X1  g366(.A(G1971), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n694), .A2(G23), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n589), .B2(new_n694), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT33), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1976), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n596), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT86), .Z(new_n801));
  NAND4_X1  g376(.A1(new_n791), .A2(new_n792), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n704), .A2(G25), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n468), .A2(G131), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n483), .A2(G119), .ZN(new_n807));
  OR2_X1    g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G107), .C2(new_n482), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n805), .B1(new_n811), .B2(new_n704), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT85), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT85), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n603), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G16), .B2(G24), .ZN(new_n818));
  INV_X1    g393(.A(G1986), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT88), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n815), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n803), .A2(new_n804), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n786), .A2(new_n825), .A3(new_n826), .ZN(G150));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n828));
  XNOR2_X1  g403(.A(G150), .B(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n619), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n518), .A2(new_n832), .B1(new_n520), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n513), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n565), .B(new_n837), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n831), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n837), .A2(new_n841), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(new_n479), .B(new_n635), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n487), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n468), .A2(G142), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n483), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n482), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n810), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n628), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n628), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n761), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n761), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n737), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n714), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n864));
  NAND2_X1  g439(.A1(G164), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n491), .A2(new_n493), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n505), .B(new_n506), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n499), .A4(new_n497), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT97), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n863), .A2(new_n870), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n861), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n859), .A3(new_n860), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n848), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n876), .A3(new_n848), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n616), .A2(new_n611), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n619), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n616), .B2(new_n611), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n611), .A2(new_n579), .A3(new_n891), .A4(new_n581), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G299), .B(new_n611), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(KEYINPUT100), .A3(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n890), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n611), .A2(G559), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n838), .B(new_n899), .Z(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n896), .B2(new_n900), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n589), .B(new_n603), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(G305), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n904), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n902), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G868), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g490(.A(new_n914), .B1(G868), .B2(new_n837), .ZN(G331));
  NAND3_X1  g491(.A1(new_n552), .A2(new_n555), .A3(G168), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G168), .B1(new_n552), .B2(new_n555), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n838), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(G171), .A2(G286), .ZN(new_n921));
  INV_X1    g496(.A(new_n838), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n923), .A3(KEYINPUT102), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(new_n922), .A3(new_n925), .A4(new_n917), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n924), .A2(new_n898), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n920), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(KEYINPUT103), .B(new_n838), .C1(new_n918), .C2(new_n919), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n896), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n911), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT104), .B1(new_n896), .B2(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n887), .A4(new_n893), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n888), .A2(new_n938), .A3(new_n889), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n940), .A2(new_n929), .A3(new_n930), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n896), .B1(new_n924), .B2(new_n926), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n911), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  OAI211_X1 g521(.A(KEYINPUT105), .B(new_n911), .C1(new_n941), .C2(new_n942), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n934), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n931), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n924), .A2(new_n898), .A3(new_n926), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n933), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n911), .B1(new_n927), .B2(new_n931), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n946), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n934), .A2(new_n945), .A3(new_n947), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(new_n946), .ZN(new_n959));
  MUX2_X1   g534(.A(new_n956), .B(new_n959), .S(KEYINPUT44), .Z(G397));
  INV_X1    g535(.A(KEYINPUT62), .ZN(new_n961));
  INV_X1    g536(.A(G1966), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n494), .B2(new_n509), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n963), .C1(new_n494), .C2(new_n509), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT45), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT106), .B(G40), .Z(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND4_X1   g545(.A1(new_n478), .A2(new_n469), .A3(new_n472), .A4(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n964), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n962), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n965), .A2(new_n975), .A3(new_n967), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n473), .A2(new_n478), .A3(new_n970), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G2084), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT110), .B(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(G168), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT120), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n987));
  INV_X1    g562(.A(new_n967), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n966), .B1(new_n868), .B2(new_n963), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n972), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n973), .ZN(new_n991));
  AOI21_X1  g566(.A(G1966), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n993));
  OAI21_X1  g568(.A(G8), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT121), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n983), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n981), .A2(KEYINPUT121), .A3(G8), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n982), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT51), .B(new_n983), .C1(new_n981), .C2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n961), .B(new_n986), .C1(new_n998), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT124), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n976), .A2(new_n971), .A3(new_n977), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1961), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n976), .A2(KEYINPUT115), .A3(new_n971), .A4(new_n977), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n978), .B1(new_n972), .B2(new_n964), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n865), .A2(new_n869), .A3(KEYINPUT45), .A4(new_n963), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2078), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1008), .B1(KEYINPUT53), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n968), .A2(new_n973), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(new_n777), .ZN(new_n1016));
  NOR4_X1   g591(.A1(new_n968), .A2(new_n973), .A3(KEYINPUT122), .A4(G2078), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(G171), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n868), .A2(new_n975), .A3(new_n963), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT50), .B1(new_n988), .B2(new_n989), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n772), .A3(new_n1024), .A4(new_n971), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT107), .B(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1011), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n982), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT109), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  MUX2_X1   g607(.A(new_n1030), .B(new_n1031), .S(new_n1032), .Z(new_n1033));
  NOR2_X1   g608(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1027), .B1(G2090), .B2(new_n1003), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(G8), .A3(new_n1033), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n965), .A2(new_n971), .A3(new_n967), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n589), .A2(G1976), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n999), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n596), .B2(new_n1042), .ZN(new_n1043));
  NOR4_X1   g618(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT111), .A4(G1981), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1043), .A2(new_n1044), .B1(new_n1042), .B2(new_n596), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT112), .ZN(new_n1049));
  OAI221_X1 g624(.A(new_n1049), .B1(new_n1042), .B2(new_n596), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1047), .A2(new_n999), .A3(new_n1050), .A4(new_n1037), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1037), .A2(new_n999), .A3(new_n1038), .A4(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1040), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1036), .A2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1020), .A2(new_n1034), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1001), .A2(new_n1002), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n986), .B1(new_n998), .B2(new_n1000), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1002), .B1(new_n1001), .B2(new_n1057), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT125), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1001), .A2(new_n1057), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT124), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1060), .A4(new_n1058), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1051), .A2(new_n1052), .A3(new_n589), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1037), .A2(new_n999), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1069), .B2(KEYINPUT113), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1036), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1070), .A2(new_n1072), .B1(new_n1073), .B2(new_n1055), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1056), .A2(new_n1034), .ZN(new_n1075));
  AOI211_X1 g650(.A(G286), .B(new_n982), .C1(new_n974), .C2(new_n980), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT63), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1033), .B1(new_n1035), .B2(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(KEYINPUT63), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1056), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n616), .B(KEYINPUT57), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1023), .A2(new_n971), .A3(new_n1024), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1082), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1085), .A2(new_n1082), .A3(new_n1088), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n611), .ZN(new_n1091));
  INV_X1    g666(.A(G1348), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1005), .A2(new_n1092), .A3(new_n1007), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1037), .A2(G2067), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1089), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND3_X1  g673(.A1(new_n1037), .A2(KEYINPUT116), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1011), .B2(G1996), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT116), .B1(new_n1037), .B2(new_n1098), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(new_n565), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n1094), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1104), .A2(new_n619), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1090), .A2(new_n1089), .A3(KEYINPUT118), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1082), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(KEYINPUT118), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1103), .B(new_n1105), .C1(new_n1106), .C2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1082), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1089), .B2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n1082), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1095), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(new_n1104), .A3(new_n619), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1096), .B1(new_n1112), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1124));
  OR2_X1    g699(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(new_n1125), .C1(new_n1013), .C2(new_n1019), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n870), .A2(new_n963), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n972), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n482), .B1(new_n477), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1129), .B2(new_n477), .ZN(new_n1131));
  AND4_X1   g706(.A1(KEYINPUT53), .A2(new_n473), .A3(G40), .A4(new_n777), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1133), .A2(new_n1010), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1134), .B(new_n1008), .C1(KEYINPUT53), .C2(new_n1012), .ZN(new_n1135));
  AND4_X1   g710(.A1(new_n1059), .A2(new_n1126), .A3(new_n1075), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1081), .B1(new_n1123), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1063), .A2(new_n1067), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1128), .A2(new_n978), .ZN(new_n1139));
  INV_X1    g714(.A(G1996), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n714), .B(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n761), .B(G2067), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n811), .A2(new_n813), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n811), .A2(new_n813), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n603), .B(new_n819), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1139), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT46), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1142), .A2(new_n715), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1149), .A2(new_n1150), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1153), .A2(KEYINPUT126), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(KEYINPUT126), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT47), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1158), .A2(new_n1143), .B1(G2067), .B2(new_n761), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1139), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1139), .A2(new_n819), .A3(new_n603), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT48), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1160), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1157), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1148), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  NOR2_X1   g744(.A1(G227), .A2(new_n459), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1171), .B1(new_n688), .B2(new_n689), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1172), .A2(G401), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1173), .A2(new_n883), .ZN(new_n1174));
  AOI211_X1 g748(.A(new_n1170), .B(new_n1174), .C1(new_n948), .C2(new_n955), .ZN(new_n1175));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1176));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n956), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1177), .ZN(G308));
  NAND2_X1  g752(.A1(new_n956), .A2(new_n1176), .ZN(G225));
endmodule


