

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n649, n650, n651, n652, n653, n654, n655, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759;

  AND2_X1 U360 ( .A1(n338), .A2(n337), .ZN(n649) );
  AND2_X1 U361 ( .A1(n341), .A2(n340), .ZN(n657) );
  INV_X1 U362 ( .A(n723), .ZN(n337) );
  INV_X1 U363 ( .A(n723), .ZN(n340) );
  XNOR2_X1 U364 ( .A(n647), .B(n339), .ZN(n338) );
  XNOR2_X1 U365 ( .A(n655), .B(n342), .ZN(n341) );
  BUF_X1 U366 ( .A(n673), .Z(n343) );
  XNOR2_X1 U367 ( .A(n550), .B(n549), .ZN(n673) );
  XNOR2_X1 U368 ( .A(n602), .B(KEYINPUT1), .ZN(n539) );
  INV_X1 U369 ( .A(G143), .ZN(n450) );
  INV_X1 U370 ( .A(n646), .ZN(n339) );
  INV_X1 U371 ( .A(n654), .ZN(n342) );
  XNOR2_X1 U372 ( .A(n404), .B(KEYINPUT4), .ZN(n501) );
  XOR2_X1 U373 ( .A(n501), .B(n726), .Z(n516) );
  XNOR2_X1 U374 ( .A(n420), .B(KEYINPUT19), .ZN(n396) );
  XNOR2_X1 U375 ( .A(n456), .B(KEYINPUT73), .ZN(n726) );
  BUF_X1 U376 ( .A(G143), .Z(n346) );
  AND2_X2 U377 ( .A1(n401), .A2(n402), .ZN(n362) );
  XNOR2_X2 U378 ( .A(n444), .B(n443), .ZN(n706) );
  INV_X4 U379 ( .A(G116), .ZN(n426) );
  AND2_X1 U380 ( .A1(n435), .A2(n433), .ZN(n432) );
  OR2_X1 U381 ( .A1(n546), .A2(n675), .ZN(n418) );
  NOR2_X1 U382 ( .A1(n608), .A2(n600), .ZN(n597) );
  AND2_X1 U383 ( .A1(n375), .A2(n374), .ZN(n575) );
  NOR2_X1 U384 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U385 ( .A(n534), .B(n533), .ZN(n574) );
  XNOR2_X1 U386 ( .A(n652), .B(n653), .ZN(n654) );
  XNOR2_X1 U387 ( .A(n645), .B(KEYINPUT59), .ZN(n646) );
  XNOR2_X1 U388 ( .A(n484), .B(n425), .ZN(n424) );
  XNOR2_X1 U389 ( .A(n423), .B(G104), .ZN(n475) );
  XNOR2_X1 U390 ( .A(G122), .B(G113), .ZN(n423) );
  XNOR2_X1 U391 ( .A(G146), .B(G125), .ZN(n471) );
  XNOR2_X1 U392 ( .A(G101), .B(KEYINPUT68), .ZN(n404) );
  XNOR2_X1 U393 ( .A(G119), .B(KEYINPUT3), .ZN(n456) );
  XNOR2_X1 U394 ( .A(KEYINPUT16), .B(G110), .ZN(n425) );
  XNOR2_X1 U395 ( .A(n344), .B(n345), .ZN(n580) );
  NOR2_X1 U396 ( .A1(n651), .A2(n622), .ZN(n344) );
  NAND2_X1 U397 ( .A1(n460), .A2(G210), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n424), .B(n475), .ZN(n725) );
  BUF_X1 U399 ( .A(n391), .Z(n347) );
  BUF_X1 U400 ( .A(n624), .Z(n348) );
  XNOR2_X2 U401 ( .A(n499), .B(n422), .ZN(n551) );
  NAND2_X1 U402 ( .A1(n387), .A2(n388), .ZN(n415) );
  NOR2_X1 U403 ( .A1(n675), .A2(n389), .ZN(n388) );
  INV_X1 U404 ( .A(KEYINPUT104), .ZN(n389) );
  NOR2_X1 U405 ( .A1(n380), .A2(n378), .ZN(n437) );
  AND2_X1 U406 ( .A1(n379), .A2(n438), .ZN(n378) );
  NAND2_X1 U407 ( .A1(n383), .A2(n381), .ZN(n380) );
  NOR2_X1 U408 ( .A1(n440), .A2(n439), .ZN(n438) );
  XNOR2_X1 U409 ( .A(n471), .B(KEYINPUT10), .ZN(n521) );
  AND2_X1 U410 ( .A1(n354), .A2(n384), .ZN(n383) );
  INV_X1 U411 ( .A(n701), .ZN(n370) );
  INV_X1 U412 ( .A(KEYINPUT85), .ZN(n411) );
  NOR2_X1 U413 ( .A1(n573), .A2(n572), .ZN(n589) );
  XNOR2_X1 U414 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n594) );
  XNOR2_X1 U415 ( .A(n521), .B(n520), .ZN(n740) );
  XNOR2_X1 U416 ( .A(n487), .B(G122), .ZN(n429) );
  XNOR2_X1 U417 ( .A(n518), .B(n508), .ZN(n624) );
  XNOR2_X1 U418 ( .A(n405), .B(n501), .ZN(n505) );
  NAND2_X1 U419 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U420 ( .A(n462), .B(n463), .ZN(n464) );
  XNOR2_X1 U421 ( .A(n461), .B(KEYINPUT75), .ZN(n462) );
  XOR2_X1 U422 ( .A(KEYINPUT90), .B(KEYINPUT14), .Z(n463) );
  NAND2_X1 U423 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U424 ( .A(n532), .B(KEYINPUT25), .ZN(n533) );
  XNOR2_X1 U425 ( .A(n445), .B(KEYINPUT28), .ZN(n603) );
  NOR2_X1 U426 ( .A1(n584), .A2(n585), .ZN(n445) );
  INV_X1 U427 ( .A(KEYINPUT92), .ZN(n422) );
  INV_X1 U428 ( .A(n577), .ZN(n393) );
  INV_X1 U429 ( .A(KEYINPUT22), .ZN(n410) );
  XNOR2_X1 U430 ( .A(KEYINPUT89), .B(KEYINPUT15), .ZN(n458) );
  INV_X1 U431 ( .A(G237), .ZN(n459) );
  INV_X1 U432 ( .A(G902), .ZN(n479) );
  XNOR2_X1 U433 ( .A(G137), .B(G113), .ZN(n511) );
  XOR2_X1 U434 ( .A(KEYINPUT5), .B(G116), .Z(n512) );
  XNOR2_X1 U435 ( .A(n408), .B(G140), .ZN(n519) );
  INV_X1 U436 ( .A(G137), .ZN(n408) );
  XOR2_X1 U437 ( .A(KEYINPUT74), .B(KEYINPUT93), .Z(n523) );
  XNOR2_X1 U438 ( .A(G128), .B(KEYINPUT24), .ZN(n522) );
  XNOR2_X1 U439 ( .A(G119), .B(G110), .ZN(n525) );
  NOR2_X1 U440 ( .A1(G953), .A2(G237), .ZN(n513) );
  XOR2_X1 U441 ( .A(KEYINPUT70), .B(G131), .Z(n507) );
  XNOR2_X1 U442 ( .A(n519), .B(n406), .ZN(n405) );
  XNOR2_X1 U443 ( .A(n407), .B(G110), .ZN(n406) );
  INV_X1 U444 ( .A(G104), .ZN(n407) );
  INV_X1 U445 ( .A(G107), .ZN(n502) );
  XNOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n452) );
  INV_X1 U447 ( .A(KEYINPUT48), .ZN(n441) );
  NAND2_X1 U448 ( .A1(n353), .A2(n360), .ZN(n400) );
  AND2_X1 U449 ( .A1(n751), .A2(G952), .ZN(n386) );
  OR2_X1 U450 ( .A1(n575), .A2(KEYINPUT71), .ZN(n373) );
  XOR2_X1 U451 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n552) );
  XNOR2_X1 U452 ( .A(n595), .B(n594), .ZN(n596) );
  BUF_X1 U453 ( .A(n580), .Z(n609) );
  OR2_X1 U454 ( .A1(n555), .A2(n545), .ZN(n641) );
  INV_X1 U455 ( .A(n619), .ZN(n748) );
  XNOR2_X1 U456 ( .A(n447), .B(n446), .ZN(n720) );
  XNOR2_X1 U457 ( .A(n528), .B(n530), .ZN(n447) );
  INV_X1 U458 ( .A(n740), .ZN(n446) );
  XNOR2_X1 U459 ( .A(n428), .B(n427), .ZN(n716) );
  XNOR2_X1 U460 ( .A(n506), .B(n490), .ZN(n427) );
  XNOR2_X1 U461 ( .A(n486), .B(n429), .ZN(n428) );
  INV_X1 U462 ( .A(KEYINPUT2), .ZN(n620) );
  NAND2_X1 U463 ( .A1(n464), .A2(G952), .ZN(n688) );
  NOR2_X1 U464 ( .A1(n421), .A2(n669), .ZN(n542) );
  INV_X1 U465 ( .A(KEYINPUT80), .ZN(n443) );
  AND2_X1 U466 ( .A1(n398), .A2(n591), .ZN(n701) );
  XNOR2_X1 U467 ( .A(n371), .B(KEYINPUT67), .ZN(n398) );
  NOR2_X1 U468 ( .A1(n593), .A2(n660), .ZN(n372) );
  INV_X1 U469 ( .A(KEYINPUT95), .ZN(n358) );
  XNOR2_X1 U470 ( .A(n394), .B(KEYINPUT84), .ZN(n535) );
  XNOR2_X1 U471 ( .A(n628), .B(n627), .ZN(n630) );
  INV_X1 U472 ( .A(G122), .ZN(n390) );
  OR2_X1 U473 ( .A1(n571), .A2(n466), .ZN(n349) );
  AND2_X1 U474 ( .A1(n660), .A2(n561), .ZN(n350) );
  AND2_X1 U475 ( .A1(n415), .A2(n411), .ZN(n351) );
  AND2_X1 U476 ( .A1(n431), .A2(n437), .ZN(n352) );
  AND2_X1 U477 ( .A1(n416), .A2(n351), .ZN(n353) );
  OR2_X1 U478 ( .A1(n640), .A2(KEYINPUT81), .ZN(n354) );
  AND2_X1 U479 ( .A1(n587), .A2(n376), .ZN(n355) );
  INV_X2 U480 ( .A(G953), .ZN(n751) );
  XNOR2_X1 U481 ( .A(KEYINPUT87), .B(KEYINPUT0), .ZN(n356) );
  XOR2_X1 U482 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n357) );
  INV_X1 U483 ( .A(KEYINPUT81), .ZN(n439) );
  BUF_X1 U484 ( .A(n650), .Z(n719) );
  XNOR2_X1 U485 ( .A(n359), .B(n358), .ZN(n697) );
  NOR2_X1 U486 ( .A1(n551), .A2(n538), .ZN(n359) );
  AND2_X1 U487 ( .A1(n560), .A2(n414), .ZN(n360) );
  NAND2_X1 U488 ( .A1(n560), .A2(n414), .ZN(n413) );
  NAND2_X1 U489 ( .A1(n413), .A2(KEYINPUT85), .ZN(n401) );
  NAND2_X1 U490 ( .A1(n361), .A2(n596), .ZN(n608) );
  XNOR2_X1 U491 ( .A(n592), .B(KEYINPUT76), .ZN(n361) );
  NAND2_X1 U492 ( .A1(n362), .A2(n400), .ZN(n399) );
  AND2_X1 U493 ( .A1(n363), .A2(n366), .ZN(n403) );
  NAND2_X1 U494 ( .A1(n364), .A2(KEYINPUT44), .ZN(n363) );
  NOR2_X1 U495 ( .A1(n757), .A2(KEYINPUT69), .ZN(n365) );
  INV_X1 U496 ( .A(n757), .ZN(n369) );
  NAND2_X1 U497 ( .A1(n365), .A2(n370), .ZN(n364) );
  NAND2_X1 U498 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U499 ( .A1(n397), .A2(n367), .ZN(n366) );
  NOR2_X1 U500 ( .A1(n368), .A2(KEYINPUT44), .ZN(n367) );
  NAND2_X1 U501 ( .A1(n409), .A2(n372), .ZN(n371) );
  XNOR2_X2 U502 ( .A(n500), .B(n410), .ZN(n409) );
  NAND2_X1 U503 ( .A1(n576), .A2(n373), .ZN(n584) );
  XNOR2_X1 U504 ( .A(n589), .B(KEYINPUT72), .ZN(n374) );
  INV_X1 U505 ( .A(n574), .ZN(n375) );
  NAND2_X1 U506 ( .A1(n706), .A2(n587), .ZN(n382) );
  NAND2_X1 U507 ( .A1(n706), .A2(n355), .ZN(n384) );
  INV_X1 U508 ( .A(KEYINPUT47), .ZN(n376) );
  NAND2_X1 U509 ( .A1(n382), .A2(KEYINPUT47), .ZN(n379) );
  NAND2_X1 U510 ( .A1(n382), .A2(n377), .ZN(n381) );
  AND2_X1 U511 ( .A1(n439), .A2(KEYINPUT47), .ZN(n377) );
  NAND2_X1 U512 ( .A1(n464), .A2(n386), .ZN(n385) );
  XNOR2_X1 U513 ( .A(n385), .B(KEYINPUT91), .ZN(n571) );
  XNOR2_X2 U514 ( .A(n419), .B(n356), .ZN(n499) );
  INV_X1 U515 ( .A(n546), .ZN(n387) );
  NAND2_X1 U516 ( .A1(n391), .A2(KEYINPUT44), .ZN(n560) );
  XNOR2_X1 U517 ( .A(n347), .B(n390), .ZN(G24) );
  XNOR2_X1 U518 ( .A(n391), .B(KEYINPUT69), .ZN(n397) );
  XNOR2_X2 U519 ( .A(n559), .B(n558), .ZN(n391) );
  NAND2_X1 U520 ( .A1(n409), .A2(n392), .ZN(n394) );
  NOR2_X1 U521 ( .A1(n660), .A2(n393), .ZN(n392) );
  XNOR2_X1 U522 ( .A(n395), .B(n357), .ZN(n731) );
  NAND2_X1 U523 ( .A1(n399), .A2(n403), .ZN(n395) );
  XNOR2_X2 U524 ( .A(n666), .B(KEYINPUT6), .ZN(n577) );
  NAND2_X1 U525 ( .A1(n396), .A2(n349), .ZN(n419) );
  AND2_X1 U526 ( .A1(n396), .A2(n602), .ZN(n586) );
  NAND2_X1 U527 ( .A1(n412), .A2(KEYINPUT85), .ZN(n402) );
  XNOR2_X2 U528 ( .A(n741), .B(G146), .ZN(n518) );
  XNOR2_X2 U529 ( .A(n506), .B(n507), .ZN(n741) );
  XNOR2_X2 U530 ( .A(n485), .B(G134), .ZN(n506) );
  NOR2_X1 U531 ( .A1(n756), .A2(n759), .ZN(n606) );
  XNOR2_X1 U532 ( .A(n606), .B(KEYINPUT46), .ZN(n442) );
  NOR2_X2 U533 ( .A1(n547), .A2(n577), .ZN(n550) );
  NAND2_X1 U534 ( .A1(n539), .A2(n659), .ZN(n547) );
  XNOR2_X2 U535 ( .A(n450), .B(G128), .ZN(n485) );
  NAND2_X1 U536 ( .A1(n416), .A2(n415), .ZN(n412) );
  NAND2_X1 U537 ( .A1(n417), .A2(n418), .ZN(n416) );
  NAND2_X1 U538 ( .A1(n350), .A2(n409), .ZN(n562) );
  NAND2_X1 U539 ( .A1(n644), .A2(KEYINPUT104), .ZN(n414) );
  NOR2_X1 U540 ( .A1(n644), .A2(KEYINPUT104), .ZN(n417) );
  NAND2_X1 U541 ( .A1(n580), .A2(n677), .ZN(n420) );
  INV_X1 U542 ( .A(n499), .ZN(n421) );
  XNOR2_X2 U543 ( .A(n426), .B(G107), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n505), .B(n504), .ZN(n508) );
  NAND2_X1 U545 ( .A1(n432), .A2(n430), .ZN(n618) );
  NAND2_X1 U546 ( .A1(n352), .A2(n442), .ZN(n430) );
  AND2_X1 U547 ( .A1(n588), .A2(KEYINPUT48), .ZN(n431) );
  NAND2_X1 U548 ( .A1(n434), .A2(n441), .ZN(n433) );
  NAND2_X1 U549 ( .A1(n437), .A2(n588), .ZN(n434) );
  NAND2_X1 U550 ( .A1(n436), .A2(n441), .ZN(n435) );
  INV_X1 U551 ( .A(n442), .ZN(n436) );
  INV_X1 U552 ( .A(n640), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n603), .A2(n586), .ZN(n444) );
  NOR2_X1 U554 ( .A1(n697), .A2(n712), .ZN(n546) );
  AND2_X1 U555 ( .A1(n513), .A2(G210), .ZN(n448) );
  AND2_X1 U556 ( .A1(n630), .A2(n636), .ZN(G54) );
  XNOR2_X1 U557 ( .A(n514), .B(n448), .ZN(n515) );
  XNOR2_X1 U558 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U559 ( .A(n516), .B(n515), .ZN(n517) );
  INV_X1 U560 ( .A(KEYINPUT23), .ZN(n524) );
  XNOR2_X1 U561 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U562 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U563 ( .A(n568), .B(n567), .ZN(n593) );
  XNOR2_X1 U564 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n581) );
  XNOR2_X1 U565 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U566 ( .A(n723), .ZN(n636) );
  INV_X1 U567 ( .A(KEYINPUT35), .ZN(n558) );
  XNOR2_X1 U568 ( .A(n485), .B(n471), .ZN(n454) );
  NAND2_X1 U569 ( .A1(n751), .A2(G224), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U571 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U572 ( .A(n725), .B(n455), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n457), .B(n516), .ZN(n651) );
  XNOR2_X1 U574 ( .A(n458), .B(n479), .ZN(n493) );
  INV_X1 U575 ( .A(n493), .ZN(n622) );
  NAND2_X1 U576 ( .A1(n479), .A2(n459), .ZN(n460) );
  NAND2_X1 U577 ( .A1(n460), .A2(G214), .ZN(n677) );
  AND2_X1 U578 ( .A1(n464), .A2(G953), .ZN(n465) );
  NAND2_X1 U579 ( .A1(G902), .A2(n465), .ZN(n569) );
  NOR2_X1 U580 ( .A1(n569), .A2(G898), .ZN(n466) );
  XNOR2_X1 U581 ( .A(n507), .B(n346), .ZN(n470) );
  XOR2_X1 U582 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n468) );
  XNOR2_X1 U583 ( .A(G140), .B(KEYINPUT11), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U585 ( .A(n470), .B(n469), .ZN(n473) );
  INV_X1 U586 ( .A(n521), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n473), .B(n472), .ZN(n478) );
  NAND2_X1 U588 ( .A1(G214), .A2(n513), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n474), .B(KEYINPUT12), .ZN(n476) );
  XNOR2_X1 U590 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U591 ( .A(n478), .B(n477), .ZN(n645) );
  NAND2_X1 U592 ( .A1(n645), .A2(n479), .ZN(n481) );
  XNOR2_X1 U593 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n481), .B(n480), .ZN(n555) );
  XNOR2_X1 U595 ( .A(KEYINPUT102), .B(G478), .ZN(n492) );
  XOR2_X1 U596 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n483) );
  XNOR2_X1 U597 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n482) );
  XNOR2_X1 U598 ( .A(n483), .B(n482), .ZN(n487) );
  XOR2_X1 U599 ( .A(KEYINPUT101), .B(n484), .Z(n486) );
  XOR2_X1 U600 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n489) );
  NAND2_X1 U601 ( .A1(G234), .A2(n751), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n489), .B(n488), .ZN(n529) );
  NAND2_X1 U603 ( .A1(G217), .A2(n529), .ZN(n490) );
  NOR2_X1 U604 ( .A1(G902), .A2(n716), .ZN(n491) );
  XNOR2_X1 U605 ( .A(n492), .B(n491), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n680) );
  NAND2_X1 U607 ( .A1(n493), .A2(G234), .ZN(n495) );
  XNOR2_X1 U608 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n531) );
  NAND2_X1 U610 ( .A1(n531), .A2(G221), .ZN(n497) );
  INV_X1 U611 ( .A(KEYINPUT21), .ZN(n496) );
  XNOR2_X1 U612 ( .A(n497), .B(n496), .ZN(n663) );
  INV_X1 U613 ( .A(n663), .ZN(n573) );
  NOR2_X1 U614 ( .A1(n680), .A2(n573), .ZN(n498) );
  NAND2_X1 U615 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND2_X1 U616 ( .A1(G227), .A2(n751), .ZN(n503) );
  NOR2_X1 U617 ( .A1(n624), .A2(G902), .ZN(n510) );
  INV_X1 U618 ( .A(G469), .ZN(n509) );
  XNOR2_X2 U619 ( .A(n510), .B(n509), .ZN(n602) );
  BUF_X1 U620 ( .A(n539), .Z(n660) );
  XNOR2_X1 U621 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U622 ( .A(n518), .B(n517), .ZN(n632) );
  NOR2_X2 U623 ( .A1(n632), .A2(G902), .ZN(n568) );
  INV_X1 U624 ( .A(G472), .ZN(n566) );
  XNOR2_X2 U625 ( .A(n568), .B(n566), .ZN(n666) );
  INV_X1 U626 ( .A(n519), .ZN(n520) );
  XNOR2_X1 U627 ( .A(n523), .B(n522), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U629 ( .A1(n529), .A2(G221), .ZN(n530) );
  NOR2_X1 U630 ( .A1(n720), .A2(G902), .ZN(n534) );
  NAND2_X1 U631 ( .A1(n531), .A2(G217), .ZN(n532) );
  INV_X1 U632 ( .A(n574), .ZN(n591) );
  NOR2_X2 U633 ( .A1(n535), .A2(n591), .ZN(n644) );
  AND2_X1 U634 ( .A1(n574), .A2(n663), .ZN(n659) );
  INV_X1 U635 ( .A(n659), .ZN(n536) );
  NOR2_X1 U636 ( .A1(n666), .A2(n536), .ZN(n537) );
  NAND2_X1 U637 ( .A1(n602), .A2(n537), .ZN(n538) );
  INV_X1 U638 ( .A(n547), .ZN(n540) );
  NAND2_X1 U639 ( .A1(n666), .A2(n540), .ZN(n669) );
  XOR2_X1 U640 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n541) );
  XNOR2_X1 U641 ( .A(n542), .B(n541), .ZN(n712) );
  INV_X1 U642 ( .A(n554), .ZN(n545) );
  NAND2_X1 U643 ( .A1(n555), .A2(n545), .ZN(n544) );
  INV_X1 U644 ( .A(KEYINPUT103), .ZN(n543) );
  XNOR2_X1 U645 ( .A(n544), .B(n543), .ZN(n696) );
  NAND2_X1 U646 ( .A1(n696), .A2(n641), .ZN(n587) );
  INV_X1 U647 ( .A(n587), .ZN(n675) );
  XNOR2_X1 U648 ( .A(KEYINPUT33), .B(KEYINPUT88), .ZN(n548) );
  XNOR2_X1 U649 ( .A(n548), .B(KEYINPUT106), .ZN(n549) );
  NOR2_X1 U650 ( .A1(n673), .A2(n551), .ZN(n553) );
  XNOR2_X1 U651 ( .A(n553), .B(n552), .ZN(n557) );
  OR2_X1 U652 ( .A1(n555), .A2(n554), .ZN(n607) );
  XOR2_X1 U653 ( .A(n607), .B(KEYINPUT77), .Z(n556) );
  NOR2_X2 U654 ( .A1(n557), .A2(n556), .ZN(n559) );
  XOR2_X1 U655 ( .A(KEYINPUT79), .B(n577), .Z(n561) );
  NOR2_X1 U656 ( .A1(n574), .A2(n562), .ZN(n564) );
  XNOR2_X1 U657 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n563) );
  XNOR2_X1 U658 ( .A(n564), .B(n563), .ZN(n757) );
  INV_X1 U659 ( .A(KEYINPUT105), .ZN(n565) );
  INV_X1 U660 ( .A(n593), .ZN(n585) );
  NOR2_X1 U661 ( .A1(G900), .A2(n569), .ZN(n570) );
  NOR2_X1 U662 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U663 ( .A1(KEYINPUT71), .A2(n575), .ZN(n576) );
  OR2_X1 U664 ( .A1(n584), .A2(n577), .ZN(n578) );
  NOR2_X1 U665 ( .A1(n578), .A2(n641), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n579), .A2(n677), .ZN(n613) );
  INV_X1 U667 ( .A(n609), .ZN(n615) );
  NOR2_X1 U668 ( .A1(n613), .A2(n615), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n583), .A2(n660), .ZN(n714) );
  XOR2_X1 U670 ( .A(n714), .B(KEYINPUT83), .Z(n588) );
  NAND2_X1 U671 ( .A1(n589), .A2(n602), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n593), .A2(n677), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n609), .B(KEYINPUT38), .ZN(n600) );
  XNOR2_X1 U674 ( .A(KEYINPUT39), .B(n597), .ZN(n611) );
  NOR2_X1 U675 ( .A1(n611), .A2(n641), .ZN(n599) );
  XNOR2_X1 U676 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n599), .B(n598), .ZN(n756) );
  INV_X1 U678 ( .A(n600), .ZN(n678) );
  NAND2_X1 U679 ( .A1(n678), .A2(n677), .ZN(n674) );
  NOR2_X1 U680 ( .A1(n680), .A2(n674), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT41), .ZN(n689) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n689), .A2(n604), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT42), .ZN(n759) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n640) );
  NOR2_X1 U687 ( .A1(n696), .A2(n611), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT109), .ZN(n755) );
  NOR2_X1 U689 ( .A1(n660), .A2(n613), .ZN(n614) );
  XOR2_X1 U690 ( .A(n614), .B(KEYINPUT43), .Z(n616) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n643) );
  AND2_X1 U692 ( .A1(n755), .A2(n643), .ZN(n617) );
  NOR2_X2 U693 ( .A1(n731), .A2(n619), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n658) );
  NAND2_X1 U695 ( .A1(n658), .A2(n622), .ZN(n623) );
  XNOR2_X2 U696 ( .A(n623), .B(KEYINPUT65), .ZN(n650) );
  NAND2_X1 U697 ( .A1(n719), .A2(G469), .ZN(n628) );
  XOR2_X1 U698 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n626) );
  XNOR2_X1 U699 ( .A(n348), .B(KEYINPUT117), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  INV_X1 U701 ( .A(G952), .ZN(n629) );
  AND2_X1 U702 ( .A1(n629), .A2(G953), .ZN(n723) );
  NAND2_X1 U703 ( .A1(n650), .A2(G472), .ZN(n634) );
  XNOR2_X1 U704 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n635) );
  INV_X1 U707 ( .A(n635), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U710 ( .A(n346), .B(KEYINPUT113), .Z(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(G45) );
  INV_X1 U712 ( .A(n641), .ZN(n709) );
  NAND2_X1 U713 ( .A1(n697), .A2(n709), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(G104), .ZN(G6) );
  XNOR2_X1 U715 ( .A(n643), .B(G140), .ZN(G42) );
  XOR2_X1 U716 ( .A(n644), .B(G101), .Z(G3) );
  NAND2_X1 U717 ( .A1(n650), .A2(G475), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n649), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n650), .A2(G210), .ZN(n655) );
  BUF_X1 U720 ( .A(n651), .Z(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n653) );
  XNOR2_X1 U722 ( .A(n657), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U723 ( .A(n658), .Z(n694) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U725 ( .A(n661), .B(KEYINPUT115), .ZN(n662) );
  XNOR2_X1 U726 ( .A(n662), .B(KEYINPUT50), .ZN(n668) );
  NOR2_X1 U727 ( .A1(n663), .A2(n574), .ZN(n664) );
  XOR2_X1 U728 ( .A(KEYINPUT49), .B(n664), .Z(n665) );
  NOR2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U732 ( .A(KEYINPUT51), .B(n671), .ZN(n672) );
  NOR2_X1 U733 ( .A1(n689), .A2(n672), .ZN(n685) );
  NOR2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U735 ( .A(KEYINPUT116), .B(n676), .ZN(n682) );
  NOR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U737 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U738 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U739 ( .A1(n343), .A2(n683), .ZN(n684) );
  NOR2_X1 U740 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n686), .B(KEYINPUT52), .ZN(n687) );
  NOR2_X1 U742 ( .A1(n688), .A2(n687), .ZN(n691) );
  NOR2_X1 U743 ( .A1(n343), .A2(n689), .ZN(n690) );
  NOR2_X1 U744 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U745 ( .A1(n692), .A2(n751), .ZN(n693) );
  NOR2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U747 ( .A(n695), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U748 ( .A(n696), .ZN(n711) );
  NAND2_X1 U749 ( .A1(n697), .A2(n711), .ZN(n699) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n698) );
  XNOR2_X1 U751 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U752 ( .A(G107), .B(n700), .ZN(G9) );
  XOR2_X1 U753 ( .A(G110), .B(n701), .Z(G12) );
  XOR2_X1 U754 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n703) );
  NAND2_X1 U755 ( .A1(n711), .A2(n706), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n705) );
  XOR2_X1 U757 ( .A(G128), .B(KEYINPUT111), .Z(n704) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(G30) );
  NAND2_X1 U759 ( .A1(n706), .A2(n709), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT114), .ZN(n708) );
  XNOR2_X1 U761 ( .A(G146), .B(n708), .ZN(G48) );
  NAND2_X1 U762 ( .A1(n712), .A2(n709), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n710), .B(G113), .ZN(G15) );
  NAND2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(G116), .ZN(G18) );
  XOR2_X1 U766 ( .A(G125), .B(KEYINPUT37), .Z(n715) );
  XNOR2_X1 U767 ( .A(n714), .B(n715), .ZN(G27) );
  NAND2_X1 U768 ( .A1(n719), .A2(G478), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U770 ( .A1(n723), .A2(n718), .ZN(G63) );
  NAND2_X1 U771 ( .A1(n719), .A2(G217), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(G66) );
  XOR2_X1 U774 ( .A(G101), .B(KEYINPUT121), .Z(n724) );
  XNOR2_X1 U775 ( .A(n725), .B(n724), .ZN(n727) );
  XNOR2_X1 U776 ( .A(n726), .B(n727), .ZN(n729) );
  NOR2_X1 U777 ( .A1(n751), .A2(G898), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(KEYINPUT120), .B(n730), .ZN(n739) );
  OR2_X1 U780 ( .A1(n731), .A2(G953), .ZN(n737) );
  XOR2_X1 U781 ( .A(KEYINPUT61), .B(KEYINPUT119), .Z(n733) );
  NAND2_X1 U782 ( .A1(G224), .A2(G953), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(KEYINPUT118), .B(n734), .ZN(n735) );
  NAND2_X1 U785 ( .A1(n735), .A2(G898), .ZN(n736) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(G69) );
  XOR2_X1 U788 ( .A(KEYINPUT122), .B(n740), .Z(n743) );
  XNOR2_X1 U789 ( .A(n741), .B(KEYINPUT4), .ZN(n742) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(n749) );
  XNOR2_X1 U791 ( .A(G227), .B(n749), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(KEYINPUT124), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  XOR2_X1 U794 ( .A(KEYINPUT125), .B(n746), .Z(n747) );
  NAND2_X1 U795 ( .A1(G953), .A2(n747), .ZN(n754) );
  XNOR2_X1 U796 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n750), .B(KEYINPUT123), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n754), .A2(n753), .ZN(G72) );
  XNOR2_X1 U800 ( .A(G134), .B(n755), .ZN(G36) );
  XOR2_X1 U801 ( .A(n756), .B(G131), .Z(G33) );
  XOR2_X1 U802 ( .A(G119), .B(n757), .Z(n758) );
  XNOR2_X1 U803 ( .A(KEYINPUT126), .B(n758), .ZN(G21) );
  XOR2_X1 U804 ( .A(G137), .B(n759), .Z(G39) );
endmodule

