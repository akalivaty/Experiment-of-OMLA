

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751;

  NOR2_X1 U365 ( .A1(n630), .A2(n362), .ZN(n668) );
  AND2_X1 U366 ( .A1(n606), .A2(n605), .ZN(n547) );
  OR2_X1 U367 ( .A1(n602), .A2(n601), .ZN(n346) );
  OR2_X1 U368 ( .A1(n501), .A2(n500), .ZN(n531) );
  BUF_X1 U369 ( .A(n558), .Z(n637) );
  XNOR2_X1 U370 ( .A(G113), .B(KEYINPUT74), .ZN(n395) );
  NOR2_X1 U371 ( .A1(n629), .A2(n608), .ZN(n604) );
  NOR2_X1 U372 ( .A1(n524), .A2(n647), .ZN(n525) );
  INV_X1 U373 ( .A(G953), .ZN(n739) );
  NOR2_X2 U374 ( .A1(n595), .A2(n573), .ZN(n579) );
  XNOR2_X2 U375 ( .A(n572), .B(n571), .ZN(n595) );
  AND2_X2 U376 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X2 U377 ( .A(n348), .B(KEYINPUT67), .ZN(n374) );
  XNOR2_X2 U378 ( .A(n375), .B(KEYINPUT67), .ZN(n694) );
  XNOR2_X2 U379 ( .A(n737), .B(G146), .ZN(n380) );
  XNOR2_X2 U380 ( .A(n471), .B(n357), .ZN(n737) );
  NOR2_X1 U381 ( .A1(n542), .A2(n482), .ZN(n483) );
  NOR2_X2 U382 ( .A1(n531), .A2(n503), .ZN(n391) );
  NOR2_X1 U383 ( .A1(G902), .A2(n611), .ZN(n444) );
  XNOR2_X1 U384 ( .A(n442), .B(n441), .ZN(n611) );
  OR2_X1 U385 ( .A1(n689), .A2(G902), .ZN(n493) );
  XNOR2_X1 U386 ( .A(n394), .B(G131), .ZN(n429) );
  XNOR2_X1 U387 ( .A(G119), .B(G116), .ZN(n396) );
  OR2_X2 U388 ( .A1(n458), .A2(n718), .ZN(n542) );
  NAND2_X2 U389 ( .A1(n379), .A2(KEYINPUT70), .ZN(n376) );
  NAND2_X1 U390 ( .A1(n598), .A2(n347), .ZN(n345) );
  NAND2_X1 U391 ( .A1(n345), .A2(n346), .ZN(n382) );
  AND2_X1 U392 ( .A1(n599), .A2(n383), .ZN(n347) );
  NAND2_X1 U393 ( .A1(n377), .A2(n376), .ZN(n348) );
  NAND2_X1 U394 ( .A1(n377), .A2(n376), .ZN(n349) );
  NAND2_X1 U395 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X2 U396 ( .A1(n378), .A2(KEYINPUT2), .ZN(n377) );
  NOR2_X2 U397 ( .A1(n529), .A2(n528), .ZN(n648) );
  XNOR2_X2 U398 ( .A(n350), .B(n351), .ZN(n558) );
  NOR2_X1 U399 ( .A1(n673), .A2(G902), .ZN(n350) );
  XOR2_X1 U400 ( .A(G472), .B(KEYINPUT77), .Z(n351) );
  BUF_X1 U401 ( .A(n373), .Z(n352) );
  BUF_X1 U402 ( .A(n588), .Z(n353) );
  INV_X1 U403 ( .A(n597), .ZN(n354) );
  BUF_X1 U404 ( .A(n695), .Z(n355) );
  XOR2_X1 U405 ( .A(G137), .B(G140), .Z(n486) );
  XOR2_X1 U406 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n431) );
  INV_X1 U407 ( .A(KEYINPUT72), .ZN(n394) );
  XNOR2_X1 U408 ( .A(G902), .B(KEYINPUT15), .ZN(n608) );
  XNOR2_X1 U409 ( .A(G137), .B(G101), .ZN(n399) );
  XNOR2_X1 U410 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n465) );
  NOR2_X1 U411 ( .A1(n511), .A2(n635), .ZN(n426) );
  XNOR2_X1 U412 ( .A(n499), .B(n494), .ZN(n540) );
  INV_X1 U413 ( .A(KEYINPUT39), .ZN(n361) );
  INV_X1 U414 ( .A(KEYINPUT0), .ZN(n553) );
  NOR2_X1 U415 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U416 ( .A(n455), .B(n454), .ZN(n679) );
  XNOR2_X1 U417 ( .A(n380), .B(n490), .ZN(n689) );
  NAND2_X1 U418 ( .A1(n614), .A2(G953), .ZN(n699) );
  XOR2_X1 U419 ( .A(KEYINPUT65), .B(KEYINPUT4), .Z(n356) );
  XOR2_X1 U420 ( .A(n429), .B(G134), .Z(n357) );
  XOR2_X1 U421 ( .A(KEYINPUT96), .B(G110), .Z(n358) );
  AND2_X1 U422 ( .A1(n601), .A2(n602), .ZN(n359) );
  XOR2_X1 U423 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n602) );
  INV_X1 U424 ( .A(n363), .ZN(n523) );
  BUF_X1 U425 ( .A(n748), .Z(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n525), .ZN(n539) );
  NOR2_X1 U427 ( .A1(n547), .A2(KEYINPUT2), .ZN(n362) );
  NOR2_X1 U428 ( .A1(n547), .A2(KEYINPUT2), .ZN(n629) );
  NOR2_X1 U429 ( .A1(n540), .A2(n631), .ZN(n562) );
  NOR2_X2 U430 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X2 U431 ( .A(n475), .B(n364), .ZN(n363) );
  AND2_X1 U432 ( .A1(n476), .A2(G210), .ZN(n364) );
  NAND2_X1 U433 ( .A1(n435), .A2(n366), .ZN(n367) );
  NAND2_X1 U434 ( .A1(n365), .A2(n434), .ZN(n368) );
  NAND2_X1 U435 ( .A1(n367), .A2(n368), .ZN(n442) );
  INV_X1 U436 ( .A(n435), .ZN(n365) );
  INV_X1 U437 ( .A(n434), .ZN(n366) );
  INV_X1 U438 ( .A(n632), .ZN(n369) );
  BUF_X2 U439 ( .A(n540), .Z(n632) );
  OR2_X1 U440 ( .A1(n497), .A2(n558), .ZN(n498) );
  INV_X1 U441 ( .A(n523), .ZN(n370) );
  AND2_X1 U442 ( .A1(n390), .A2(n389), .ZN(n371) );
  AND2_X1 U443 ( .A1(n594), .A2(n704), .ZN(n389) );
  XNOR2_X2 U444 ( .A(n526), .B(KEYINPUT40), .ZN(n751) );
  OR2_X1 U445 ( .A1(n621), .A2(n609), .ZN(n378) );
  NAND2_X1 U446 ( .A1(n384), .A2(n381), .ZN(n372) );
  NOR2_X2 U447 ( .A1(n670), .A2(G953), .ZN(n672) );
  XNOR2_X1 U448 ( .A(n349), .B(KEYINPUT67), .ZN(n373) );
  NAND2_X1 U449 ( .A1(n604), .A2(n603), .ZN(n379) );
  NAND2_X1 U450 ( .A1(n599), .A2(n598), .ZN(n387) );
  NAND2_X1 U451 ( .A1(n595), .A2(KEYINPUT71), .ZN(n599) );
  XNOR2_X1 U452 ( .A(n380), .B(n404), .ZN(n673) );
  NAND2_X1 U453 ( .A1(n384), .A2(n381), .ZN(n607) );
  NAND2_X1 U454 ( .A1(n382), .A2(n371), .ZN(n381) );
  INV_X1 U455 ( .A(n602), .ZN(n383) );
  AND2_X2 U456 ( .A1(n385), .A2(n386), .ZN(n384) );
  NAND2_X1 U457 ( .A1(n388), .A2(n602), .ZN(n385) );
  NAND2_X1 U458 ( .A1(n387), .A2(n359), .ZN(n386) );
  NAND2_X1 U459 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U460 ( .A1(n580), .A2(KEYINPUT44), .ZN(n390) );
  NOR2_X1 U461 ( .A1(n656), .A2(n655), .ZN(n392) );
  XNOR2_X1 U462 ( .A(KEYINPUT88), .B(KEYINPUT46), .ZN(n534) );
  XOR2_X1 U463 ( .A(KEYINPUT62), .B(n673), .Z(n674) );
  INV_X1 U464 ( .A(KEYINPUT60), .ZN(n616) );
  XNOR2_X2 U465 ( .A(G143), .B(KEYINPUT66), .ZN(n393) );
  XNOR2_X2 U466 ( .A(n393), .B(G128), .ZN(n448) );
  XNOR2_X2 U467 ( .A(n448), .B(n356), .ZN(n471) );
  XNOR2_X1 U468 ( .A(n396), .B(n395), .ZN(n398) );
  XNOR2_X1 U469 ( .A(KEYINPUT75), .B(KEYINPUT3), .ZN(n397) );
  XNOR2_X1 U470 ( .A(n398), .B(n397), .ZN(n463) );
  NOR2_X1 U471 ( .A1(G953), .A2(G237), .ZN(n436) );
  NAND2_X1 U472 ( .A1(n436), .A2(G210), .ZN(n400) );
  XNOR2_X1 U473 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U474 ( .A(KEYINPUT79), .B(KEYINPUT5), .ZN(n401) );
  XNOR2_X1 U475 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n463), .B(n403), .ZN(n404) );
  XNOR2_X1 U477 ( .A(n558), .B(KEYINPUT6), .ZN(n574) );
  NAND2_X1 U478 ( .A1(G237), .A2(G234), .ZN(n405) );
  XNOR2_X1 U479 ( .A(n405), .B(KEYINPUT94), .ZN(n406) );
  XNOR2_X1 U480 ( .A(KEYINPUT14), .B(n406), .ZN(n409) );
  AND2_X1 U481 ( .A1(G953), .A2(G902), .ZN(n407) );
  NAND2_X1 U482 ( .A1(n409), .A2(n407), .ZN(n548) );
  XOR2_X1 U483 ( .A(n548), .B(KEYINPUT107), .Z(n408) );
  NOR2_X1 U484 ( .A1(G900), .A2(n408), .ZN(n410) );
  NAND2_X1 U485 ( .A1(G952), .A2(n409), .ZN(n659) );
  NOR2_X1 U486 ( .A1(n659), .A2(G953), .ZN(n550) );
  NOR2_X1 U487 ( .A1(n410), .A2(n550), .ZN(n511) );
  XNOR2_X1 U488 ( .A(G128), .B(G119), .ZN(n411) );
  XNOR2_X1 U489 ( .A(n358), .B(n411), .ZN(n413) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n412) );
  XNOR2_X1 U491 ( .A(n413), .B(n412), .ZN(n417) );
  NAND2_X1 U492 ( .A1(n739), .A2(G234), .ZN(n415) );
  XNOR2_X1 U493 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n414) );
  XNOR2_X1 U494 ( .A(n415), .B(n414), .ZN(n446) );
  NAND2_X1 U495 ( .A1(G221), .A2(n446), .ZN(n416) );
  XNOR2_X1 U496 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X2 U497 ( .A(G146), .B(G125), .ZN(n466) );
  XNOR2_X1 U498 ( .A(n466), .B(KEYINPUT10), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n486), .B(n435), .ZN(n736) );
  XNOR2_X1 U500 ( .A(n418), .B(n736), .ZN(n685) );
  INV_X1 U501 ( .A(G902), .ZN(n474) );
  NAND2_X1 U502 ( .A1(n685), .A2(n474), .ZN(n423) );
  XOR2_X1 U503 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n421) );
  NAND2_X1 U504 ( .A1(n608), .A2(G234), .ZN(n419) );
  XNOR2_X1 U505 ( .A(n419), .B(KEYINPUT20), .ZN(n424) );
  AND2_X1 U506 ( .A1(n424), .A2(G217), .ZN(n420) );
  XNOR2_X1 U507 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X2 U508 ( .A(n423), .B(n422), .ZN(n635) );
  AND2_X1 U509 ( .A1(n424), .A2(G221), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n425), .B(KEYINPUT21), .ZN(n634) );
  NAND2_X1 U511 ( .A1(n426), .A2(n634), .ZN(n497) );
  INV_X1 U512 ( .A(n497), .ZN(n427) );
  NAND2_X1 U513 ( .A1(n574), .A2(n427), .ZN(n428) );
  XNOR2_X1 U514 ( .A(n428), .B(KEYINPUT108), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n429), .B(KEYINPUT99), .ZN(n433) );
  XNOR2_X1 U516 ( .A(G140), .B(KEYINPUT11), .ZN(n430) );
  XNOR2_X1 U517 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U518 ( .A(n433), .B(n432), .ZN(n434) );
  NAND2_X1 U519 ( .A1(n436), .A2(G214), .ZN(n438) );
  XNOR2_X1 U520 ( .A(G143), .B(G122), .ZN(n437) );
  XNOR2_X1 U521 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U522 ( .A(G104), .B(G113), .Z(n439) );
  XNOR2_X1 U523 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U524 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n443) );
  XNOR2_X1 U525 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U526 ( .A(n445), .B(G475), .ZN(n527) );
  AND2_X1 U527 ( .A1(n446), .A2(G217), .ZN(n447) );
  XNOR2_X1 U528 ( .A(n448), .B(n447), .ZN(n455) );
  XOR2_X1 U529 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n450) );
  XNOR2_X1 U530 ( .A(G107), .B(G134), .ZN(n449) );
  XNOR2_X1 U531 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U532 ( .A(n451), .B(KEYINPUT7), .Z(n453) );
  XNOR2_X1 U533 ( .A(G116), .B(G122), .ZN(n452) );
  XNOR2_X1 U534 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U535 ( .A1(n679), .A2(n474), .ZN(n457) );
  XOR2_X1 U536 ( .A(G478), .B(KEYINPUT103), .Z(n456) );
  XNOR2_X1 U537 ( .A(n457), .B(n456), .ZN(n528) );
  OR2_X1 U538 ( .A1(n527), .A2(n528), .ZN(n718) );
  XNOR2_X1 U539 ( .A(G101), .B(G104), .ZN(n459) );
  INV_X1 U540 ( .A(n459), .ZN(n461) );
  XNOR2_X1 U541 ( .A(G107), .B(G110), .ZN(n460) );
  XNOR2_X1 U542 ( .A(n461), .B(n460), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT16), .B(G122), .ZN(n462) );
  XNOR2_X1 U544 ( .A(n484), .B(n462), .ZN(n464) );
  XNOR2_X1 U545 ( .A(n464), .B(n463), .ZN(n730) );
  XNOR2_X1 U546 ( .A(n466), .B(n465), .ZN(n469) );
  NAND2_X1 U547 ( .A1(n739), .A2(G224), .ZN(n467) );
  XNOR2_X1 U548 ( .A(n467), .B(KEYINPUT81), .ZN(n468) );
  XNOR2_X1 U549 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U550 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U551 ( .A(n730), .B(n472), .ZN(n695) );
  NAND2_X1 U552 ( .A1(n695), .A2(n608), .ZN(n475) );
  INV_X1 U553 ( .A(G237), .ZN(n473) );
  NAND2_X1 U554 ( .A1(n474), .A2(n473), .ZN(n476) );
  NAND2_X1 U555 ( .A1(n476), .A2(G214), .ZN(n477) );
  XNOR2_X1 U556 ( .A(n477), .B(KEYINPUT93), .ZN(n646) );
  INV_X1 U557 ( .A(n646), .ZN(n478) );
  NAND2_X1 U558 ( .A1(n363), .A2(n478), .ZN(n480) );
  INV_X1 U559 ( .A(KEYINPUT90), .ZN(n479) );
  XNOR2_X2 U560 ( .A(n480), .B(n479), .ZN(n502) );
  BUF_X1 U561 ( .A(n502), .Z(n481) );
  INV_X1 U562 ( .A(n481), .ZN(n482) );
  XNOR2_X1 U563 ( .A(n483), .B(KEYINPUT36), .ZN(n495) );
  BUF_X1 U564 ( .A(n484), .Z(n485) );
  XOR2_X1 U565 ( .A(n486), .B(KEYINPUT80), .Z(n488) );
  NAND2_X1 U566 ( .A1(G227), .A2(n739), .ZN(n487) );
  XNOR2_X1 U567 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U568 ( .A(n485), .B(n489), .ZN(n490) );
  INV_X1 U569 ( .A(KEYINPUT73), .ZN(n491) );
  XNOR2_X1 U570 ( .A(n491), .B(G469), .ZN(n492) );
  XNOR2_X2 U571 ( .A(n493), .B(n492), .ZN(n499) );
  XNOR2_X1 U572 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n494) );
  NAND2_X1 U573 ( .A1(n495), .A2(n369), .ZN(n496) );
  XNOR2_X2 U574 ( .A(n496), .B(KEYINPUT112), .ZN(n748) );
  XNOR2_X1 U575 ( .A(n498), .B(KEYINPUT28), .ZN(n501) );
  INV_X1 U576 ( .A(n499), .ZN(n500) );
  XNOR2_X2 U577 ( .A(n502), .B(KEYINPUT19), .ZN(n552) );
  BUF_X1 U578 ( .A(n552), .Z(n503) );
  NAND2_X1 U579 ( .A1(n527), .A2(n528), .ZN(n504) );
  XOR2_X1 U580 ( .A(n504), .B(KEYINPUT104), .Z(n712) );
  INV_X1 U581 ( .A(n712), .ZN(n721) );
  NAND2_X1 U582 ( .A1(n721), .A2(n718), .ZN(n650) );
  NAND2_X1 U583 ( .A1(n391), .A2(n650), .ZN(n518) );
  NAND2_X1 U584 ( .A1(n518), .A2(KEYINPUT47), .ZN(n516) );
  OR2_X2 U585 ( .A1(n558), .A2(n646), .ZN(n505) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n506) );
  NAND2_X1 U587 ( .A1(n505), .A2(n506), .ZN(n510) );
  INV_X1 U588 ( .A(n505), .ZN(n508) );
  INV_X1 U589 ( .A(n506), .ZN(n507) );
  NAND2_X1 U590 ( .A1(n508), .A2(n507), .ZN(n509) );
  NAND2_X1 U591 ( .A1(n510), .A2(n509), .ZN(n513) );
  NAND2_X1 U592 ( .A1(n635), .A2(n634), .ZN(n631) );
  INV_X1 U593 ( .A(n631), .ZN(n561) );
  NAND2_X1 U594 ( .A1(n499), .A2(n561), .ZN(n589) );
  NOR2_X1 U595 ( .A1(n589), .A2(n511), .ZN(n512) );
  NAND2_X1 U596 ( .A1(n513), .A2(n512), .ZN(n524) );
  INV_X1 U597 ( .A(n528), .ZN(n514) );
  NOR2_X1 U598 ( .A1(n527), .A2(n514), .ZN(n569) );
  NAND2_X1 U599 ( .A1(n569), .A2(n370), .ZN(n515) );
  OR2_X1 U600 ( .A1(n524), .A2(n515), .ZN(n618) );
  NAND2_X1 U601 ( .A1(n516), .A2(n618), .ZN(n517) );
  XNOR2_X1 U602 ( .A(n517), .B(KEYINPUT84), .ZN(n521) );
  NOR2_X1 U603 ( .A1(KEYINPUT47), .A2(n518), .ZN(n519) );
  XNOR2_X1 U604 ( .A(n519), .B(KEYINPUT78), .ZN(n520) );
  NOR2_X1 U605 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U606 ( .A1(n748), .A2(n522), .ZN(n537) );
  XOR2_X1 U607 ( .A(KEYINPUT38), .B(n523), .Z(n647) );
  INV_X1 U608 ( .A(n718), .ZN(n716) );
  NAND2_X1 U609 ( .A1(n539), .A2(n716), .ZN(n526) );
  NOR2_X1 U610 ( .A1(n647), .A2(n646), .ZN(n651) );
  INV_X1 U611 ( .A(n527), .ZN(n529) );
  NAND2_X1 U612 ( .A1(n651), .A2(n648), .ZN(n530) );
  XOR2_X1 U613 ( .A(KEYINPUT41), .B(n530), .Z(n662) );
  NOR2_X1 U614 ( .A1(n662), .A2(n531), .ZN(n533) );
  XNOR2_X1 U615 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n532) );
  XNOR2_X1 U616 ( .A(n533), .B(n532), .ZN(n750) );
  NAND2_X1 U617 ( .A1(n751), .A2(n750), .ZN(n535) );
  XNOR2_X1 U618 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U619 ( .A(n538), .B(KEYINPUT48), .ZN(n606) );
  NAND2_X1 U620 ( .A1(n539), .A2(n712), .ZN(n724) );
  NAND2_X1 U621 ( .A1(n632), .A2(n478), .ZN(n541) );
  OR2_X1 U622 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U623 ( .A(n543), .B(KEYINPUT43), .ZN(n544) );
  NAND2_X1 U624 ( .A1(n544), .A2(n523), .ZN(n545) );
  XNOR2_X1 U625 ( .A(n545), .B(KEYINPUT109), .ZN(n747) );
  INV_X1 U626 ( .A(n747), .ZN(n546) );
  AND2_X1 U627 ( .A1(n724), .A2(n546), .ZN(n605) );
  NOR2_X1 U628 ( .A1(n548), .A2(G898), .ZN(n549) );
  NOR2_X2 U629 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X2 U630 ( .A(n554), .B(n553), .ZN(n584) );
  NAND2_X1 U631 ( .A1(n648), .A2(n634), .ZN(n555) );
  NOR2_X1 U632 ( .A1(n584), .A2(n555), .ZN(n557) );
  XOR2_X1 U633 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n556) );
  XNOR2_X1 U634 ( .A(n557), .B(n556), .ZN(n575) );
  INV_X1 U635 ( .A(n637), .ZN(n590) );
  NOR2_X1 U636 ( .A1(n590), .A2(n635), .ZN(n559) );
  NAND2_X1 U637 ( .A1(n632), .A2(n559), .ZN(n560) );
  NOR2_X1 U638 ( .A1(n575), .A2(n560), .ZN(n620) );
  OR2_X1 U639 ( .A1(n620), .A2(KEYINPUT71), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n584), .B(KEYINPUT95), .ZN(n588) );
  NAND2_X1 U641 ( .A1(n562), .A2(n574), .ZN(n566) );
  XNOR2_X1 U642 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n564) );
  XNOR2_X1 U643 ( .A(KEYINPUT76), .B(KEYINPUT91), .ZN(n563) );
  XNOR2_X1 U644 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U645 ( .A(n566), .B(n565), .ZN(n655) );
  INV_X1 U646 ( .A(n655), .ZN(n663) );
  NAND2_X1 U647 ( .A1(n588), .A2(n663), .ZN(n568) );
  INV_X1 U648 ( .A(KEYINPUT34), .ZN(n567) );
  XNOR2_X1 U649 ( .A(n568), .B(n567), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U651 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n571) );
  NOR2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n581) );
  NOR2_X1 U653 ( .A1(n632), .A2(n635), .ZN(n576) );
  NAND2_X1 U654 ( .A1(n581), .A2(n576), .ZN(n578) );
  XOR2_X1 U655 ( .A(KEYINPUT83), .B(KEYINPUT32), .Z(n577) );
  XNOR2_X2 U656 ( .A(n578), .B(n577), .ZN(n619) );
  NAND2_X1 U657 ( .A1(n579), .A2(n619), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n581), .A2(n632), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n582), .B(KEYINPUT89), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n583), .A2(n635), .ZN(n704) );
  OR2_X1 U661 ( .A1(n637), .A2(n631), .ZN(n585) );
  OR2_X1 U662 ( .A1(n632), .A2(n585), .ZN(n642) );
  NOR2_X1 U663 ( .A1(n584), .A2(n642), .ZN(n587) );
  XNOR2_X1 U664 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n586) );
  XNOR2_X1 U665 ( .A(n587), .B(n586), .ZN(n720) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n353), .A2(n591), .ZN(n709) );
  NAND2_X1 U668 ( .A1(n720), .A2(n709), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n592), .A2(n650), .ZN(n593) );
  XOR2_X1 U670 ( .A(KEYINPUT105), .B(n593), .Z(n594) );
  INV_X1 U671 ( .A(n595), .ZN(n597) );
  NOR2_X1 U672 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U674 ( .A(n620), .ZN(n600) );
  AND2_X1 U675 ( .A1(n619), .A2(n600), .ZN(n601) );
  INV_X1 U676 ( .A(KEYINPUT2), .ZN(n622) );
  NAND2_X1 U677 ( .A1(n372), .A2(n622), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n738) );
  NOR2_X1 U679 ( .A1(n607), .A2(n738), .ZN(n621) );
  NOR2_X1 U680 ( .A1(n608), .A2(KEYINPUT70), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n694), .A2(G475), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n610) );
  XNOR2_X1 U683 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U685 ( .A(G952), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n699), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(G60) );
  XNOR2_X1 U688 ( .A(n618), .B(G143), .ZN(G45) );
  XNOR2_X1 U689 ( .A(n619), .B(G119), .ZN(G21) );
  XOR2_X1 U690 ( .A(G110), .B(n620), .Z(G12) );
  OR2_X1 U691 ( .A1(n621), .A2(n622), .ZN(n624) );
  INV_X1 U692 ( .A(n372), .ZN(n725) );
  NAND2_X1 U693 ( .A1(n725), .A2(n622), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n625), .A2(KEYINPUT86), .ZN(n628) );
  NOR2_X1 U696 ( .A1(KEYINPUT2), .A2(KEYINPUT86), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n372), .A2(n626), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U699 ( .A(KEYINPUT50), .B(n633), .Z(n640) );
  NOR2_X1 U700 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U701 ( .A(n636), .B(KEYINPUT49), .ZN(n638) );
  NAND2_X1 U702 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U703 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U704 ( .A(n641), .B(KEYINPUT117), .ZN(n643) );
  NAND2_X1 U705 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U706 ( .A(KEYINPUT51), .B(n644), .ZN(n645) );
  NOR2_X1 U707 ( .A1(n645), .A2(n662), .ZN(n657) );
  NAND2_X1 U708 ( .A1(n647), .A2(n646), .ZN(n649) );
  AND2_X1 U709 ( .A1(n649), .A2(n648), .ZN(n654) );
  NAND2_X1 U710 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U711 ( .A(KEYINPUT118), .B(n652), .Z(n653) );
  NOR2_X1 U712 ( .A1(n654), .A2(n653), .ZN(n656) );
  OR2_X1 U713 ( .A1(n657), .A2(n392), .ZN(n658) );
  XNOR2_X1 U714 ( .A(n658), .B(KEYINPUT52), .ZN(n661) );
  INV_X1 U715 ( .A(n659), .ZN(n660) );
  NAND2_X1 U716 ( .A1(n661), .A2(n660), .ZN(n666) );
  INV_X1 U717 ( .A(n662), .ZN(n664) );
  NAND2_X1 U718 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U719 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U720 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U721 ( .A(n669), .B(KEYINPUT119), .ZN(n670) );
  XNOR2_X1 U722 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n671) );
  XNOR2_X1 U723 ( .A(n672), .B(n671), .ZN(G75) );
  NAND2_X1 U724 ( .A1(n694), .A2(G472), .ZN(n675) );
  XNOR2_X1 U725 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U726 ( .A1(n676), .A2(n699), .ZN(n678) );
  XNOR2_X1 U727 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n677) );
  XNOR2_X1 U728 ( .A(n678), .B(n677), .ZN(G57) );
  INV_X1 U729 ( .A(KEYINPUT124), .ZN(n683) );
  NAND2_X1 U730 ( .A1(n373), .A2(G478), .ZN(n680) );
  XNOR2_X1 U731 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U732 ( .A1(n681), .A2(n699), .ZN(n682) );
  XNOR2_X1 U733 ( .A(n682), .B(n683), .ZN(G63) );
  XOR2_X1 U734 ( .A(n354), .B(G122), .Z(G24) );
  NAND2_X1 U735 ( .A1(n374), .A2(G217), .ZN(n684) );
  XOR2_X1 U736 ( .A(n685), .B(n684), .Z(n686) );
  INV_X1 U737 ( .A(n699), .ZN(n692) );
  NOR2_X1 U738 ( .A1(n686), .A2(n692), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n352), .A2(G469), .ZN(n691) );
  XOR2_X1 U740 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n687) );
  XNOR2_X1 U741 ( .A(n687), .B(KEYINPUT58), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U743 ( .A(n691), .B(n690), .ZN(n693) );
  NOR2_X1 U744 ( .A1(n693), .A2(n692), .ZN(G54) );
  NAND2_X1 U745 ( .A1(n374), .A2(G210), .ZN(n698) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n696) );
  XNOR2_X1 U747 ( .A(n355), .B(n696), .ZN(n697) );
  XNOR2_X1 U748 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U749 ( .A1(n700), .A2(n699), .ZN(n703) );
  XOR2_X1 U750 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n701) );
  XNOR2_X1 U751 ( .A(n701), .B(KEYINPUT87), .ZN(n702) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(G51) );
  XNOR2_X1 U753 ( .A(n704), .B(G101), .ZN(G3) );
  NOR2_X1 U754 ( .A1(n709), .A2(n718), .ZN(n706) );
  XNOR2_X1 U755 ( .A(G104), .B(KEYINPUT113), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n706), .B(n705), .ZN(G6) );
  XOR2_X1 U757 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n708) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT27), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(n711) );
  NOR2_X1 U760 ( .A1(n709), .A2(n721), .ZN(n710) );
  XOR2_X1 U761 ( .A(n711), .B(n710), .Z(G9) );
  XOR2_X1 U762 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n714) );
  NAND2_X1 U763 ( .A1(n712), .A2(n391), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U765 ( .A(G128), .B(n715), .Z(G30) );
  NAND2_X1 U766 ( .A1(n391), .A2(n716), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n717), .B(G146), .ZN(G48) );
  NOR2_X1 U768 ( .A1(n720), .A2(n718), .ZN(n719) );
  XOR2_X1 U769 ( .A(G113), .B(n719), .Z(G15) );
  NOR2_X1 U770 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U771 ( .A(KEYINPUT116), .B(n722), .Z(n723) );
  XNOR2_X1 U772 ( .A(G116), .B(n723), .ZN(G18) );
  XNOR2_X1 U773 ( .A(G134), .B(n724), .ZN(G36) );
  NAND2_X1 U774 ( .A1(n725), .A2(n739), .ZN(n729) );
  NAND2_X1 U775 ( .A1(G953), .A2(G224), .ZN(n726) );
  XNOR2_X1 U776 ( .A(KEYINPUT61), .B(n726), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G898), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n735) );
  BUF_X1 U779 ( .A(n730), .Z(n731) );
  XOR2_X1 U780 ( .A(KEYINPUT125), .B(n731), .Z(n733) );
  NOR2_X1 U781 ( .A1(G898), .A2(n739), .ZN(n732) );
  NOR2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n738), .B(n741), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n746) );
  XNOR2_X1 U787 ( .A(n741), .B(G227), .ZN(n742) );
  XNOR2_X1 U788 ( .A(n742), .B(KEYINPUT126), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(G900), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n744), .A2(G953), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n746), .A2(n745), .ZN(G72) );
  XOR2_X1 U792 ( .A(G140), .B(n747), .Z(G42) );
  XOR2_X1 U793 ( .A(G125), .B(n360), .Z(n749) );
  XNOR2_X1 U794 ( .A(KEYINPUT37), .B(n749), .ZN(G27) );
  XNOR2_X1 U795 ( .A(G137), .B(n750), .ZN(G39) );
  XNOR2_X1 U796 ( .A(G131), .B(n751), .ZN(G33) );
endmodule

