

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715;

  INV_X1 U372 ( .A(KEYINPUT3), .ZN(n390) );
  NOR2_X2 U373 ( .A1(n569), .A2(n568), .ZN(n702) );
  AND2_X2 U374 ( .A1(n714), .A2(n715), .ZN(n526) );
  NOR2_X2 U375 ( .A1(n552), .A2(n551), .ZN(n553) );
  BUF_X2 U376 ( .A(n507), .Z(n547) );
  NOR2_X1 U377 ( .A1(n627), .A2(n481), .ZN(n432) );
  INV_X1 U378 ( .A(n527), .ZN(n471) );
  INV_X1 U379 ( .A(G143), .ZN(n359) );
  XNOR2_X1 U380 ( .A(n558), .B(n557), .ZN(n569) );
  OR2_X1 U381 ( .A1(n496), .A2(KEYINPUT44), .ZN(n497) );
  XNOR2_X1 U382 ( .A(n359), .B(G128), .ZN(n413) );
  XNOR2_X1 U383 ( .A(n556), .B(KEYINPUT83), .ZN(n557) );
  XOR2_X1 U384 ( .A(G137), .B(G140), .Z(n371) );
  INV_X1 U385 ( .A(n534), .ZN(n350) );
  XNOR2_X1 U386 ( .A(n520), .B(KEYINPUT1), .ZN(n468) );
  BUF_X1 U387 ( .A(n604), .Z(n351) );
  XNOR2_X1 U388 ( .A(n360), .B(KEYINPUT4), .ZN(n361) );
  NOR2_X1 U389 ( .A1(n514), .A2(n640), .ZN(n515) );
  XNOR2_X1 U390 ( .A(n388), .B(n362), .ZN(n701) );
  XNOR2_X1 U391 ( .A(n371), .B(KEYINPUT91), .ZN(n362) );
  INV_X2 U392 ( .A(G953), .ZN(n704) );
  NOR2_X1 U393 ( .A1(n667), .A2(n666), .ZN(n671) );
  XNOR2_X1 U394 ( .A(n547), .B(KEYINPUT38), .ZN(n628) );
  XNOR2_X1 U395 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n501) );
  NOR2_X1 U396 ( .A1(n484), .A2(n462), .ZN(n632) );
  XNOR2_X1 U397 ( .A(n431), .B(KEYINPUT0), .ZN(n464) );
  INV_X1 U398 ( .A(KEYINPUT28), .ZN(n518) );
  BUF_X1 U399 ( .A(n464), .Z(n481) );
  XNOR2_X1 U400 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U401 ( .A(n701), .B(n353), .ZN(n677) );
  XNOR2_X1 U402 ( .A(n368), .B(n395), .ZN(n353) );
  XNOR2_X1 U403 ( .A(n585), .B(KEYINPUT87), .ZN(n685) );
  XNOR2_X1 U404 ( .A(n533), .B(KEYINPUT36), .ZN(n535) );
  INV_X1 U405 ( .A(KEYINPUT84), .ZN(n488) );
  NOR2_X1 U406 ( .A1(G953), .A2(n672), .ZN(n674) );
  XNOR2_X1 U407 ( .A(n413), .B(G134), .ZN(n447) );
  NOR2_X1 U408 ( .A1(n677), .A2(G902), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n679), .B(n678), .ZN(n680) );
  BUF_X1 U410 ( .A(n675), .Z(n681) );
  AND2_X2 U411 ( .A1(n580), .A2(n663), .ZN(n675) );
  NAND2_X1 U412 ( .A1(n574), .A2(n573), .ZN(n580) );
  AND2_X1 U413 ( .A1(n535), .A2(n534), .ZN(n354) );
  XOR2_X1 U414 ( .A(n370), .B(n700), .Z(n355) );
  AND2_X1 U415 ( .A1(G214), .A2(n438), .ZN(n356) );
  OR2_X1 U416 ( .A1(n619), .A2(n614), .ZN(n357) );
  XOR2_X1 U417 ( .A(n582), .B(n581), .Z(n358) );
  INV_X1 U418 ( .A(n628), .ZN(n630) );
  INV_X1 U419 ( .A(KEYINPUT67), .ZN(n540) );
  XNOR2_X1 U420 ( .A(n541), .B(KEYINPUT47), .ZN(n552) );
  INV_X1 U421 ( .A(KEYINPUT75), .ZN(n396) );
  XNOR2_X1 U422 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U423 ( .A(n700), .B(n356), .ZN(n439) );
  XNOR2_X1 U424 ( .A(n399), .B(n398), .ZN(n582) );
  NOR2_X1 U425 ( .A1(n620), .A2(n530), .ZN(n531) );
  XNOR2_X1 U426 ( .A(n502), .B(n501), .ZN(n543) );
  INV_X1 U427 ( .A(n468), .ZN(n534) );
  INV_X1 U428 ( .A(n685), .ZN(n586) );
  NAND2_X1 U429 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U430 ( .A(G131), .B(KEYINPUT68), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n447), .B(n361), .ZN(n388) );
  INV_X1 U432 ( .A(KEYINPUT65), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n363), .B(G101), .ZN(n410) );
  XOR2_X1 U434 ( .A(G146), .B(n410), .Z(n395) );
  XNOR2_X2 U435 ( .A(G110), .B(G107), .ZN(n365) );
  INV_X1 U436 ( .A(G104), .ZN(n364) );
  XNOR2_X2 U437 ( .A(n365), .B(n364), .ZN(n405) );
  NAND2_X1 U438 ( .A1(G227), .A2(n704), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n366), .B(KEYINPUT92), .ZN(n367) );
  XNOR2_X1 U440 ( .A(n405), .B(n367), .ZN(n368) );
  XNOR2_X2 U441 ( .A(n352), .B(G469), .ZN(n520) );
  NAND2_X1 U442 ( .A1(G234), .A2(n704), .ZN(n369) );
  XOR2_X1 U443 ( .A(KEYINPUT8), .B(n369), .Z(n454) );
  NAND2_X1 U444 ( .A1(G221), .A2(n454), .ZN(n370) );
  XNOR2_X2 U445 ( .A(G146), .B(G125), .ZN(n409) );
  XNOR2_X1 U446 ( .A(n409), .B(KEYINPUT10), .ZN(n700) );
  XNOR2_X1 U447 ( .A(G119), .B(G110), .ZN(n372) );
  XNOR2_X1 U448 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U449 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n374) );
  XNOR2_X1 U450 ( .A(G128), .B(KEYINPUT23), .ZN(n373) );
  XNOR2_X1 U451 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U452 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U453 ( .A(n355), .B(n377), .ZN(n592) );
  INV_X1 U454 ( .A(G902), .ZN(n420) );
  NAND2_X1 U455 ( .A1(n592), .A2(n420), .ZN(n383) );
  XOR2_X1 U456 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n381) );
  XNOR2_X1 U457 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n378) );
  XNOR2_X1 U458 ( .A(n378), .B(G902), .ZN(n418) );
  NAND2_X1 U459 ( .A1(n418), .A2(G234), .ZN(n379) );
  XNOR2_X1 U460 ( .A(n379), .B(KEYINPUT20), .ZN(n384) );
  NAND2_X1 U461 ( .A1(n384), .A2(G217), .ZN(n380) );
  XNOR2_X1 U462 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X2 U463 ( .A(n383), .B(n382), .ZN(n514) );
  XOR2_X1 U464 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n386) );
  NAND2_X1 U465 ( .A1(n384), .A2(G221), .ZN(n385) );
  XNOR2_X1 U466 ( .A(n386), .B(n385), .ZN(n640) );
  XOR2_X1 U467 ( .A(KEYINPUT96), .B(n640), .Z(n463) );
  NAND2_X1 U468 ( .A1(n514), .A2(n463), .ZN(n387) );
  XNOR2_X1 U469 ( .A(n387), .B(KEYINPUT66), .ZN(n647) );
  NOR2_X2 U470 ( .A1(n468), .A2(n647), .ZN(n478) );
  XOR2_X1 U471 ( .A(G137), .B(KEYINPUT5), .Z(n389) );
  XNOR2_X1 U472 ( .A(n388), .B(n389), .ZN(n399) );
  XNOR2_X1 U473 ( .A(n390), .B(G119), .ZN(n392) );
  XNOR2_X1 U474 ( .A(G116), .B(G113), .ZN(n391) );
  XNOR2_X1 U475 ( .A(n392), .B(n391), .ZN(n407) );
  NOR2_X1 U476 ( .A1(G953), .A2(G237), .ZN(n438) );
  AND2_X1 U477 ( .A1(n438), .A2(G210), .ZN(n393) );
  XNOR2_X1 U478 ( .A(n407), .B(n393), .ZN(n394) );
  XNOR2_X1 U479 ( .A(n395), .B(n394), .ZN(n397) );
  NAND2_X1 U480 ( .A1(n582), .A2(n420), .ZN(n400) );
  XNOR2_X2 U481 ( .A(n400), .B(G472), .ZN(n480) );
  XNOR2_X1 U482 ( .A(n480), .B(KEYINPUT6), .ZN(n527) );
  NAND2_X1 U483 ( .A1(n478), .A2(n471), .ZN(n402) );
  INV_X1 U484 ( .A(KEYINPUT33), .ZN(n401) );
  XNOR2_X1 U485 ( .A(n402), .B(n401), .ZN(n627) );
  XNOR2_X1 U486 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n403) );
  XNOR2_X1 U487 ( .A(n403), .B(G122), .ZN(n404) );
  XNOR2_X1 U488 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U489 ( .A(n407), .B(n406), .ZN(n686) );
  XNOR2_X1 U490 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n408) );
  XNOR2_X1 U491 ( .A(n409), .B(n408), .ZN(n411) );
  XNOR2_X1 U492 ( .A(n411), .B(n410), .ZN(n416) );
  NAND2_X1 U493 ( .A1(n704), .A2(G224), .ZN(n412) );
  XNOR2_X1 U494 ( .A(n412), .B(KEYINPUT4), .ZN(n414) );
  XNOR2_X1 U495 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U496 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U497 ( .A(n686), .B(n417), .ZN(n604) );
  INV_X1 U498 ( .A(n418), .ZN(n572) );
  OR2_X2 U499 ( .A1(n604), .A2(n572), .ZN(n423) );
  INV_X1 U500 ( .A(G237), .ZN(n419) );
  NAND2_X1 U501 ( .A1(n420), .A2(n419), .ZN(n424) );
  NAND2_X1 U502 ( .A1(n424), .A2(G210), .ZN(n421) );
  XNOR2_X1 U503 ( .A(n421), .B(KEYINPUT78), .ZN(n422) );
  XNOR2_X1 U504 ( .A(n423), .B(n422), .ZN(n507) );
  NAND2_X1 U505 ( .A1(n424), .A2(G214), .ZN(n561) );
  INV_X1 U506 ( .A(n561), .ZN(n629) );
  OR2_X2 U507 ( .A1(n507), .A2(n629), .ZN(n532) );
  XNOR2_X2 U508 ( .A(n532), .B(KEYINPUT19), .ZN(n537) );
  NAND2_X1 U509 ( .A1(G234), .A2(G237), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n425), .B(KEYINPUT14), .ZN(n428) );
  NAND2_X1 U511 ( .A1(n428), .A2(G952), .ZN(n426) );
  XOR2_X1 U512 ( .A(KEYINPUT89), .B(n426), .Z(n660) );
  INV_X1 U513 ( .A(n660), .ZN(n427) );
  NAND2_X1 U514 ( .A1(n427), .A2(n704), .ZN(n506) );
  NAND2_X1 U515 ( .A1(G902), .A2(n428), .ZN(n503) );
  XOR2_X1 U516 ( .A(G898), .B(KEYINPUT90), .Z(n694) );
  NAND2_X1 U517 ( .A1(G953), .A2(n694), .ZN(n689) );
  OR2_X1 U518 ( .A1(n503), .A2(n689), .ZN(n429) );
  NAND2_X1 U519 ( .A1(n506), .A2(n429), .ZN(n430) );
  NAND2_X1 U520 ( .A1(n537), .A2(n430), .ZN(n431) );
  XNOR2_X1 U521 ( .A(n432), .B(KEYINPUT34), .ZN(n460) );
  XOR2_X1 U522 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n434) );
  XNOR2_X1 U523 ( .A(G131), .B(KEYINPUT99), .ZN(n433) );
  XNOR2_X1 U524 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U525 ( .A(n435), .B(G140), .Z(n437) );
  XNOR2_X1 U526 ( .A(G122), .B(G104), .ZN(n436) );
  XNOR2_X1 U527 ( .A(n437), .B(n436), .ZN(n440) );
  XOR2_X1 U528 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n442) );
  XNOR2_X1 U529 ( .A(G143), .B(G113), .ZN(n441) );
  XNOR2_X1 U530 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U531 ( .A(n444), .B(n443), .ZN(n597) );
  NOR2_X1 U532 ( .A1(G902), .A2(n597), .ZN(n446) );
  XNOR2_X1 U533 ( .A(KEYINPUT13), .B(G475), .ZN(n445) );
  XNOR2_X1 U534 ( .A(n446), .B(n445), .ZN(n484) );
  INV_X1 U535 ( .A(n484), .ZN(n459) );
  XOR2_X1 U536 ( .A(KEYINPUT7), .B(G107), .Z(n449) );
  XNOR2_X1 U537 ( .A(G116), .B(G122), .ZN(n448) );
  XNOR2_X1 U538 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U539 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n451) );
  XNOR2_X1 U540 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n450) );
  XNOR2_X1 U541 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U542 ( .A(n453), .B(n452), .Z(n456) );
  NAND2_X1 U543 ( .A1(G217), .A2(n454), .ZN(n455) );
  XNOR2_X1 U544 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n447), .B(n457), .ZN(n682) );
  NOR2_X1 U546 ( .A1(n682), .A2(G902), .ZN(n458) );
  XNOR2_X1 U547 ( .A(n458), .B(G478), .ZN(n485) );
  NOR2_X1 U548 ( .A1(n459), .A2(n485), .ZN(n548) );
  NAND2_X1 U549 ( .A1(n460), .A2(n548), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n461), .B(KEYINPUT35), .ZN(n712) );
  INV_X1 U551 ( .A(n485), .ZN(n462) );
  NAND2_X1 U552 ( .A1(n632), .A2(n463), .ZN(n465) );
  NOR2_X1 U553 ( .A1(n465), .A2(n464), .ZN(n467) );
  XOR2_X1 U554 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n466) );
  XNOR2_X1 U555 ( .A(n467), .B(n466), .ZN(n472) );
  BUF_X2 U556 ( .A(n480), .Z(n645) );
  NOR2_X1 U557 ( .A1(n645), .A2(n514), .ZN(n469) );
  NAND2_X1 U558 ( .A1(n350), .A2(n469), .ZN(n470) );
  NOR2_X1 U559 ( .A1(n472), .A2(n470), .ZN(n589) );
  NOR2_X1 U560 ( .A1(n712), .A2(n589), .ZN(n477) );
  XNOR2_X1 U561 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n476) );
  NOR2_X1 U562 ( .A1(n472), .A2(n471), .ZN(n487) );
  XNOR2_X1 U563 ( .A(n514), .B(KEYINPUT104), .ZN(n641) );
  NOR2_X1 U564 ( .A1(n468), .A2(n641), .ZN(n473) );
  XNOR2_X1 U565 ( .A(n473), .B(KEYINPUT106), .ZN(n474) );
  NAND2_X1 U566 ( .A1(n487), .A2(n474), .ZN(n475) );
  XOR2_X1 U567 ( .A(n476), .B(n475), .Z(n713) );
  NAND2_X1 U568 ( .A1(n477), .A2(n713), .ZN(n496) );
  NAND2_X1 U569 ( .A1(n496), .A2(KEYINPUT44), .ZN(n494) );
  NAND2_X1 U570 ( .A1(n478), .A2(n645), .ZN(n652) );
  NOR2_X1 U571 ( .A1(n652), .A2(n481), .ZN(n479) );
  XNOR2_X1 U572 ( .A(n479), .B(KEYINPUT31), .ZN(n623) );
  NOR2_X2 U573 ( .A1(n647), .A2(n520), .ZN(n542) );
  INV_X1 U574 ( .A(n480), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n542), .A2(n517), .ZN(n482) );
  NOR2_X1 U576 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U577 ( .A(n483), .B(KEYINPUT97), .ZN(n610) );
  NAND2_X1 U578 ( .A1(n623), .A2(n610), .ZN(n486) );
  NAND2_X1 U579 ( .A1(n484), .A2(n485), .ZN(n620) );
  OR2_X1 U580 ( .A1(n485), .A2(n484), .ZN(n622) );
  NAND2_X1 U581 ( .A1(n620), .A2(n622), .ZN(n635) );
  NAND2_X1 U582 ( .A1(n486), .A2(n635), .ZN(n491) );
  NAND2_X1 U583 ( .A1(n487), .A2(n350), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U585 ( .A1(n490), .A2(n641), .ZN(n591) );
  NAND2_X1 U586 ( .A1(n491), .A2(n591), .ZN(n492) );
  XNOR2_X1 U587 ( .A(n492), .B(KEYINPUT105), .ZN(n493) );
  NAND2_X1 U588 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U589 ( .A(n495), .B(KEYINPUT85), .ZN(n498) );
  NAND2_X1 U590 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U591 ( .A(n499), .B(KEYINPUT45), .ZN(n577) );
  NAND2_X1 U592 ( .A1(n577), .A2(n572), .ZN(n500) );
  XNOR2_X1 U593 ( .A(n500), .B(KEYINPUT81), .ZN(n571) );
  NAND2_X1 U594 ( .A1(n561), .A2(n645), .ZN(n502) );
  NOR2_X1 U595 ( .A1(G900), .A2(n503), .ZN(n504) );
  NAND2_X1 U596 ( .A1(G953), .A2(n504), .ZN(n505) );
  NAND2_X1 U597 ( .A1(n506), .A2(n505), .ZN(n545) );
  AND2_X1 U598 ( .A1(n545), .A2(n628), .ZN(n508) );
  NAND2_X1 U599 ( .A1(n542), .A2(n508), .ZN(n509) );
  NOR2_X1 U600 ( .A1(n543), .A2(n509), .ZN(n511) );
  XNOR2_X1 U601 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n510) );
  XOR2_X1 U602 ( .A(n511), .B(n510), .Z(n559) );
  NOR2_X1 U603 ( .A1(n620), .A2(n559), .ZN(n513) );
  XNOR2_X1 U604 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n714) );
  NAND2_X1 U606 ( .A1(n545), .A2(n515), .ZN(n516) );
  XNOR2_X1 U607 ( .A(KEYINPUT70), .B(n516), .ZN(n528) );
  NOR2_X1 U608 ( .A1(n528), .A2(n517), .ZN(n519) );
  XNOR2_X1 U609 ( .A(n519), .B(n518), .ZN(n521) );
  NOR2_X2 U610 ( .A1(n521), .A2(n520), .ZN(n538) );
  NAND2_X1 U611 ( .A1(n628), .A2(n561), .ZN(n522) );
  XOR2_X1 U612 ( .A(KEYINPUT112), .B(n522), .Z(n634) );
  NAND2_X1 U613 ( .A1(n632), .A2(n634), .ZN(n523) );
  XNOR2_X1 U614 ( .A(KEYINPUT41), .B(n523), .ZN(n654) );
  NAND2_X1 U615 ( .A1(n538), .A2(n654), .ZN(n524) );
  XNOR2_X1 U616 ( .A(n524), .B(KEYINPUT42), .ZN(n715) );
  INV_X1 U617 ( .A(KEYINPUT46), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n526), .B(n525), .ZN(n536) );
  NOR2_X1 U619 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U620 ( .A(n529), .B(KEYINPUT107), .ZN(n530) );
  XOR2_X1 U621 ( .A(KEYINPUT108), .B(n531), .Z(n563) );
  NOR2_X1 U622 ( .A1(n563), .A2(n532), .ZN(n533) );
  NOR2_X1 U623 ( .A1(n536), .A2(n354), .ZN(n555) );
  NOR2_X1 U624 ( .A1(n539), .A2(n620), .ZN(n619) );
  NOR2_X1 U625 ( .A1(n539), .A2(n622), .ZN(n614) );
  NAND2_X1 U626 ( .A1(n357), .A2(n540), .ZN(n541) );
  INV_X1 U627 ( .A(n542), .ZN(n544) );
  NOR2_X1 U628 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U629 ( .A1(n546), .A2(n545), .ZN(n550) );
  INV_X1 U630 ( .A(n547), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n566), .A2(n548), .ZN(n549) );
  NOR2_X1 U632 ( .A1(n550), .A2(n549), .ZN(n617) );
  XNOR2_X1 U633 ( .A(KEYINPUT80), .B(n617), .ZN(n551) );
  XNOR2_X1 U634 ( .A(n553), .B(KEYINPUT74), .ZN(n554) );
  NAND2_X1 U635 ( .A1(n555), .A2(n554), .ZN(n558) );
  XNOR2_X1 U636 ( .A(KEYINPUT48), .B(KEYINPUT69), .ZN(n556) );
  OR2_X1 U637 ( .A1(n559), .A2(n622), .ZN(n560) );
  XOR2_X1 U638 ( .A(KEYINPUT113), .B(n560), .Z(n711) );
  XNOR2_X1 U639 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n350), .A2(n561), .ZN(n562) );
  NOR2_X1 U641 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U642 ( .A(n565), .B(n564), .ZN(n567) );
  NAND2_X1 U643 ( .A1(n567), .A2(n547), .ZN(n590) );
  NAND2_X1 U644 ( .A1(n711), .A2(n590), .ZN(n568) );
  XNOR2_X1 U645 ( .A(n702), .B(KEYINPUT76), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n572), .A2(KEYINPUT2), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n702), .A2(KEYINPUT2), .ZN(n576) );
  INV_X1 U649 ( .A(KEYINPUT82), .ZN(n575) );
  XNOR2_X1 U650 ( .A(n576), .B(n575), .ZN(n579) );
  BUF_X1 U651 ( .A(n577), .Z(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n663) );
  NAND2_X1 U653 ( .A1(n675), .A2(G472), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n581) );
  XNOR2_X1 U655 ( .A(n583), .B(n358), .ZN(n587) );
  INV_X1 U656 ( .A(G952), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n584), .A2(G953), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n588), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U660 ( .A(G110), .B(n589), .Z(G12) );
  XNOR2_X1 U661 ( .A(n590), .B(G140), .ZN(G42) );
  XNOR2_X1 U662 ( .A(n591), .B(G101), .ZN(G3) );
  NAND2_X1 U663 ( .A1(n681), .A2(G217), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT123), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X1 U666 ( .A1(n595), .A2(n685), .ZN(G66) );
  NAND2_X1 U667 ( .A1(n675), .A2(G475), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT64), .B(KEYINPUT59), .Z(n596) );
  XNOR2_X1 U669 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n599), .B(n598), .ZN(n600) );
  NOR2_X2 U671 ( .A1(n600), .A2(n685), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U673 ( .A1(n675), .A2(G210), .ZN(n606) );
  XOR2_X1 U674 ( .A(KEYINPUT86), .B(KEYINPUT54), .Z(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT55), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n351), .B(n603), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X2 U678 ( .A1(n607), .A2(n685), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U680 ( .A1(n610), .A2(n620), .ZN(n609) );
  XOR2_X1 U681 ( .A(G104), .B(n609), .Z(G6) );
  NOR2_X1 U682 ( .A1(n610), .A2(n622), .ZN(n612) );
  XNOR2_X1 U683 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U685 ( .A(G107), .B(n613), .ZN(G9) );
  XOR2_X1 U686 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n616) );
  XNOR2_X1 U687 ( .A(n614), .B(G128), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(G30) );
  XOR2_X1 U689 ( .A(G143), .B(n617), .Z(n618) );
  XNOR2_X1 U690 ( .A(KEYINPUT116), .B(n618), .ZN(G45) );
  XOR2_X1 U691 ( .A(G146), .B(n619), .Z(G48) );
  NOR2_X1 U692 ( .A1(n623), .A2(n620), .ZN(n621) );
  XOR2_X1 U693 ( .A(G113), .B(n621), .Z(G15) );
  NOR2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n625) );
  XNOR2_X1 U695 ( .A(G116), .B(KEYINPUT117), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(G18) );
  XNOR2_X1 U697 ( .A(G125), .B(n354), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U701 ( .A(KEYINPUT119), .B(n633), .Z(n637) );
  NAND2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U703 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U704 ( .A(KEYINPUT120), .B(n638), .Z(n639) );
  NOR2_X1 U705 ( .A1(n627), .A2(n639), .ZN(n657) );
  INV_X1 U706 ( .A(n640), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U708 ( .A(KEYINPUT49), .B(n643), .Z(n644) );
  NOR2_X1 U709 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U710 ( .A(KEYINPUT118), .B(n646), .ZN(n650) );
  NAND2_X1 U711 ( .A1(n350), .A2(n647), .ZN(n648) );
  XNOR2_X1 U712 ( .A(KEYINPUT50), .B(n648), .ZN(n649) );
  NAND2_X1 U713 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U714 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U715 ( .A(KEYINPUT51), .B(n653), .ZN(n655) );
  INV_X1 U716 ( .A(n654), .ZN(n668) );
  NOR2_X1 U717 ( .A1(n655), .A2(n668), .ZN(n656) );
  NOR2_X1 U718 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U719 ( .A(n658), .B(KEYINPUT52), .ZN(n659) );
  NOR2_X1 U720 ( .A1(n660), .A2(n659), .ZN(n667) );
  AND2_X1 U721 ( .A1(n702), .A2(n578), .ZN(n662) );
  XOR2_X1 U722 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n661) );
  NOR2_X1 U723 ( .A1(n662), .A2(n661), .ZN(n665) );
  INV_X1 U724 ( .A(n663), .ZN(n664) );
  NOR2_X1 U725 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U726 ( .A1(n668), .A2(n627), .ZN(n669) );
  XNOR2_X1 U727 ( .A(n669), .B(KEYINPUT121), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U729 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n673) );
  XNOR2_X1 U730 ( .A(n674), .B(n673), .ZN(G75) );
  NAND2_X1 U731 ( .A1(n681), .A2(G469), .ZN(n679) );
  XOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n676) );
  XNOR2_X1 U733 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U734 ( .A1(n685), .A2(n680), .ZN(G54) );
  NAND2_X1 U735 ( .A1(n681), .A2(G478), .ZN(n683) );
  XNOR2_X1 U736 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U737 ( .A1(n685), .A2(n684), .ZN(G63) );
  XOR2_X1 U738 ( .A(G101), .B(KEYINPUT125), .Z(n687) );
  XNOR2_X1 U739 ( .A(n686), .B(n687), .ZN(n688) );
  NAND2_X1 U740 ( .A1(n689), .A2(n688), .ZN(n698) );
  INV_X1 U741 ( .A(n578), .ZN(n690) );
  NOR2_X1 U742 ( .A1(n690), .A2(G953), .ZN(n696) );
  XOR2_X1 U743 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n692) );
  NAND2_X1 U744 ( .A1(G224), .A2(G953), .ZN(n691) );
  XNOR2_X1 U745 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U748 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U749 ( .A(KEYINPUT126), .B(n699), .ZN(G69) );
  XNOR2_X1 U750 ( .A(n701), .B(n700), .ZN(n706) );
  INV_X1 U751 ( .A(n706), .ZN(n703) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U753 ( .A1(n705), .A2(n704), .ZN(n710) );
  XNOR2_X1 U754 ( .A(G227), .B(n706), .ZN(n707) );
  NAND2_X1 U755 ( .A1(n707), .A2(G900), .ZN(n708) );
  NAND2_X1 U756 ( .A1(n708), .A2(G953), .ZN(n709) );
  NAND2_X1 U757 ( .A1(n710), .A2(n709), .ZN(G72) );
  XNOR2_X1 U758 ( .A(G134), .B(n711), .ZN(G36) );
  XOR2_X1 U759 ( .A(G122), .B(n712), .Z(G24) );
  XNOR2_X1 U760 ( .A(G119), .B(n713), .ZN(G21) );
  XNOR2_X1 U761 ( .A(n714), .B(G131), .ZN(G33) );
  XNOR2_X1 U762 ( .A(G137), .B(n715), .ZN(G39) );
endmodule

