//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT0), .A3(G128), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT0), .B(G128), .Z(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(new_n207), .A3(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n197), .A2(G143), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n201), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT84), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n216), .A3(G125), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G224), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n206), .A2(new_n215), .A3(new_n220), .A4(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(KEYINPUT5), .A3(G119), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G116), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(KEYINPUT66), .A3(G119), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n229), .A2(new_n230), .B1(G116), .B2(new_n228), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n231), .B2(KEYINPUT5), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT2), .B(G113), .Z(new_n233));
  AOI22_X1  g047(.A1(new_n232), .A2(G113), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n235));
  INV_X1    g049(.A(G107), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n238));
  INV_X1    g052(.A(G101), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G107), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n235), .A2(new_n242), .A3(new_n236), .A4(G104), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n239), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n236), .A2(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(KEYINPUT78), .A3(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n247), .A2(KEYINPUT78), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n234), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n255), .A3(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n231), .B(new_n233), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(G110), .B(G122), .Z(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT82), .ZN(new_n265));
  INV_X1    g079(.A(new_n260), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n251), .A2(new_n258), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n251), .B2(new_n258), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n269), .B2(KEYINPUT6), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n251), .A2(new_n258), .A3(new_n266), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n261), .A2(new_n265), .A3(KEYINPUT6), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n224), .B(new_n264), .C1(new_n270), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT85), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n271), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT82), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n263), .B1(new_n277), .B2(new_n272), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n224), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n218), .B1(new_n283), .B2(new_n221), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n218), .B(KEYINPUT86), .C1(new_n283), .C2(new_n221), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n234), .B(new_n250), .Z(new_n289));
  XNOR2_X1  g103(.A(new_n260), .B(KEYINPUT8), .ZN(new_n290));
  OAI221_X1 g104(.A(new_n271), .B1(new_n223), .B2(new_n283), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n282), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n188), .B1(new_n281), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n188), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n295), .B(new_n292), .C1(new_n275), .C2(new_n280), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT87), .ZN(new_n298));
  INV_X1    g112(.A(G221), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT9), .B(G234), .Z(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n282), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n219), .A2(G227), .ZN(new_n302));
  INV_X1    g116(.A(G140), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(G110), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n250), .A2(KEYINPUT10), .A3(new_n214), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n248), .B2(new_n249), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT79), .A3(new_n214), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n254), .A2(new_n256), .ZN(new_n315));
  INV_X1    g129(.A(new_n204), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT64), .B(G143), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n207), .B1(new_n317), .B2(new_n197), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n197), .B1(new_n191), .B2(new_n193), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n318), .A2(new_n209), .B1(new_n190), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n208), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n250), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n315), .A2(new_n316), .B1(new_n322), .B2(new_n311), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT11), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G137), .ZN(new_n326));
  INV_X1    g140(.A(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT11), .A3(G134), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n327), .B2(G134), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(KEYINPUT65), .A3(G137), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n330), .B1(new_n329), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n314), .A2(new_n323), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n337), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n250), .A2(new_n214), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n248), .A2(new_n249), .B1(new_n320), .B2(new_n208), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n322), .B1(new_n250), .B2(new_n214), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n348), .A2(new_n343), .A3(new_n344), .A4(new_n339), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n307), .B1(new_n338), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n312), .A2(KEYINPUT79), .A3(new_n214), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT79), .B1(new_n312), .B2(new_n214), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n316), .A2(new_n256), .A3(new_n254), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(KEYINPUT10), .B2(new_n341), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n339), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n314), .A2(new_n323), .A3(new_n337), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n306), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(KEYINPUT81), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT81), .B1(new_n351), .B2(new_n359), .ZN(new_n362));
  OAI21_X1  g176(.A(G469), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G469), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n282), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n337), .B1(new_n314), .B2(new_n323), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n307), .B1(new_n338), .B2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n358), .A2(new_n349), .A3(new_n347), .A4(new_n306), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n365), .B1(new_n369), .B2(new_n364), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n301), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n298), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(KEYINPUT26), .B(G101), .Z(new_n373));
  INV_X1    g187(.A(G237), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n219), .A3(G210), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT28), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n196), .B(new_n203), .C1(new_n335), .C2(new_n336), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n325), .A2(G137), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n327), .A2(G134), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR4_X1   g198(.A1(new_n319), .A2(KEYINPUT1), .A3(new_n209), .A4(new_n190), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n211), .B1(new_n198), .B2(new_n200), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n381), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT69), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n380), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n257), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n380), .B2(new_n387), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n379), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n380), .A2(new_n387), .A3(new_n390), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n390), .B1(new_n380), .B2(new_n387), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT28), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n378), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n394), .A2(KEYINPUT68), .A3(new_n378), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT68), .B1(new_n394), .B2(new_n378), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n380), .A2(new_n387), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n380), .A2(new_n387), .A3(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n257), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT31), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n394), .A2(new_n378), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT68), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n394), .A2(KEYINPUT68), .A3(new_n378), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n407), .A3(KEYINPUT31), .A4(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n399), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G472), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n282), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n407), .A2(new_n394), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(new_n378), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n393), .A2(new_n397), .A3(new_n378), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n282), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT71), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n396), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT70), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n394), .B(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n379), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n393), .ZN(new_n430));
  INV_X1    g244(.A(new_n378), .ZN(new_n431));
  NOR4_X1   g245(.A1(new_n429), .A2(new_n420), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G472), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n411), .A2(new_n407), .A3(new_n412), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n413), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n437), .B2(new_n399), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT32), .A3(new_n416), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n419), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G125), .B(G140), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT16), .ZN(new_n442));
  INV_X1    g256(.A(G125), .ZN(new_n443));
  OR3_X1    g257(.A1(new_n443), .A2(KEYINPUT16), .A3(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(G146), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n228), .A2(G128), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n209), .A2(G119), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n450), .B2(new_n447), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT24), .B(G110), .Z(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(KEYINPUT23), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT73), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n449), .C1(KEYINPUT23), .C2(new_n447), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G110), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n457), .A2(G110), .B1(new_n452), .B2(new_n453), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n442), .A2(G146), .A3(new_n444), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT74), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n441), .A2(new_n197), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G137), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n467), .B(new_n468), .Z(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n459), .A2(new_n465), .A3(new_n469), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G217), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(G234), .B2(new_n282), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(G902), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT75), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n282), .A3(new_n472), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT25), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n471), .A2(new_n481), .A3(new_n282), .A4(new_n472), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n484), .A3(new_n476), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n440), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n374), .A2(new_n219), .A3(G143), .A4(G214), .ZN(new_n489));
  INV_X1    g303(.A(G214), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n490), .A2(G237), .A3(G953), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n317), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT17), .A3(G131), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(G131), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n330), .B(new_n489), .C1(new_n317), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n446), .B(new_n493), .C1(KEYINPUT17), .C2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n441), .B(new_n197), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n489), .C1(new_n317), .C2(new_n491), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n495), .A2(new_n500), .A3(KEYINPUT88), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT88), .B1(new_n495), .B2(new_n500), .ZN(new_n502));
  OAI221_X1 g316(.A(new_n498), .B1(new_n499), .B2(new_n494), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(G104), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n505), .B(KEYINPUT90), .Z(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n441), .B(KEYINPUT19), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n197), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n463), .A2(new_n496), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n503), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n505), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n510), .B2(new_n503), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n282), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n517), .A2(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(KEYINPUT20), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n507), .ZN(new_n521));
  INV_X1    g335(.A(new_n505), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n497), .B2(new_n503), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n282), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G475), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n317), .A2(new_n209), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n189), .A2(G128), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n527), .A2(G134), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n194), .A2(G128), .ZN(new_n530));
  INV_X1    g344(.A(new_n528), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n325), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT91), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G134), .B1(new_n527), .B2(new_n528), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(new_n325), .A3(new_n531), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(G116), .B(G122), .Z(new_n538));
  OR2_X1    g352(.A1(new_n538), .A2(G107), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n225), .A2(KEYINPUT14), .A3(G122), .ZN(new_n540));
  OAI211_X1 g354(.A(G107), .B(new_n540), .C1(new_n538), .C2(KEYINPUT14), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n533), .A2(new_n537), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n530), .A2(KEYINPUT13), .A3(new_n531), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(G134), .C1(KEYINPUT13), .C2(new_n530), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n538), .B(G107), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n536), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n300), .A2(G217), .A3(new_n219), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n542), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n542), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G902), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G478), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n553), .B(G478), .C1(new_n551), .C2(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT92), .B1(new_n555), .B2(new_n556), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G952), .ZN(new_n562));
  AOI211_X1 g376(.A(G953), .B(new_n562), .C1(G234), .C2(G237), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n282), .B(new_n219), .C1(G234), .C2(G237), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT21), .B(G898), .Z(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n526), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n372), .A2(new_n488), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  OAI211_X1 g386(.A(new_n187), .B(new_n568), .C1(new_n294), .C2(new_n296), .ZN(new_n573));
  INV_X1    g387(.A(new_n550), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n542), .A2(new_n546), .A3(new_n548), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT33), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n549), .B2(new_n550), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n578), .A3(G478), .A4(new_n282), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT93), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n552), .A2(G478), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n526), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n573), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n301), .ZN(new_n585));
  INV_X1    g399(.A(new_n370), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n351), .A2(new_n359), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n364), .B1(new_n589), .B2(new_n360), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n585), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n415), .A2(new_n282), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n417), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n591), .A2(new_n594), .A3(new_n486), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n584), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT94), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT34), .B(G104), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  AOI22_X1  g413(.A1(new_n518), .A2(new_n519), .B1(G475), .B2(new_n524), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n561), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT95), .B1(new_n573), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n187), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n274), .A2(KEYINPUT85), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n279), .B1(new_n278), .B2(new_n224), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n293), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n295), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n281), .A2(new_n188), .A3(new_n293), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  INV_X1    g424(.A(new_n601), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n568), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n595), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT35), .B(G107), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  INV_X1    g432(.A(new_n594), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n559), .A2(new_n560), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n470), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n466), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n476), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n483), .A2(new_n623), .ZN(new_n624));
  AND4_X1   g438(.A1(new_n620), .A2(new_n600), .A3(new_n568), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n372), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT37), .B(G110), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G12));
  AND2_X1   g443(.A1(new_n371), .A2(new_n440), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT99), .B(G900), .Z(new_n631));
  OR3_X1    g445(.A1(new_n566), .A2(KEYINPUT100), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n566), .B2(new_n631), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n564), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT101), .Z(new_n635));
  NOR2_X1   g449(.A1(new_n601), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n630), .A2(new_n636), .A3(new_n609), .A4(new_n624), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  NAND2_X1  g452(.A1(new_n607), .A2(new_n608), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT38), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n635), .B(KEYINPUT39), .Z(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT40), .B1(new_n591), .B2(new_n642), .ZN(new_n643));
  OR3_X1    g457(.A1(new_n591), .A2(KEYINPUT40), .A3(new_n642), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n620), .A2(new_n600), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n378), .B1(new_n426), .B2(new_n428), .ZN(new_n647));
  INV_X1    g461(.A(new_n434), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n282), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(G472), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n419), .A2(new_n439), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n624), .A2(new_n603), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n645), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n194), .ZN(G45));
  INV_X1    g470(.A(new_n635), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n526), .A2(new_n582), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n630), .A2(new_n659), .A3(new_n609), .A4(new_n624), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  NAND2_X1  g475(.A1(new_n440), .A2(new_n487), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n358), .A2(new_n349), .A3(new_n347), .A4(new_n306), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n306), .B1(new_n357), .B2(new_n358), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n364), .B(new_n282), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT102), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n369), .A2(new_n364), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n369), .A2(KEYINPUT102), .A3(new_n364), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n585), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n584), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  OR2_X1    g488(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  INV_X1    g489(.A(new_n669), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n301), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n488), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n602), .B2(new_n612), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT103), .B(G116), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G18));
  NAND4_X1  g495(.A1(new_n625), .A2(new_n609), .A3(new_n677), .A4(new_n440), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  OAI21_X1  g497(.A(new_n431), .B1(new_n429), .B2(new_n430), .ZN(new_n684));
  AOI211_X1 g498(.A(G472), .B(G902), .C1(new_n684), .C2(new_n437), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT104), .B1(new_n438), .B2(new_n416), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n398), .B1(new_n436), .B2(new_n413), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n687), .B(G472), .C1(new_n688), .C2(G902), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n685), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n487), .A3(new_n568), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n297), .A2(new_n670), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n646), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n692), .A2(new_n693), .A3(new_n696), .A4(new_n646), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  NOR3_X1   g513(.A1(new_n297), .A2(new_n670), .A3(new_n658), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n684), .A2(new_n437), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n416), .A3(new_n282), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n687), .B1(new_n592), .B2(G472), .ZN(new_n703));
  INV_X1    g517(.A(new_n689), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n624), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n690), .A2(new_n707), .A3(new_n624), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NOR3_X1   g525(.A1(new_n294), .A2(new_n296), .A3(new_n603), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n365), .B(KEYINPUT107), .Z(new_n713));
  NAND3_X1  g527(.A1(new_n351), .A2(G469), .A3(new_n359), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n665), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n585), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n488), .A2(new_n712), .A3(new_n659), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n439), .A2(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n417), .A2(KEYINPUT109), .A3(new_n418), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT109), .B1(new_n417), .B2(new_n418), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n419), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n439), .A4(new_n722), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n728), .A3(new_n433), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n607), .A2(new_n187), .A3(new_n608), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n658), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n716), .A2(new_n719), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n487), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n720), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  NAND4_X1  g549(.A1(new_n488), .A2(new_n712), .A3(new_n636), .A4(new_n717), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT110), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n662), .A2(new_n730), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n636), .A4(new_n717), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  NAND3_X1  g556(.A1(new_n351), .A2(KEYINPUT45), .A3(new_n359), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n589), .A2(new_n360), .ZN(new_n744));
  OAI211_X1 g558(.A(G469), .B(new_n743), .C1(new_n744), .C2(KEYINPUT45), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n713), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n665), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n745), .B2(new_n713), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n585), .B(new_n641), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n600), .A2(new_n582), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT111), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n594), .A2(new_n624), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n749), .B1(new_n757), .B2(KEYINPUT44), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n730), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  NOR3_X1   g576(.A1(new_n730), .A2(new_n658), .A3(new_n440), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n486), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n764), .B1(new_n763), .B2(new_n486), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n747), .A2(new_n748), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(KEYINPUT47), .A3(new_n585), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT47), .B1(new_n768), .B2(new_n585), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n765), .B(new_n767), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  NOR2_X1   g587(.A1(new_n640), .A2(new_n486), .ZN(new_n774));
  INV_X1    g588(.A(new_n651), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n750), .A2(new_n301), .A3(new_n603), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n668), .A2(new_n669), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT49), .Z(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n640), .A2(new_n187), .A3(new_n670), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT116), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n487), .A2(new_n752), .A3(new_n563), .A4(new_n690), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT50), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n730), .A2(new_n670), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n487), .A2(new_n786), .A3(new_n563), .A4(new_n775), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n600), .A3(new_n581), .A4(new_n580), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n768), .A2(new_n585), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n769), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n777), .A2(new_n585), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n712), .B(new_n782), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n752), .A2(new_n563), .A3(new_n709), .A4(new_n786), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n785), .A2(KEYINPUT51), .A3(new_n788), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n788), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n799), .B2(new_n784), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n371), .A2(new_n440), .ZN(new_n802));
  INV_X1    g616(.A(new_n624), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n802), .A2(new_n297), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n804), .A2(new_n636), .B1(new_n700), .B2(new_n709), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n717), .A2(new_n651), .A3(new_n803), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n609), .A3(new_n657), .A4(new_n646), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n660), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n710), .A2(new_n637), .A3(new_n660), .A4(new_n807), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n720), .A2(new_n733), .B1(new_n737), .B2(new_n740), .ZN(new_n813));
  INV_X1    g627(.A(new_n583), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n707), .B1(new_n690), .B2(new_n624), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n814), .B(new_n717), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n803), .A2(new_n557), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n630), .A2(new_n600), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n657), .A3(new_n712), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n672), .A2(new_n682), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n679), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n813), .A2(new_n821), .A3(new_n698), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n812), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n600), .A2(new_n557), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n297), .A2(KEYINPUT87), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n297), .A2(KEYINPUT87), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n568), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n298), .A2(new_n831), .A3(new_n568), .A4(new_n826), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n832), .A3(new_n595), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n568), .B(new_n814), .C1(new_n827), .C2(new_n828), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n298), .A2(new_n836), .A3(new_n568), .A4(new_n814), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n837), .A3(new_n595), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n571), .A2(new_n833), .A3(new_n838), .A4(new_n626), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n825), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n734), .A2(new_n741), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n635), .B(new_n730), .C1(new_n817), .C2(new_n819), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n808), .A2(new_n811), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n823), .A2(new_n698), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n833), .A2(new_n838), .A3(new_n571), .A4(new_n626), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT54), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n782), .A2(new_n693), .ZN(new_n851));
  INV_X1    g665(.A(new_n824), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n839), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n844), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n729), .A2(new_n487), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n563), .A3(new_n752), .A4(new_n786), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT48), .Z(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n562), .A3(G953), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n850), .A2(new_n851), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n787), .A2(new_n814), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n801), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(G952), .A2(G953), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n779), .B1(new_n863), .B2(new_n864), .ZN(G75));
  XNOR2_X1  g679(.A(new_n278), .B(KEYINPUT117), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(G210), .B(G902), .C1(new_n840), .C2(new_n849), .ZN(new_n869));
  NOR2_X1   g683(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n869), .A2(new_n224), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n224), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n870), .ZN(new_n874));
  INV_X1    g688(.A(new_n224), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n869), .A2(new_n224), .A3(new_n870), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n867), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n219), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n873), .A2(new_n878), .A3(new_n880), .ZN(G51));
  XOR2_X1   g695(.A(new_n713), .B(KEYINPUT57), .Z(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n850), .B2(new_n856), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n856), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n367), .A2(new_n368), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n282), .B1(new_n853), .B2(new_n854), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(new_n745), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n879), .B1(new_n888), .B2(new_n891), .ZN(G54));
  NAND3_X1  g706(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n893));
  INV_X1    g707(.A(new_n515), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .A4(new_n515), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n880), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n899), .A3(new_n880), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(G60));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n850), .B2(new_n856), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n576), .A2(new_n578), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n880), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n884), .A2(new_n885), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n903), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n905), .ZN(G63));
  NAND2_X1  g723(.A1(new_n853), .A2(new_n854), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n474), .A2(new_n282), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n622), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n913), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n853), .B2(new_n854), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n914), .B(new_n880), .C1(new_n473), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT61), .B1(new_n917), .B2(KEYINPUT121), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G66));
  AOI21_X1  g735(.A(new_n219), .B1(new_n567), .B2(G224), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n823), .A2(new_n698), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n848), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT123), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n922), .B1(new_n926), .B2(new_n219), .ZN(new_n927));
  INV_X1    g741(.A(G898), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n866), .B1(new_n928), .B2(G953), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G69));
  INV_X1    g744(.A(new_n749), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(new_n609), .A3(new_n646), .A4(new_n857), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n932), .A2(new_n813), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n772), .A3(new_n761), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n805), .A2(new_n660), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT125), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n766), .B1(new_n791), .B2(new_n769), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n937), .A2(new_n765), .B1(new_n758), .B2(new_n760), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n939));
  INV_X1    g753(.A(new_n935), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n938), .A2(new_n933), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n405), .A2(new_n406), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n508), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n219), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(G227), .A2(G900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G953), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n640), .A2(new_n644), .ZN(new_n948));
  INV_X1    g762(.A(new_n652), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n643), .A4(new_n653), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n940), .A2(new_n950), .A3(KEYINPUT62), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n655), .B2(new_n935), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n591), .A2(new_n642), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n738), .B(new_n955), .C1(new_n814), .C2(new_n826), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n938), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n938), .A2(new_n954), .A3(KEYINPUT124), .A4(new_n956), .ZN(new_n960));
  AOI21_X1  g774(.A(G953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n945), .B(new_n947), .C1(new_n961), .C2(new_n944), .ZN(new_n962));
  XOR2_X1   g776(.A(KEYINPUT126), .B(G900), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n944), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(G953), .A3(new_n946), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n962), .A2(KEYINPUT127), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n434), .B1(new_n421), .B2(new_n378), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n910), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n972), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n959), .A2(new_n960), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n925), .ZN(new_n977));
  INV_X1    g791(.A(new_n421), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n378), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n880), .B(new_n974), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n925), .A2(new_n941), .A3(new_n936), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n378), .B(new_n978), .C1(new_n981), .C2(new_n972), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n982), .ZN(G57));
endmodule


