

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739;

  NOR2_X1 U367 ( .A1(n562), .A2(n690), .ZN(n533) );
  AND2_X1 U368 ( .A1(n365), .A2(n505), .ZN(n499) );
  XNOR2_X1 U369 ( .A(n503), .B(KEYINPUT106), .ZN(n562) );
  INV_X1 U370 ( .A(n670), .ZN(n509) );
  OR2_X1 U371 ( .A1(n660), .A2(G902), .ZN(n404) );
  OR2_X1 U372 ( .A1(n546), .A2(n690), .ZN(n583) );
  XNOR2_X1 U373 ( .A(n394), .B(KEYINPUT64), .ZN(n395) );
  XNOR2_X2 U374 ( .A(n344), .B(n553), .ZN(n652) );
  NAND2_X2 U375 ( .A1(n550), .A2(n549), .ZN(n344) );
  BUF_X2 U376 ( .A(n623), .Z(n666) );
  NAND2_X1 U377 ( .A1(n350), .A2(n366), .ZN(n370) );
  XNOR2_X1 U378 ( .A(G128), .B(G110), .ZN(n405) );
  NOR2_X1 U379 ( .A1(n556), .A2(n687), .ZN(n558) );
  INV_X2 U380 ( .A(G953), .ZN(n733) );
  XNOR2_X1 U381 ( .A(n377), .B(KEYINPUT32), .ZN(n651) );
  AND2_X4 U382 ( .A1(n604), .A2(n352), .ZN(n346) );
  XNOR2_X2 U383 ( .A(n395), .B(n476), .ZN(n444) );
  XNOR2_X1 U384 ( .A(n370), .B(KEYINPUT35), .ZN(n525) );
  INV_X1 U385 ( .A(n506), .ZN(n512) );
  NAND2_X1 U386 ( .A1(n505), .A2(n504), .ZN(n681) );
  OR2_X1 U387 ( .A1(n494), .A2(n493), .ZN(n377) );
  XNOR2_X1 U388 ( .A(n378), .B(n492), .ZN(n494) );
  OR2_X1 U389 ( .A1(n696), .A2(n501), .ZN(n369) );
  XNOR2_X1 U390 ( .A(n449), .B(n448), .ZN(n546) );
  XNOR2_X2 U391 ( .A(G101), .B(KEYINPUT67), .ZN(n423) );
  XNOR2_X1 U392 ( .A(G143), .B(G128), .ZN(n476) );
  BUF_X1 U393 ( .A(n562), .Z(n345) );
  NAND2_X1 U394 ( .A1(n346), .A2(G217), .ZN(n648) );
  NAND2_X1 U395 ( .A1(n346), .A2(G210), .ZN(n609) );
  NAND2_X1 U396 ( .A1(n346), .A2(G475), .ZN(n638) );
  NAND2_X1 U397 ( .A1(n346), .A2(G472), .ZN(n644) );
  NAND2_X1 U398 ( .A1(n346), .A2(G478), .ZN(n657) );
  NAND2_X1 U399 ( .A1(n346), .A2(G469), .ZN(n663) );
  XNOR2_X2 U400 ( .A(n347), .B(n348), .ZN(n503) );
  NOR2_X1 U401 ( .A1(n642), .A2(G902), .ZN(n347) );
  XOR2_X1 U402 ( .A(n434), .B(n433), .Z(n348) );
  AND2_X2 U403 ( .A1(n369), .A2(n368), .ZN(n350) );
  XNOR2_X2 U404 ( .A(n730), .B(G146), .ZN(n432) );
  XNOR2_X2 U405 ( .A(n444), .B(n396), .ZN(n730) );
  NAND2_X1 U406 ( .A1(n491), .A2(n349), .ZN(n378) );
  AND2_X1 U407 ( .A1(n581), .A2(n509), .ZN(n365) );
  AND2_X1 U408 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U409 ( .A1(KEYINPUT80), .A2(G953), .ZN(n388) );
  NAND2_X1 U410 ( .A1(n390), .A2(KEYINPUT80), .ZN(n389) );
  INV_X1 U411 ( .A(G224), .ZN(n390) );
  NAND2_X1 U412 ( .A1(n385), .A2(n733), .ZN(n384) );
  AND2_X1 U413 ( .A1(n386), .A2(G224), .ZN(n385) );
  XNOR2_X1 U414 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n440) );
  XNOR2_X1 U415 ( .A(G110), .B(KEYINPUT16), .ZN(n436) );
  NOR2_X1 U416 ( .A1(n391), .A2(n372), .ZN(n363) );
  BUF_X1 U417 ( .A(n546), .Z(n598) );
  XNOR2_X1 U418 ( .A(n545), .B(n544), .ZN(n570) );
  XNOR2_X1 U419 ( .A(n471), .B(G475), .ZN(n472) );
  INV_X1 U420 ( .A(KEYINPUT46), .ZN(n376) );
  XNOR2_X2 U421 ( .A(G119), .B(G113), .ZN(n424) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n459) );
  XNOR2_X1 U423 ( .A(G113), .B(G143), .ZN(n461) );
  NAND2_X1 U424 ( .A1(n532), .A2(KEYINPUT2), .ZN(n392) );
  XNOR2_X1 U425 ( .A(n499), .B(n354), .ZN(n696) );
  XNOR2_X1 U426 ( .A(n598), .B(n547), .ZN(n555) );
  BUF_X1 U427 ( .A(n503), .Z(n510) );
  XNOR2_X1 U428 ( .A(G107), .B(G110), .ZN(n400) );
  NAND2_X1 U429 ( .A1(n387), .A2(n384), .ZN(n442) );
  BUF_X1 U430 ( .A(n696), .Z(n705) );
  XNOR2_X1 U431 ( .A(n373), .B(n356), .ZN(n358) );
  XNOR2_X1 U432 ( .A(n610), .B(KEYINPUT91), .ZN(n658) );
  XNOR2_X1 U433 ( .A(n566), .B(KEYINPUT42), .ZN(n621) );
  NAND2_X1 U434 ( .A1(n588), .A2(n505), .ZN(n616) );
  OR2_X1 U435 ( .A1(n595), .A2(n583), .ZN(n587) );
  BUF_X1 U436 ( .A(n525), .Z(n654) );
  AND2_X1 U437 ( .A1(n570), .A2(n569), .ZN(n635) );
  INV_X1 U438 ( .A(n505), .ZN(n672) );
  NAND2_X2 U439 ( .A1(n358), .A2(n600), .ZN(n602) );
  AND2_X1 U440 ( .A1(n693), .A2(n559), .ZN(n349) );
  AND2_X1 U441 ( .A1(n512), .A2(n501), .ZN(n351) );
  OR2_X1 U442 ( .A1(n603), .A2(n602), .ZN(n352) );
  AND2_X1 U443 ( .A1(n523), .A2(n622), .ZN(n353) );
  XOR2_X1 U444 ( .A(n498), .B(KEYINPUT33), .Z(n354) );
  XOR2_X1 U445 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n355) );
  INV_X1 U446 ( .A(n725), .ZN(n549) );
  INV_X1 U447 ( .A(n727), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n593), .B(KEYINPUT48), .ZN(n356) );
  AND2_X1 U449 ( .A1(n532), .A2(KEYINPUT84), .ZN(n357) );
  XNOR2_X2 U450 ( .A(n602), .B(KEYINPUT75), .ZN(n364) );
  NAND2_X1 U451 ( .A1(n361), .A2(n359), .ZN(n604) );
  NAND2_X1 U452 ( .A1(n364), .A2(n360), .ZN(n359) );
  AND2_X1 U453 ( .A1(n666), .A2(n357), .ZN(n360) );
  XNOR2_X2 U454 ( .A(n531), .B(n530), .ZN(n623) );
  NAND2_X1 U455 ( .A1(n362), .A2(n371), .ZN(n361) );
  NAND2_X1 U456 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X2 U457 ( .A(n571), .B(KEYINPUT1), .ZN(n505) );
  XNOR2_X2 U458 ( .A(n404), .B(G469), .ZN(n571) );
  XNOR2_X2 U459 ( .A(n503), .B(KEYINPUT6), .ZN(n581) );
  NOR2_X1 U460 ( .A1(n367), .A2(n568), .ZN(n366) );
  NOR2_X1 U461 ( .A1(n512), .A2(n501), .ZN(n367) );
  NAND2_X1 U462 ( .A1(n696), .A2(n351), .ZN(n368) );
  NAND2_X1 U463 ( .A1(n392), .A2(KEYINPUT84), .ZN(n371) );
  INV_X1 U464 ( .A(n392), .ZN(n372) );
  NAND2_X1 U465 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U466 ( .A1(n592), .A2(n591), .ZN(n374) );
  XNOR2_X1 U467 ( .A(n567), .B(n376), .ZN(n375) );
  NAND2_X1 U468 ( .A1(n572), .A2(n457), .ZN(n458) );
  XNOR2_X2 U469 ( .A(n583), .B(KEYINPUT19), .ZN(n572) );
  NAND2_X1 U470 ( .A1(n380), .A2(n379), .ZN(n382) );
  INV_X1 U471 ( .A(n524), .ZN(n379) );
  INV_X1 U472 ( .A(n525), .ZN(n380) );
  NAND2_X1 U473 ( .A1(n381), .A2(n353), .ZN(n383) );
  NAND2_X1 U474 ( .A1(n382), .A2(KEYINPUT44), .ZN(n381) );
  XNOR2_X1 U475 ( .A(n383), .B(KEYINPUT89), .ZN(n529) );
  INV_X1 U476 ( .A(KEYINPUT80), .ZN(n386) );
  NAND2_X1 U477 ( .A1(n623), .A2(n532), .ZN(n391) );
  NAND2_X1 U478 ( .A1(n550), .A2(n393), .ZN(n634) );
  XNOR2_X2 U479 ( .A(n548), .B(n355), .ZN(n550) );
  INV_X1 U480 ( .A(KEYINPUT99), .ZN(n513) );
  XNOR2_X1 U481 ( .A(n514), .B(n513), .ZN(n517) );
  NAND2_X1 U482 ( .A1(n517), .A2(n686), .ZN(n523) );
  XNOR2_X1 U483 ( .A(n467), .B(n466), .ZN(n470) );
  XNOR2_X1 U484 ( .A(n473), .B(n472), .ZN(n516) );
  XNOR2_X2 U485 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n394) );
  INV_X1 U486 ( .A(G137), .ZN(n411) );
  XNOR2_X1 U487 ( .A(n411), .B(G134), .ZN(n396) );
  NAND2_X1 U488 ( .A1(n733), .A2(G227), .ZN(n397) );
  XNOR2_X1 U489 ( .A(n397), .B(KEYINPUT79), .ZN(n398) );
  XNOR2_X1 U490 ( .A(G131), .B(G140), .ZN(n468) );
  XNOR2_X1 U491 ( .A(n398), .B(n468), .ZN(n402) );
  XNOR2_X1 U492 ( .A(G101), .B(G104), .ZN(n399) );
  XNOR2_X1 U493 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U494 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U495 ( .A(n432), .B(n403), .ZN(n660) );
  XNOR2_X1 U496 ( .A(n405), .B(KEYINPUT24), .ZN(n407) );
  XNOR2_X1 U497 ( .A(KEYINPUT96), .B(KEYINPUT23), .ZN(n406) );
  XNOR2_X1 U498 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X2 U499 ( .A(G146), .B(G125), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n441), .B(KEYINPUT10), .ZN(n469) );
  XNOR2_X1 U501 ( .A(n408), .B(n469), .ZN(n417) );
  NAND2_X1 U502 ( .A1(G234), .A2(n733), .ZN(n410) );
  INV_X1 U503 ( .A(KEYINPUT8), .ZN(n409) );
  XNOR2_X1 U504 ( .A(n410), .B(n409), .ZN(n474) );
  NAND2_X1 U505 ( .A1(n474), .A2(G221), .ZN(n415) );
  XNOR2_X1 U506 ( .A(n411), .B(G140), .ZN(n413) );
  XNOR2_X1 U507 ( .A(G119), .B(KEYINPUT68), .ZN(n412) );
  XNOR2_X1 U508 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U509 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U510 ( .A(n417), .B(n416), .ZN(n647) );
  INV_X1 U511 ( .A(G902), .ZN(n486) );
  NAND2_X1 U512 ( .A1(n647), .A2(n486), .ZN(n422) );
  XNOR2_X1 U513 ( .A(G902), .B(KEYINPUT15), .ZN(n601) );
  NAND2_X1 U514 ( .A1(n601), .A2(G234), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n418), .B(KEYINPUT20), .ZN(n489) );
  NAND2_X1 U516 ( .A1(n489), .A2(G217), .ZN(n420) );
  XNOR2_X1 U517 ( .A(KEYINPUT78), .B(KEYINPUT25), .ZN(n419) );
  XNOR2_X1 U518 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X2 U519 ( .A(n422), .B(n421), .ZN(n497) );
  NAND2_X1 U520 ( .A1(n505), .A2(n497), .ZN(n435) );
  XNOR2_X1 U521 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U522 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n425) );
  XNOR2_X1 U523 ( .A(n426), .B(n425), .ZN(n439) );
  NAND2_X1 U524 ( .A1(n459), .A2(G210), .ZN(n427) );
  XNOR2_X1 U525 ( .A(n427), .B(G131), .ZN(n429) );
  XNOR2_X1 U526 ( .A(G116), .B(KEYINPUT5), .ZN(n428) );
  XNOR2_X1 U527 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U528 ( .A(n439), .B(n430), .Z(n431) );
  XNOR2_X1 U529 ( .A(n432), .B(n431), .ZN(n642) );
  XNOR2_X1 U530 ( .A(G472), .B(KEYINPUT97), .ZN(n434) );
  INV_X1 U531 ( .A(KEYINPUT71), .ZN(n433) );
  OR2_X1 U532 ( .A1(n435), .A2(n581), .ZN(n493) );
  XNOR2_X2 U533 ( .A(G116), .B(G107), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(n436), .ZN(n437) );
  XNOR2_X1 U535 ( .A(G122), .B(G104), .ZN(n464) );
  XNOR2_X1 U536 ( .A(n437), .B(n464), .ZN(n438) );
  XNOR2_X1 U537 ( .A(n439), .B(n438), .ZN(n628) );
  XNOR2_X1 U538 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U539 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U540 ( .A(n444), .B(n445), .ZN(n446) );
  XNOR2_X1 U541 ( .A(n628), .B(n446), .ZN(n607) );
  INV_X1 U542 ( .A(n601), .ZN(n532) );
  OR2_X2 U543 ( .A1(n607), .A2(n532), .ZN(n449) );
  INV_X1 U544 ( .A(G237), .ZN(n447) );
  NAND2_X1 U545 ( .A1(n486), .A2(n447), .ZN(n450) );
  NAND2_X1 U546 ( .A1(n450), .A2(G210), .ZN(n448) );
  AND2_X1 U547 ( .A1(n450), .A2(G214), .ZN(n690) );
  NAND2_X1 U548 ( .A1(G237), .A2(G234), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n451), .B(KEYINPUT14), .ZN(n455) );
  NAND2_X1 U550 ( .A1(G952), .A2(n455), .ZN(n452) );
  XOR2_X1 U551 ( .A(KEYINPUT93), .B(n452), .Z(n702) );
  NOR2_X1 U552 ( .A1(n702), .A2(G953), .ZN(n453) );
  XNOR2_X1 U553 ( .A(n453), .B(KEYINPUT94), .ZN(n539) );
  NOR2_X1 U554 ( .A1(G898), .A2(n733), .ZN(n454) );
  XNOR2_X1 U555 ( .A(KEYINPUT95), .B(n454), .ZN(n629) );
  NAND2_X1 U556 ( .A1(G902), .A2(n455), .ZN(n535) );
  NOR2_X1 U557 ( .A1(n629), .A2(n535), .ZN(n456) );
  OR2_X1 U558 ( .A1(n539), .A2(n456), .ZN(n457) );
  XNOR2_X1 U559 ( .A(n458), .B(KEYINPUT0), .ZN(n500) );
  INV_X1 U560 ( .A(n500), .ZN(n491) );
  NAND2_X1 U561 ( .A1(n459), .A2(G214), .ZN(n460) );
  XOR2_X1 U562 ( .A(n461), .B(n460), .Z(n467) );
  XOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n463) );
  XNOR2_X1 U564 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n462) );
  XNOR2_X1 U565 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U566 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n469), .B(n468), .ZN(n731) );
  XNOR2_X1 U568 ( .A(n470), .B(n731), .ZN(n636) );
  NOR2_X1 U569 ( .A1(G902), .A2(n636), .ZN(n473) );
  XNOR2_X1 U570 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n471) );
  NAND2_X1 U571 ( .A1(n474), .A2(G217), .ZN(n478) );
  XNOR2_X1 U572 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U573 ( .A(n478), .B(n477), .ZN(n485) );
  XOR2_X1 U574 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n480) );
  XNOR2_X1 U575 ( .A(G134), .B(KEYINPUT7), .ZN(n479) );
  XNOR2_X1 U576 ( .A(n480), .B(n479), .ZN(n483) );
  XNOR2_X1 U577 ( .A(G122), .B(KEYINPUT105), .ZN(n481) );
  XNOR2_X1 U578 ( .A(n481), .B(KEYINPUT103), .ZN(n482) );
  XNOR2_X1 U579 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U580 ( .A(n485), .B(n484), .ZN(n655) );
  NAND2_X1 U581 ( .A1(n655), .A2(n486), .ZN(n488) );
  INV_X1 U582 ( .A(G478), .ZN(n487) );
  XNOR2_X1 U583 ( .A(n488), .B(n487), .ZN(n515) );
  INV_X1 U584 ( .A(n515), .ZN(n502) );
  NOR2_X1 U585 ( .A1(n516), .A2(n502), .ZN(n693) );
  NAND2_X1 U586 ( .A1(n489), .A2(G221), .ZN(n490) );
  XNOR2_X1 U587 ( .A(n490), .B(KEYINPUT21), .ZN(n675) );
  INV_X1 U588 ( .A(n675), .ZN(n559) );
  XNOR2_X1 U589 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n492) );
  INV_X1 U590 ( .A(n494), .ZN(n519) );
  NAND2_X1 U591 ( .A1(n345), .A2(n497), .ZN(n495) );
  NOR2_X1 U592 ( .A1(n495), .A2(n505), .ZN(n496) );
  NAND2_X1 U593 ( .A1(n519), .A2(n496), .ZN(n618) );
  NAND2_X1 U594 ( .A1(n651), .A2(n618), .ZN(n524) );
  OR2_X1 U595 ( .A1(n497), .A2(n675), .ZN(n670) );
  INV_X1 U596 ( .A(KEYINPUT69), .ZN(n498) );
  BUF_X1 U597 ( .A(n500), .Z(n506) );
  XOR2_X1 U598 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n501) );
  NAND2_X1 U599 ( .A1(n516), .A2(n502), .ZN(n568) );
  XOR2_X1 U600 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n508) );
  NOR2_X1 U601 ( .A1(n510), .A2(n670), .ZN(n504) );
  NOR2_X2 U602 ( .A1(n506), .A2(n681), .ZN(n507) );
  XOR2_X2 U603 ( .A(n508), .B(n507), .Z(n728) );
  NAND2_X1 U604 ( .A1(n571), .A2(n509), .ZN(n534) );
  INV_X1 U605 ( .A(n510), .ZN(n678) );
  NOR2_X1 U606 ( .A1(n534), .A2(n678), .ZN(n511) );
  NAND2_X1 U607 ( .A1(n512), .A2(n511), .ZN(n715) );
  NAND2_X1 U608 ( .A1(n728), .A2(n715), .ZN(n514) );
  OR2_X1 U609 ( .A1(n516), .A2(n515), .ZN(n727) );
  NAND2_X1 U610 ( .A1(n516), .A2(n515), .ZN(n725) );
  NAND2_X1 U611 ( .A1(n727), .A2(n725), .ZN(n686) );
  INV_X1 U612 ( .A(n581), .ZN(n518) );
  NAND2_X1 U613 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U614 ( .A(KEYINPUT88), .B(n520), .Z(n522) );
  NOR2_X1 U615 ( .A1(n505), .A2(n497), .ZN(n521) );
  NAND2_X1 U616 ( .A1(n522), .A2(n521), .ZN(n622) );
  NOR2_X1 U617 ( .A1(n524), .A2(KEYINPUT44), .ZN(n527) );
  INV_X1 U618 ( .A(n654), .ZN(n526) );
  NAND2_X1 U619 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U620 ( .A1(n529), .A2(n528), .ZN(n531) );
  XOR2_X1 U621 ( .A(KEYINPUT85), .B(KEYINPUT45), .Z(n530) );
  XNOR2_X1 U622 ( .A(n533), .B(KEYINPUT30), .ZN(n543) );
  INV_X1 U623 ( .A(n534), .ZN(n540) );
  NOR2_X1 U624 ( .A1(G900), .A2(n535), .ZN(n536) );
  NAND2_X1 U625 ( .A1(G953), .A2(n536), .ZN(n537) );
  XNOR2_X1 U626 ( .A(n537), .B(KEYINPUT107), .ZN(n538) );
  OR2_X1 U627 ( .A1(n539), .A2(n538), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n540), .A2(n560), .ZN(n541) );
  XNOR2_X1 U629 ( .A(n541), .B(KEYINPUT77), .ZN(n542) );
  NAND2_X1 U630 ( .A1(n543), .A2(n542), .ZN(n545) );
  INV_X1 U631 ( .A(KEYINPUT76), .ZN(n544) );
  XNOR2_X1 U632 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n547) );
  NAND2_X1 U633 ( .A1(n570), .A2(n555), .ZN(n548) );
  XNOR2_X1 U634 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n552) );
  INV_X1 U635 ( .A(KEYINPUT110), .ZN(n551) );
  XNOR2_X1 U636 ( .A(n552), .B(n551), .ZN(n553) );
  INV_X1 U637 ( .A(n693), .ZN(n556) );
  INV_X1 U638 ( .A(n555), .ZN(n691) );
  OR2_X1 U639 ( .A1(n691), .A2(n690), .ZN(n687) );
  INV_X1 U640 ( .A(KEYINPUT41), .ZN(n557) );
  XNOR2_X1 U641 ( .A(n558), .B(n557), .ZN(n704) );
  AND2_X1 U642 ( .A1(n704), .A2(n571), .ZN(n565) );
  AND2_X1 U643 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n497), .A2(n561), .ZN(n580) );
  OR2_X1 U645 ( .A1(n345), .A2(n580), .ZN(n564) );
  XNOR2_X1 U646 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n564), .B(n563), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n565), .A2(n574), .ZN(n566) );
  NAND2_X1 U649 ( .A1(n652), .A2(n621), .ZN(n567) );
  NOR2_X1 U650 ( .A1(n568), .A2(n598), .ZN(n569) );
  XNOR2_X1 U651 ( .A(n635), .B(KEYINPUT83), .ZN(n576) );
  AND2_X1 U652 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U653 ( .A1(n574), .A2(n573), .ZN(n722) );
  NAND2_X1 U654 ( .A1(n722), .A2(n686), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n578), .A2(KEYINPUT47), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U657 ( .A(n577), .B(KEYINPUT82), .ZN(n592) );
  NOR2_X1 U658 ( .A1(n578), .A2(KEYINPUT47), .ZN(n579) );
  XNOR2_X1 U659 ( .A(n579), .B(KEYINPUT73), .ZN(n590) );
  NOR2_X1 U660 ( .A1(n725), .A2(n580), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n595) );
  XNOR2_X1 U662 ( .A(KEYINPUT112), .B(KEYINPUT36), .ZN(n585) );
  INV_X1 U663 ( .A(KEYINPUT90), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U665 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n616), .B(KEYINPUT86), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U668 ( .A(KEYINPUT66), .ZN(n593) );
  OR2_X1 U669 ( .A1(n505), .A2(n690), .ZN(n594) );
  OR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U671 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n597), .B(n596), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n620) );
  AND2_X1 U674 ( .A1(n634), .A2(n620), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n623), .A2(KEYINPUT2), .ZN(n603) );
  XOR2_X1 U676 ( .A(KEYINPUT81), .B(KEYINPUT54), .Z(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT55), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n609), .B(n608), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n733), .A2(G952), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n658), .ZN(n613) );
  INV_X1 U682 ( .A(KEYINPUT56), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(G51) );
  XNOR2_X1 U684 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(G125), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(G27) );
  XNOR2_X1 U687 ( .A(G110), .B(KEYINPUT114), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(G12) );
  XNOR2_X1 U689 ( .A(G140), .B(KEYINPUT118), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(G42) );
  XNOR2_X1 U691 ( .A(n621), .B(G137), .ZN(G39) );
  XNOR2_X1 U692 ( .A(n622), .B(G101), .ZN(G3) );
  NAND2_X1 U693 ( .A1(n666), .A2(n733), .ZN(n627) );
  NAND2_X1 U694 ( .A1(G953), .A2(G224), .ZN(n624) );
  XNOR2_X1 U695 ( .A(KEYINPUT61), .B(n624), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n625), .A2(G898), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n633) );
  INV_X1 U698 ( .A(n628), .ZN(n631) );
  INV_X1 U699 ( .A(n629), .ZN(n630) );
  NOR2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U701 ( .A(n633), .B(n632), .ZN(G69) );
  XNOR2_X1 U702 ( .A(n634), .B(G134), .ZN(G36) );
  XOR2_X1 U703 ( .A(G143), .B(n635), .Z(G45) );
  XNOR2_X1 U704 ( .A(n636), .B(KEYINPUT59), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n639), .A2(n658), .ZN(n641) );
  XNOR2_X1 U707 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(G60) );
  XOR2_X1 U709 ( .A(KEYINPUT62), .B(n642), .Z(n643) );
  XNOR2_X1 U710 ( .A(n644), .B(n643), .ZN(n645) );
  NAND2_X1 U711 ( .A1(n645), .A2(n658), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n646), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U713 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n649), .A2(n658), .ZN(n650) );
  XNOR2_X1 U715 ( .A(n650), .B(KEYINPUT125), .ZN(G66) );
  XNOR2_X1 U716 ( .A(n651), .B(G119), .ZN(G21) );
  XNOR2_X1 U717 ( .A(n652), .B(G131), .ZN(G33) );
  XNOR2_X1 U718 ( .A(G122), .B(KEYINPUT127), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n654), .B(n653), .ZN(G24) );
  XOR2_X1 U720 ( .A(KEYINPUT124), .B(n655), .Z(n656) );
  XNOR2_X1 U721 ( .A(n657), .B(n656), .ZN(n659) );
  INV_X1 U722 ( .A(n658), .ZN(n664) );
  NOR2_X1 U723 ( .A1(n659), .A2(n664), .ZN(G63) );
  XOR2_X1 U724 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n661) );
  XNOR2_X1 U725 ( .A(n660), .B(n661), .ZN(n662) );
  XNOR2_X1 U726 ( .A(n663), .B(n662), .ZN(n665) );
  NOR2_X1 U727 ( .A1(n665), .A2(n664), .ZN(G54) );
  INV_X1 U728 ( .A(n666), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n667), .A2(n602), .ZN(n668) );
  XNOR2_X1 U730 ( .A(n668), .B(KEYINPUT2), .ZN(n710) );
  NAND2_X1 U731 ( .A1(n672), .A2(n670), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n669), .A2(KEYINPUT50), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n509), .A2(KEYINPUT50), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n680) );
  NAND2_X1 U736 ( .A1(n497), .A2(n675), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n676), .B(KEYINPUT49), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n682) );
  AND2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(n683), .Z(n684) );
  XNOR2_X1 U742 ( .A(KEYINPUT119), .B(n684), .ZN(n685) );
  NAND2_X1 U743 ( .A1(n685), .A2(n704), .ZN(n699) );
  INV_X1 U744 ( .A(n686), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U746 ( .A(KEYINPUT120), .B(n689), .Z(n695) );
  NAND2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U750 ( .A1(n697), .A2(n705), .ZN(n698) );
  NAND2_X1 U751 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U752 ( .A(KEYINPUT52), .B(n700), .Z(n701) );
  NOR2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U754 ( .A(KEYINPUT121), .B(n703), .Z(n708) );
  NAND2_X1 U755 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U756 ( .A1(n706), .A2(n733), .ZN(n707) );
  NOR2_X1 U757 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U758 ( .A1(n710), .A2(n709), .ZN(n712) );
  XOR2_X1 U759 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n711) );
  XNOR2_X1 U760 ( .A(n712), .B(n711), .ZN(G75) );
  NOR2_X1 U761 ( .A1(n715), .A2(n725), .ZN(n714) );
  XNOR2_X1 U762 ( .A(G104), .B(KEYINPUT113), .ZN(n713) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(G6) );
  NOR2_X1 U764 ( .A1(n715), .A2(n727), .ZN(n717) );
  XNOR2_X1 U765 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n716) );
  XNOR2_X1 U766 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U767 ( .A(G107), .B(n718), .ZN(G9) );
  NAND2_X1 U768 ( .A1(n722), .A2(n393), .ZN(n720) );
  XOR2_X1 U769 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U771 ( .A(G128), .B(n721), .Z(G30) );
  NAND2_X1 U772 ( .A1(n722), .A2(n549), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n723), .B(KEYINPUT116), .ZN(n724) );
  XNOR2_X1 U774 ( .A(G146), .B(n724), .ZN(G48) );
  NOR2_X1 U775 ( .A1(n728), .A2(n725), .ZN(n726) );
  XOR2_X1 U776 ( .A(G113), .B(n726), .Z(G15) );
  NOR2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U778 ( .A(G116), .B(n729), .Z(G18) );
  XNOR2_X1 U779 ( .A(n731), .B(KEYINPUT126), .ZN(n732) );
  XOR2_X1 U780 ( .A(n730), .B(n732), .Z(n735) );
  XNOR2_X1 U781 ( .A(n602), .B(n735), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n739) );
  XNOR2_X1 U783 ( .A(n735), .B(G227), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(G953), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(G72) );
endmodule

