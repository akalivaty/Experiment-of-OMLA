//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n203), .B1(G155gat), .B2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n202), .A2(new_n204), .B1(KEYINPUT74), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G155gat), .B(G162gat), .Z(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G113gat), .B(G120gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT4), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n216), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n208), .B(new_n209), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT4), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n216), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT5), .ZN(new_n228));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n227), .A2(KEYINPUT76), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n222), .A2(new_n229), .A3(new_n226), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT5), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n212), .B(new_n216), .ZN(new_n235));
  INV_X1    g034(.A(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(KEYINPUT5), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT83), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT83), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n241), .A3(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT75), .B(KEYINPUT0), .Z(new_n244));
  XNOR2_X1  g043(.A(G1gat), .B(G29gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G57gat), .B(G85gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT79), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n222), .A2(new_n226), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT80), .B(KEYINPUT39), .Z(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n236), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n249), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT81), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n236), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(KEYINPUT39), .C1(new_n236), .C2(new_n235), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n256), .A2(KEYINPUT81), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n252), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT40), .ZN(new_n263));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264));
  INV_X1    g063(.A(G211gat), .ZN(new_n265));
  INV_X1    g064(.A(G218gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(KEYINPUT22), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT71), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT27), .B(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  OR2_X1    g078(.A1(KEYINPUT65), .A2(KEYINPUT26), .ZN(new_n280));
  NAND2_X1  g079(.A1(KEYINPUT65), .A2(KEYINPUT26), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(new_n279), .B2(KEYINPUT26), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n283), .B(new_n284), .C1(new_n282), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n278), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n288), .A2(KEYINPUT64), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n290), .B1(new_n288), .B2(KEYINPUT64), .ZN(new_n292));
  NOR2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n284), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT25), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(new_n290), .B2(new_n288), .ZN(new_n302));
  OR3_X1    g101(.A1(new_n302), .A2(new_n298), .A3(KEYINPUT25), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n273), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n303), .A2(new_n299), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n272), .B1(new_n307), .B2(new_n289), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n270), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G92gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(G64gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n304), .A2(new_n273), .ZN(new_n315));
  INV_X1    g114(.A(new_n270), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n307), .B2(new_n289), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n273), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n309), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n305), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n272), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n323), .B2(new_n315), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n306), .A2(new_n308), .A3(new_n270), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n309), .A2(new_n318), .A3(KEYINPUT30), .A4(new_n314), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT40), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n252), .B(new_n329), .C1(new_n260), .C2(new_n261), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n251), .A2(new_n263), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT77), .A2(G22gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT31), .B(G50gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  MUX2_X1   g134(.A(G22gat), .B(new_n332), .S(new_n335), .Z(new_n336));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n337), .B(KEYINPUT78), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n336), .B(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT3), .B1(new_n316), .B2(new_n305), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n219), .B2(new_n224), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n340), .A2(new_n219), .B1(new_n316), .B2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n248), .B1(new_n234), .B2(new_n238), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT6), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n249), .B1(new_n240), .B2(new_n242), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n234), .A2(new_n248), .A3(new_n238), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT6), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n347), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT37), .B1(new_n324), .B2(new_n325), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT37), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n309), .A2(new_n354), .A3(new_n318), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n313), .A3(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n356), .A2(KEYINPUT38), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(KEYINPUT38), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n319), .A3(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n331), .B(new_n345), .C1(new_n352), .C2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n289), .A2(new_n218), .A3(new_n299), .A4(new_n303), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n307), .A2(KEYINPUT67), .A3(new_n218), .A4(new_n289), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n304), .A2(new_n216), .ZN(new_n365));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(KEYINPUT34), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(KEYINPUT34), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT69), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(KEYINPUT69), .A3(new_n369), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n374));
  XNOR2_X1  g173(.A(G15gat), .B(G43gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND3_X1  g176(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n378));
  INV_X1    g177(.A(new_n366), .ZN(new_n379));
  AOI221_X4 g178(.A(new_n374), .B1(KEYINPUT33), .B2(new_n377), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT33), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  INV_X1    g181(.A(new_n377), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n372), .B(new_n373), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  OR3_X1    g184(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n386));
  INV_X1    g185(.A(new_n380), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n386), .A2(new_n371), .A3(new_n370), .A4(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT36), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT70), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT68), .B1(new_n384), .B2(new_n380), .ZN(new_n393));
  INV_X1    g192(.A(new_n370), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT68), .B(new_n370), .C1(new_n384), .C2(new_n380), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(KEYINPUT36), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n385), .A2(new_n388), .A3(KEYINPUT70), .A4(new_n389), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n347), .B1(new_n351), .B2(new_n346), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n327), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n321), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT73), .B1(new_n326), .B2(new_n327), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n345), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n360), .A2(new_n399), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n395), .A2(new_n345), .A3(new_n396), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT35), .B1(new_n409), .B2(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n385), .B2(new_n388), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n328), .A2(KEYINPUT35), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n352), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(G43gat), .B(G50gat), .Z(new_n416));
  INV_X1    g215(.A(KEYINPUT15), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n418));
  NOR3_X1   g217(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n416), .A2(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT87), .ZN(new_n424));
  NAND2_X1  g223(.A1(G29gat), .A2(G36gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G43gat), .B(G50gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(KEYINPUT15), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT15), .B(new_n427), .C1(new_n423), .C2(new_n426), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G15gat), .B(G22gat), .Z(new_n434));
  INV_X1    g233(.A(G1gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G22gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n435), .A2(KEYINPUT88), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT16), .B1(new_n439), .B2(G1gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G8gat), .ZN(new_n444));
  INV_X1    g243(.A(G8gat), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n436), .A2(new_n441), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n429), .A2(KEYINPUT17), .A3(new_n430), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n431), .ZN(new_n451));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n449), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n454), .A2(new_n455), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n461));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n468));
  XNOR2_X1  g267(.A(G169gat), .B(G197gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n464), .B(new_n465), .ZN(new_n475));
  INV_X1    g274(.A(new_n470), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(KEYINPUT12), .A3(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n449), .A2(new_n458), .A3(new_n451), .A4(new_n456), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n452), .B(KEYINPUT13), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n451), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n450), .A2(new_n431), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n460), .A2(new_n479), .A3(new_n480), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n489), .B2(new_n451), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n457), .B2(new_n459), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n491), .A2(KEYINPUT91), .A3(new_n479), .A4(new_n480), .ZN(new_n492));
  INV_X1    g291(.A(new_n479), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n480), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n488), .A2(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT21), .ZN(new_n496));
  XNOR2_X1  g295(.A(G71gat), .B(G78gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n498));
  INV_X1    g297(.A(G64gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(G57gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(G57gat), .ZN(new_n501));
  INV_X1    g300(.A(G57gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G64gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n497), .B(new_n500), .C1(new_n504), .C2(new_n498), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT93), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n504), .A2(KEYINPUT9), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n505), .A2(new_n507), .B1(new_n508), .B2(new_n497), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n447), .B1(new_n496), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT95), .ZN(new_n511));
  XNOR2_X1  g310(.A(G127gat), .B(G155gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G231gat), .A2(G233gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(KEYINPUT94), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G183gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n265), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n513), .B(new_n517), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n496), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n518), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G134gat), .B(G162gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT41), .ZN(new_n524));
  INV_X1    g323(.A(G232gat), .ZN(new_n525));
  INV_X1    g324(.A(G233gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n523), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT100), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n530));
  XNOR2_X1  g329(.A(G99gat), .B(G106gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT96), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(G85gat), .A3(G92gat), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT7), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(KEYINPUT96), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT8), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n532), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT7), .ZN(new_n547));
  AOI22_X1  g346(.A1(KEYINPUT8), .A2(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n531), .A3(new_n539), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n530), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n530), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n431), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT98), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n557));
  INV_X1    g356(.A(new_n555), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n433), .B(new_n448), .C1(new_n550), .C2(new_n551), .ZN(new_n561));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT99), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n560), .B2(new_n561), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n529), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT100), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n528), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n571), .A3(new_n565), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n497), .B1(KEYINPUT9), .B2(new_n504), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT92), .ZN(new_n575));
  AND2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n500), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n506), .B(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n574), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n550), .A2(new_n551), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G230gat), .A2(G233gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n509), .B1(new_n549), .B2(new_n546), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT101), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n539), .A2(new_n541), .A3(new_n544), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n531), .B1(new_n588), .B2(new_n547), .ZN(new_n589));
  AND4_X1   g388(.A1(new_n531), .A2(new_n547), .A3(new_n539), .A4(new_n548), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT97), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n549), .A2(new_n530), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n509), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n582), .B1(new_n590), .B2(new_n589), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT10), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NOR4_X1   g395(.A1(new_n550), .A2(new_n551), .A3(new_n509), .A4(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n584), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n586), .A2(KEYINPUT101), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n587), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n522), .A2(new_n573), .A3(new_n607), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n415), .A2(new_n495), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n400), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT102), .B(G1gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(G1324gat));
  AND2_X1   g412(.A1(new_n609), .A2(new_n328), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT42), .B1(new_n614), .B2(new_n445), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  MUX2_X1   g416(.A(KEYINPUT42), .B(new_n615), .S(new_n617), .Z(G1325gat));
  NAND2_X1  g417(.A1(new_n385), .A2(new_n388), .ZN(new_n619));
  AOI21_X1  g418(.A(G15gat), .B1(new_n609), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n399), .B(KEYINPUT104), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n609), .A2(G15gat), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(G1326gat));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n406), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT105), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT43), .B(G22gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1327gat));
  NOR3_X1   g430(.A1(new_n522), .A2(new_n495), .A3(new_n606), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n415), .A2(new_n573), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G29gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n610), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT106), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT45), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT107), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n414), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n410), .A2(KEYINPUT107), .A3(new_n413), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n573), .B1(new_n642), .B2(new_n408), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT108), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT44), .B1(new_n415), .B2(new_n573), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n410), .A2(KEYINPUT107), .A3(new_n413), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT107), .B1(new_n410), .B2(new_n413), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n408), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n573), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n649), .A2(KEYINPUT108), .A3(new_n644), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n633), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n610), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n638), .B1(new_n635), .B2(new_n656), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n634), .A2(new_n658), .A3(new_n328), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT46), .Z(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(KEYINPUT109), .A3(new_n328), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(G36gat), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT109), .B1(new_n654), .B2(new_n328), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(G1329gat));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665));
  INV_X1    g464(.A(new_n399), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n666), .B(new_n632), .C1(new_n645), .C2(new_n652), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G43gat), .ZN(new_n668));
  AOI21_X1  g467(.A(G43gat), .B1(new_n385), .B2(new_n388), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n634), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n665), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n625), .B(new_n632), .C1(new_n645), .C2(new_n652), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(G43gat), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT110), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n667), .A2(G43gat), .B1(new_n634), .B2(new_n669), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n676), .B(new_n677), .C1(new_n665), .C2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n675), .A2(new_n679), .ZN(G1330gat));
  INV_X1    g479(.A(new_n653), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n406), .A3(new_n632), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G50gat), .ZN(new_n683));
  INV_X1    g482(.A(G50gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n634), .A2(new_n684), .A3(new_n406), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT48), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n683), .A2(KEYINPUT48), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1331gat));
  INV_X1    g489(.A(new_n522), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n488), .A2(new_n492), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n494), .A2(new_n493), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR4_X1   g493(.A1(new_n691), .A2(new_n694), .A3(new_n650), .A4(new_n607), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n649), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n400), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(new_n502), .ZN(G1332gat));
  NAND3_X1  g497(.A1(new_n649), .A2(new_n328), .A3(new_n695), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT49), .B(G64gat), .Z(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(G1333gat));
  OAI21_X1  g501(.A(G71gat), .B1(new_n696), .B2(new_n624), .ZN(new_n703));
  INV_X1    g502(.A(G71gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n619), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g506(.A1(new_n696), .A2(new_n345), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT111), .B(G78gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1335gat));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n495), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n607), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n681), .A2(new_n610), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G85gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n649), .A2(new_n650), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n715), .C2(new_n711), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n643), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n607), .B1(new_n721), .B2(KEYINPUT113), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(KEYINPUT113), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n610), .A2(new_n542), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n714), .B1(new_n723), .B2(new_n724), .ZN(G1336gat));
  NAND3_X1  g524(.A1(new_n681), .A2(new_n328), .A3(new_n712), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G92gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n721), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(new_n543), .A3(new_n328), .A4(new_n606), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT52), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1337gat));
  NAND3_X1  g533(.A1(new_n681), .A2(new_n625), .A3(new_n712), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT114), .B(G99gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n736), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n619), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n723), .B2(new_n739), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n681), .A2(new_n406), .A3(new_n712), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G106gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n345), .A2(G106gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n606), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n744), .B2(KEYINPUT115), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n742), .B(new_n744), .C1(KEYINPUT115), .C2(new_n746), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n605), .B1(new_n599), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n596), .B1(new_n583), .B2(new_n585), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n552), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n751), .B1(new_n756), .B2(new_n584), .ZN(new_n757));
  INV_X1    g556(.A(new_n584), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AND4_X1   g559(.A1(new_n753), .A2(new_n598), .A3(KEYINPUT54), .A4(new_n759), .ZN(new_n761));
  OAI211_X1 g560(.A(KEYINPUT55), .B(new_n752), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n601), .A2(new_n605), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n598), .A2(KEYINPUT54), .A3(new_n759), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n757), .A2(new_n753), .A3(new_n759), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT55), .B1(new_n768), .B2(new_n752), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n764), .A2(new_n769), .A3(new_n495), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n449), .A2(new_n451), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n453), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n489), .A2(new_n451), .A3(new_n481), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n472), .B(new_n473), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n488), .B2(new_n492), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n606), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n573), .B1(new_n770), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n568), .A3(new_n572), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n779), .A2(new_n764), .A3(new_n769), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(KEYINPUT117), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n752), .B1(new_n760), .B2(new_n761), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n694), .A3(new_n763), .A4(new_n762), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n650), .B1(new_n786), .B2(new_n776), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n779), .A2(new_n764), .A3(new_n769), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n781), .A2(new_n691), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n522), .A2(new_n495), .A3(new_n573), .A4(new_n607), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n400), .A2(new_n328), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(new_n411), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G113gat), .B1(new_n798), .B2(new_n495), .ZN(new_n799));
  INV_X1    g598(.A(new_n409), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n495), .A2(G113gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1340gat));
  OAI21_X1  g602(.A(G120gat), .B1(new_n798), .B2(new_n607), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n607), .A2(G120gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n801), .B2(new_n805), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n691), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n796), .A2(new_n800), .A3(new_n522), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n797), .A2(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1342gat));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n801), .A2(G134gat), .A3(new_n573), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n650), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(G134gat), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n812), .A2(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT119), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(KEYINPUT119), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(G1343gat));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n778), .A2(KEYINPUT120), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n780), .B1(new_n787), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n691), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n821), .B(new_n345), .C1(new_n825), .C2(new_n792), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n790), .A2(new_n792), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n406), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n830), .B2(new_n821), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n666), .A2(new_n795), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n831), .A2(new_n495), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(G141gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n820), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n793), .A2(new_n794), .A3(new_n345), .ZN(new_n839));
  INV_X1    g638(.A(new_n795), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n624), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(G141gat), .A3(new_n495), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n836), .B(new_n837), .C1(new_n838), .C2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n842), .ZN(new_n844));
  OAI221_X1 g643(.A(new_n844), .B1(new_n820), .B2(KEYINPUT58), .C1(new_n835), .C2(new_n834), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n830), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(new_n792), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n522), .B1(new_n778), .B2(new_n780), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n821), .B(new_n406), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n848), .A2(new_n606), .A3(new_n832), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G148gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n606), .B(new_n832), .C1(new_n854), .C2(new_n826), .ZN(new_n855));
  INV_X1    g654(.A(G148gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(KEYINPUT59), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n853), .A2(KEYINPUT59), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n841), .A2(G148gat), .A3(new_n607), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n847), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n859), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n855), .A2(new_n857), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n852), .B2(G148gat), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT122), .B(new_n861), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n865), .ZN(G1345gat));
  INV_X1    g665(.A(new_n841), .ZN(new_n867));
  AOI21_X1  g666(.A(G155gat), .B1(new_n867), .B2(new_n522), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n831), .A2(new_n833), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n691), .A2(new_n205), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(G1346gat));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n206), .A3(new_n650), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n831), .A2(new_n573), .A3(new_n833), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n206), .ZN(G1347gat));
  NAND2_X1  g673(.A1(new_n400), .A2(new_n328), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n793), .A2(new_n794), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n800), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(G169gat), .A3(new_n495), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT123), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n411), .ZN(new_n880));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n495), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1348gat));
  INV_X1    g681(.A(G176gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n880), .A2(new_n883), .A3(new_n607), .ZN(new_n884));
  INV_X1    g683(.A(new_n877), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n606), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n883), .B2(new_n886), .ZN(G1349gat));
  OAI21_X1  g686(.A(G183gat), .B1(new_n880), .B2(new_n691), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n522), .A2(new_n274), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n877), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n885), .A2(new_n275), .A3(new_n650), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n880), .A2(new_n573), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n275), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n894), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(G1351gat));
  NAND2_X1  g698(.A1(new_n839), .A2(new_n624), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n875), .ZN(new_n901));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n694), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n625), .A2(new_n875), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n851), .B(new_n904), .C1(new_n839), .C2(new_n821), .ZN(new_n905));
  OAI21_X1  g704(.A(G197gat), .B1(new_n905), .B2(new_n495), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(G1352gat));
  NOR2_X1   g706(.A1(new_n607), .A2(G204gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT124), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(KEYINPUT62), .A3(new_n912), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n848), .A2(new_n606), .A3(new_n851), .A4(new_n904), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G204gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(G1353gat));
  OAI211_X1 g718(.A(KEYINPUT63), .B(G211gat), .C1(new_n905), .C2(new_n691), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n922));
  OAI21_X1  g721(.A(G211gat), .B1(new_n905), .B2(new_n691), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n901), .A2(new_n265), .A3(new_n522), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1354gat));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n905), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n848), .A2(new_n931), .A3(new_n851), .A4(new_n904), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n650), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G218gat), .ZN(new_n934));
  NOR4_X1   g733(.A1(new_n900), .A2(G218gat), .A3(new_n573), .A4(new_n875), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n929), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT127), .B(new_n935), .C1(new_n933), .C2(G218gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(G1355gat));
endmodule


