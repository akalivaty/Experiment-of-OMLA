

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n522), .A2(G2104), .ZN(n897) );
  NOR2_X1 U552 ( .A1(n691), .A2(n690), .ZN(n694) );
  AND2_X1 U553 ( .A1(n994), .A2(n519), .ZN(n757) );
  XNOR2_X1 U554 ( .A(n711), .B(n710), .ZN(n716) );
  XNOR2_X1 U555 ( .A(n764), .B(KEYINPUT105), .ZN(n768) );
  NOR2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U557 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n520) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n522), .ZN(n532) );
  OR2_X1 U559 ( .A1(KEYINPUT33), .A2(n754), .ZN(n517) );
  OR2_X1 U560 ( .A1(n767), .A2(n766), .ZN(n518) );
  OR2_X1 U561 ( .A1(n756), .A2(n767), .ZN(n519) );
  XNOR2_X1 U562 ( .A(n731), .B(KEYINPUT98), .ZN(n688) );
  INV_X1 U563 ( .A(n688), .ZN(n712) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n710) );
  INV_X1 U565 ( .A(KEYINPUT31), .ZN(n727) );
  XNOR2_X1 U566 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U567 ( .A1(G2084), .A2(n731), .ZN(n717) );
  NAND2_X1 U568 ( .A1(n730), .A2(n729), .ZN(n741) );
  INV_X1 U569 ( .A(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U570 ( .A1(n789), .A2(n685), .ZN(n731) );
  AND2_X1 U571 ( .A1(n768), .A2(n518), .ZN(n802) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U573 ( .A1(G651), .A2(n638), .ZN(n652) );
  NAND2_X1 U574 ( .A1(n894), .A2(G138), .ZN(n536) );
  XNOR2_X1 U575 ( .A(n521), .B(n520), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U577 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U578 ( .A1(G101), .A2(n897), .ZN(n521) );
  NAND2_X1 U579 ( .A1(G125), .A2(n532), .ZN(n523) );
  XNOR2_X1 U580 ( .A(n523), .B(KEYINPUT64), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n525), .A2(n524), .ZN(n531) );
  XNOR2_X2 U582 ( .A(n527), .B(n526), .ZN(n894) );
  NAND2_X1 U583 ( .A1(G137), .A2(n894), .ZN(n529) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U585 ( .A1(G113), .A2(n890), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U587 ( .A1(G114), .A2(n890), .ZN(n534) );
  NAND2_X1 U588 ( .A1(G126), .A2(n532), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G102), .A2(n897), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U592 ( .A(KEYINPUT91), .B(n537), .Z(n538) );
  NOR2_X1 U593 ( .A1(n539), .A2(n538), .ZN(G164) );
  XOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .Z(n638) );
  NAND2_X1 U595 ( .A1(G50), .A2(n652), .ZN(n542) );
  INV_X1 U596 ( .A(G651), .ZN(n543) );
  NOR2_X1 U597 ( .A1(G543), .A2(n543), .ZN(n540) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n540), .Z(n646) );
  NAND2_X1 U599 ( .A1(G62), .A2(n646), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n548) );
  NOR2_X1 U601 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U602 ( .A1(G88), .A2(n648), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n638), .A2(n543), .ZN(n649) );
  NAND2_X1 U604 ( .A1(G75), .A2(n649), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT85), .B(n546), .Z(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U608 ( .A(KEYINPUT86), .B(n549), .ZN(G166) );
  INV_X1 U609 ( .A(G166), .ZN(G303) );
  NAND2_X1 U610 ( .A1(G52), .A2(n652), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G64), .A2(n646), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G90), .A2(n648), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G77), .A2(n649), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U617 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U621 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n648), .A2(G89), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G76), .A2(n649), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT5), .B(n560), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n652), .A2(G51), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT75), .B(n561), .Z(n563) );
  NAND2_X1 U629 ( .A1(n646), .A2(G63), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G168) );
  XOR2_X1 U634 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U637 ( .A(G223), .B(KEYINPUT71), .ZN(n832) );
  NAND2_X1 U638 ( .A1(n832), .A2(G567), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n572) );
  NAND2_X1 U641 ( .A1(G56), .A2(n646), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n572), .B(n571), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n648), .A2(G81), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G68), .A2(n649), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n652), .A2(G43), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n990) );
  INV_X1 U651 ( .A(G860), .ZN(n604) );
  OR2_X1 U652 ( .A1(n990), .A2(n604), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G79), .A2(n649), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT74), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G92), .A2(n648), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G54), .A2(n652), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G66), .A2(n646), .ZN(n584) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n584), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U664 ( .A(KEYINPUT15), .B(n589), .ZN(n996) );
  INV_X1 U665 ( .A(n996), .ZN(n859) );
  INV_X1 U666 ( .A(G868), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n859), .A2(n600), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U669 ( .A1(n649), .A2(G78), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT68), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G65), .A2(n646), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G91), .A2(n648), .ZN(n596) );
  NAND2_X1 U674 ( .A1(G53), .A2(n652), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n997) );
  XNOR2_X1 U677 ( .A(n997), .B(KEYINPUT69), .ZN(G299) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n599) );
  XOR2_X1 U679 ( .A(KEYINPUT77), .B(n599), .Z(n602) );
  NOR2_X1 U680 ( .A1(G286), .A2(n600), .ZN(n601) );
  NOR2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U682 ( .A(KEYINPUT78), .B(n603), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n604), .A2(G559), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n605), .A2(n996), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n990), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n996), .A2(G868), .ZN(n607) );
  NOR2_X1 U688 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U689 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G123), .A2(n532), .ZN(n610) );
  XOR2_X1 U691 ( .A(KEYINPUT79), .B(n610), .Z(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G135), .A2(n894), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G99), .A2(n897), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G111), .A2(n890), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n922) );
  XNOR2_X1 U699 ( .A(n922), .B(G2096), .ZN(n619) );
  INV_X1 U700 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U702 ( .A1(G559), .A2(n996), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n990), .B(n620), .ZN(n665) );
  NOR2_X1 U704 ( .A1(n665), .A2(G860), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G93), .A2(n648), .ZN(n622) );
  NAND2_X1 U706 ( .A1(G80), .A2(n649), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n622), .A2(n621), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G67), .A2(n646), .ZN(n623) );
  XNOR2_X1 U709 ( .A(n623), .B(KEYINPUT80), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n652), .A2(G55), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n661) );
  XNOR2_X1 U713 ( .A(n628), .B(n661), .ZN(G145) );
  NAND2_X1 U714 ( .A1(G73), .A2(n649), .ZN(n629) );
  XNOR2_X1 U715 ( .A(n629), .B(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G86), .A2(n648), .ZN(n631) );
  NAND2_X1 U717 ( .A1(G48), .A2(n652), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U719 ( .A1(G61), .A2(n646), .ZN(n632) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(n632), .ZN(n633) );
  NOR2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U723 ( .A(KEYINPUT84), .B(n637), .ZN(G305) );
  NAND2_X1 U724 ( .A1(n638), .A2(G87), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n639), .B(KEYINPUT82), .ZN(n641) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U728 ( .A1(n646), .A2(n642), .ZN(n645) );
  NAND2_X1 U729 ( .A1(G49), .A2(n652), .ZN(n643) );
  XOR2_X1 U730 ( .A(KEYINPUT81), .B(n643), .Z(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(G288) );
  NAND2_X1 U732 ( .A1(n646), .A2(G60), .ZN(n647) );
  XNOR2_X1 U733 ( .A(n647), .B(KEYINPUT66), .ZN(n657) );
  NAND2_X1 U734 ( .A1(G85), .A2(n648), .ZN(n651) );
  NAND2_X1 U735 ( .A1(G72), .A2(n649), .ZN(n650) );
  NAND2_X1 U736 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U737 ( .A1(G47), .A2(n652), .ZN(n653) );
  XNOR2_X1 U738 ( .A(KEYINPUT67), .B(n653), .ZN(n654) );
  NOR2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(G290) );
  NOR2_X1 U741 ( .A1(G868), .A2(n661), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(KEYINPUT87), .ZN(n668) );
  XNOR2_X1 U743 ( .A(KEYINPUT19), .B(G288), .ZN(n659) );
  XNOR2_X1 U744 ( .A(n659), .B(G299), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n661), .B(n660), .ZN(n663) );
  XNOR2_X1 U746 ( .A(G290), .B(G303), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U748 ( .A(G305), .B(n664), .Z(n858) );
  XOR2_X1 U749 ( .A(n858), .B(n665), .Z(n666) );
  NAND2_X1 U750 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XOR2_X1 U757 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G120), .A2(G69), .ZN(n673) );
  XOR2_X1 U760 ( .A(KEYINPUT89), .B(n673), .Z(n674) );
  NOR2_X1 U761 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U762 ( .A1(G108), .A2(n675), .ZN(n836) );
  NAND2_X1 U763 ( .A1(n836), .A2(G567), .ZN(n681) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U766 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U767 ( .A1(G96), .A2(n678), .ZN(n837) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n837), .ZN(n679) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n679), .ZN(n680) );
  NAND2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n839) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U772 ( .A1(n839), .A2(n682), .ZN(n835) );
  NAND2_X1 U773 ( .A1(n835), .A2(G36), .ZN(n683) );
  XNOR2_X1 U774 ( .A(KEYINPUT90), .B(n683), .ZN(G176) );
  NAND2_X1 U775 ( .A1(G288), .A2(G1976), .ZN(n684) );
  XNOR2_X1 U776 ( .A(n684), .B(KEYINPUT103), .ZN(n1013) );
  XOR2_X1 U777 ( .A(KEYINPUT99), .B(KEYINPUT27), .Z(n687) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n789) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n788) );
  INV_X1 U780 ( .A(n788), .ZN(n685) );
  NAND2_X1 U781 ( .A1(G2072), .A2(n712), .ZN(n686) );
  XNOR2_X1 U782 ( .A(n687), .B(n686), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n688), .A2(G1956), .ZN(n689) );
  XOR2_X1 U784 ( .A(KEYINPUT100), .B(n689), .Z(n690) );
  NOR2_X1 U785 ( .A1(n694), .A2(n997), .ZN(n693) );
  INV_X1 U786 ( .A(KEYINPUT28), .ZN(n692) );
  XNOR2_X1 U787 ( .A(n693), .B(n692), .ZN(n709) );
  NAND2_X1 U788 ( .A1(n997), .A2(n694), .ZN(n707) );
  INV_X1 U789 ( .A(G1996), .ZN(n951) );
  NOR2_X1 U790 ( .A1(n731), .A2(n951), .ZN(n695) );
  XOR2_X1 U791 ( .A(n695), .B(KEYINPUT26), .Z(n697) );
  NAND2_X1 U792 ( .A1(n731), .A2(G1341), .ZN(n696) );
  NAND2_X1 U793 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U794 ( .A1(n990), .A2(n698), .ZN(n699) );
  OR2_X1 U795 ( .A1(n996), .A2(n699), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n996), .A2(n699), .ZN(n703) );
  NAND2_X1 U797 ( .A1(G2067), .A2(n712), .ZN(n701) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n731), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U805 ( .A1(n712), .A2(n944), .ZN(n714) );
  INV_X1 U806 ( .A(G1961), .ZN(n972) );
  NAND2_X1 U807 ( .A1(n972), .A2(n731), .ZN(n713) );
  NAND2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n724), .A2(G171), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n730) );
  NAND2_X1 U811 ( .A1(G8), .A2(n731), .ZN(n767) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n767), .ZN(n743) );
  INV_X1 U813 ( .A(KEYINPUT97), .ZN(n718) );
  XNOR2_X1 U814 ( .A(n718), .B(n717), .ZN(n744) );
  NOR2_X1 U815 ( .A1(n743), .A2(n744), .ZN(n720) );
  INV_X1 U816 ( .A(KEYINPUT101), .ZN(n719) );
  XNOR2_X1 U817 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U818 ( .A1(n721), .A2(G8), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n722), .B(KEYINPUT30), .ZN(n723) );
  NOR2_X1 U820 ( .A1(G168), .A2(n723), .ZN(n726) );
  NOR2_X1 U821 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U822 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n741), .A2(G286), .ZN(n738) );
  INV_X1 U824 ( .A(G8), .ZN(n736) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n767), .ZN(n733) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n731), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U828 ( .A1(G303), .A2(n734), .ZN(n735) );
  OR2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U831 ( .A(n740), .B(n739), .ZN(n748) );
  INV_X1 U832 ( .A(n741), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n760) );
  INV_X1 U837 ( .A(n760), .ZN(n752) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  NOR2_X1 U839 ( .A1(G303), .A2(G1971), .ZN(n1009) );
  XNOR2_X1 U840 ( .A(KEYINPUT102), .B(n1009), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n1003), .A2(n749), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n767), .A2(n750), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n1013), .A2(n753), .ZN(n754) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n755) );
  XNOR2_X1 U846 ( .A(KEYINPUT104), .B(n755), .ZN(n994) );
  NAND2_X1 U847 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n517), .A2(n757), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n761), .A2(n767), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XOR2_X1 U855 ( .A(n765), .B(KEYINPUT24), .Z(n766) );
  NAND2_X1 U856 ( .A1(n894), .A2(G131), .ZN(n769) );
  XOR2_X1 U857 ( .A(KEYINPUT93), .B(n769), .Z(n771) );
  NAND2_X1 U858 ( .A1(n897), .A2(G95), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(KEYINPUT94), .B(n772), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n532), .A2(G119), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT92), .B(n773), .Z(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n890), .A2(G107), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n905) );
  NAND2_X1 U866 ( .A1(G1991), .A2(n905), .ZN(n786) );
  NAND2_X1 U867 ( .A1(G141), .A2(n894), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G117), .A2(n890), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n897), .A2(G105), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n780), .Z(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n532), .A2(G129), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n871) );
  NAND2_X1 U875 ( .A1(G1996), .A2(n871), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT95), .B(n787), .Z(n936) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n817) );
  NAND2_X1 U879 ( .A1(n936), .A2(n817), .ZN(n790) );
  XOR2_X1 U880 ( .A(KEYINPUT96), .B(n790), .Z(n808) );
  INV_X1 U881 ( .A(n808), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G140), .A2(n894), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G104), .A2(n897), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n793), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G116), .A2(n890), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G128), .A2(n532), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n799), .ZN(n875) );
  XNOR2_X1 U892 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U893 ( .A1(n875), .A2(n814), .ZN(n916) );
  NAND2_X1 U894 ( .A1(n817), .A2(n916), .ZN(n812) );
  NAND2_X1 U895 ( .A1(n800), .A2(n812), .ZN(n801) );
  NOR2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n804) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n1008) );
  NAND2_X1 U898 ( .A1(n1008), .A2(n817), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n820) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n871), .ZN(n919) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n905), .ZN(n924) );
  NOR2_X1 U903 ( .A1(n805), .A2(n924), .ZN(n806) );
  XNOR2_X1 U904 ( .A(n806), .B(KEYINPUT106), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U906 ( .A(KEYINPUT107), .B(n809), .Z(n810) );
  NOR2_X1 U907 ( .A1(n919), .A2(n810), .ZN(n811) );
  XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n875), .A2(n814), .ZN(n915) );
  NAND2_X1 U911 ( .A1(n815), .A2(n915), .ZN(n816) );
  XNOR2_X1 U912 ( .A(KEYINPUT108), .B(n816), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U916 ( .A(KEYINPUT109), .B(G2451), .Z(n823) );
  XNOR2_X1 U917 ( .A(G2446), .B(G2427), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n823), .B(n822), .ZN(n830) );
  XOR2_X1 U919 ( .A(G2438), .B(G2435), .Z(n825) );
  XNOR2_X1 U920 ( .A(G2443), .B(G2430), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U922 ( .A(n826), .B(G2454), .Z(n828) );
  XNOR2_X1 U923 ( .A(G1341), .B(G1348), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(G14), .ZN(n909) );
  XOR2_X1 U927 ( .A(KEYINPUT110), .B(n909), .Z(G401) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U930 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n835), .A2(n834), .ZN(G188) );
  XNOR2_X1 U933 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G108), .ZN(G238) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n838), .B(KEYINPUT112), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  INV_X1 U941 ( .A(n839), .ZN(G319) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2090), .Z(n843) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U947 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U948 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1961), .B(G1966), .Z(n849) );
  XNOR2_X1 U952 ( .A(G1976), .B(G1971), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U954 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U955 ( .A(G1981), .B(G1956), .ZN(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U957 ( .A(KEYINPUT41), .B(G1986), .Z(n854) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U959 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(G229) );
  XNOR2_X1 U961 ( .A(G171), .B(n990), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n857), .B(G286), .ZN(n861) );
  XOR2_X1 U963 ( .A(n859), .B(n858), .Z(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n862) );
  NOR2_X1 U965 ( .A1(G37), .A2(n862), .ZN(G397) );
  NAND2_X1 U966 ( .A1(G124), .A2(n532), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n863), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G112), .A2(n890), .ZN(n864) );
  XOR2_X1 U969 ( .A(KEYINPUT113), .B(n864), .Z(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G136), .A2(n894), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G100), .A2(n897), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U974 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT119), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n871), .B(KEYINPUT46), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U978 ( .A(G160), .B(G162), .Z(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(n904) );
  NAND2_X1 U981 ( .A1(n532), .A2(G130), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n878), .B(KEYINPUT114), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G118), .A2(n890), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n897), .A2(G106), .ZN(n881) );
  XNOR2_X1 U986 ( .A(KEYINPUT115), .B(n881), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n894), .A2(G142), .ZN(n882) );
  XOR2_X1 U988 ( .A(n882), .B(KEYINPUT116), .Z(n883) );
  NOR2_X1 U989 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n885), .Z(n886) );
  XNOR2_X1 U991 ( .A(n886), .B(KEYINPUT117), .ZN(n887) );
  NOR2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U993 ( .A(n889), .B(n922), .Z(n902) );
  NAND2_X1 U994 ( .A1(G115), .A2(n890), .ZN(n892) );
  NAND2_X1 U995 ( .A1(G127), .A2(n532), .ZN(n891) );
  NAND2_X1 U996 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U997 ( .A(n893), .B(KEYINPUT47), .ZN(n896) );
  NAND2_X1 U998 ( .A1(G139), .A2(n894), .ZN(n895) );
  NAND2_X1 U999 ( .A1(n896), .A2(n895), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n897), .A2(G103), .ZN(n898) );
  XOR2_X1 U1001 ( .A(KEYINPUT118), .B(n898), .Z(n899) );
  NOR2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(n927) );
  XNOR2_X1 U1003 ( .A(G164), .B(n927), .ZN(n901) );
  XNOR2_X1 U1004 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(KEYINPUT120), .B(n908), .ZN(G395) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n909), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G397), .A2(G395), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n915), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n934) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT51), .B(n920), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n926) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1025 ( .A(G2072), .B(n927), .Z(n929) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n930), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n937), .ZN(n939) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1036 ( .A(G2090), .B(G35), .Z(n943) );
  XOR2_X1 U1037 ( .A(G34), .B(KEYINPUT54), .Z(n941) );
  XNOR2_X1 U1038 ( .A(G2084), .B(n941), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n959) );
  XNOR2_X1 U1040 ( .A(G27), .B(n944), .ZN(n956) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1042 ( .A1(G28), .A2(n945), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT121), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1048 ( .A(G32), .B(n951), .Z(n952) );
  XNOR2_X1 U1049 ( .A(KEYINPUT122), .B(n952), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1052 ( .A(n957), .B(KEYINPUT53), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(KEYINPUT123), .B(n960), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT55), .B(n961), .ZN(n963) );
  INV_X1 U1056 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(G11), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT124), .B(n965), .ZN(n1020) );
  XNOR2_X1 U1060 ( .A(G1976), .B(G23), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G1971), .B(G22), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1063 ( .A(KEYINPUT126), .B(n968), .Z(n970) );
  XNOR2_X1 U1064 ( .A(G1986), .B(G24), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT58), .B(n971), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n972), .B(G5), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n987) );
  XOR2_X1 U1069 ( .A(G1966), .B(G21), .Z(n985) );
  XOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .Z(n975) );
  XNOR2_X1 U1071 ( .A(G4), .B(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(G19), .B(G1341), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(G20), .B(G1956), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n982), .B(KEYINPUT60), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n983), .B(KEYINPUT125), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1082 ( .A(KEYINPUT61), .B(n988), .Z(n989) );
  NOR2_X1 U1083 ( .A1(G16), .A2(n989), .ZN(n1017) );
  XOR2_X1 U1084 ( .A(G16), .B(KEYINPUT56), .Z(n1015) );
  NAND2_X1 U1085 ( .A1(G303), .A2(G1971), .ZN(n992) );
  XOR2_X1 U1086 ( .A(G1341), .B(n990), .Z(n991) );
  NAND2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n1007) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G168), .ZN(n993) );
  NAND2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(n995), .B(KEYINPUT57), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n996), .B(G1348), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(n997), .B(G1956), .Z(n999) );
  XOR2_X1 U1093 ( .A(G171), .B(G1961), .Z(n998) );
  NOR2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT127), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

