//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G107), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT65), .B(G244), .Z(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G77), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n206), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n205), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n206), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n229), .B(new_n234), .C1(new_n221), .C2(new_n222), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n224), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT69), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT70), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n227), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G50), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n205), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n262), .A2(new_n263), .B1(new_n205), .B2(G68), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n257), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT11), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT78), .B1(new_n268), .B2(G68), .ZN(new_n269));
  XOR2_X1   g0069(.A(new_n269), .B(KEYINPUT12), .Z(new_n270));
  INV_X1    g0070(.A(new_n268), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n257), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n204), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G68), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n265), .A2(new_n266), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n267), .A2(new_n270), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n214), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G226), .B2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G97), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n279), .A2(new_n284), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n227), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(KEYINPUT71), .A2(G33), .A3(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n287), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(G274), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n216), .B1(new_n302), .B2(KEYINPUT76), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(KEYINPUT76), .B2(new_n302), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT13), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT77), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n300), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(KEYINPUT77), .A3(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(G169), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n308), .B1(new_n300), .B2(new_n304), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n312), .A2(KEYINPUT14), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n310), .A2(new_n317), .A3(G169), .A4(new_n311), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n277), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(G200), .A3(new_n311), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n276), .B1(new_n322), .B2(new_n309), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n295), .A2(new_n301), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G226), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G222), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G223), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n290), .C1(G77), .C2(new_n328), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n327), .A2(new_n333), .A3(new_n299), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT74), .A3(G190), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT74), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n327), .A2(new_n333), .A3(new_n299), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n321), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n260), .B1(new_n204), .B2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n272), .A2(new_n339), .B1(new_n260), .B2(new_n271), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n341), .A2(new_n262), .B1(new_n342), .B2(new_n259), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G50), .A2(G58), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n205), .B1(new_n344), .B2(new_n215), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n257), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT9), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT9), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n340), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n335), .A2(new_n338), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n337), .A2(G200), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n335), .A2(new_n338), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n349), .A2(new_n351), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(KEYINPUT73), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n352), .B(new_n353), .C1(KEYINPUT73), .C2(KEYINPUT10), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n334), .A2(new_n314), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n337), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n348), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n347), .A2(new_n268), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n273), .A2(G77), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(G77), .B2(new_n268), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT8), .B(G58), .Z(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n262), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n372), .B2(new_n257), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n328), .A2(G238), .A3(G1698), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n328), .A2(G232), .A3(new_n330), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n328), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n290), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n326), .A2(new_n219), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n299), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n373), .B1(new_n380), .B2(new_n363), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G179), .B2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(G200), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n373), .C1(new_n321), .C2(new_n380), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT72), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT72), .B1(new_n382), .B2(new_n384), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n361), .A2(KEYINPUT75), .A3(new_n365), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT79), .B1(new_n280), .B2(KEYINPUT3), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT79), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n282), .A3(G33), .ZN(new_n392));
  AND2_X1   g0192(.A1(G226), .A2(G1698), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n390), .A2(new_n392), .A3(new_n281), .A4(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n392), .A3(new_n281), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT81), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n393), .A2(new_n398), .B1(G223), .B2(new_n330), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n290), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n295), .A2(new_n301), .A3(G232), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n299), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n363), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G226), .A2(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(G223), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n407), .A2(KEYINPUT81), .B1(new_n408), .B2(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(new_n281), .A3(new_n390), .A4(new_n392), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n396), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n411), .B2(new_n290), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n405), .B1(G179), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n341), .B1(new_n204), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n272), .B1(new_n271), .B2(new_n341), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n390), .A2(new_n392), .A3(new_n281), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT7), .B1(new_n417), .B2(G20), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n397), .A2(new_n419), .A3(new_n205), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(G68), .A3(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G58), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n258), .A2(G159), .ZN(new_n427));
  OAI211_X1 g0227(.A(KEYINPUT80), .B(G20), .C1(new_n422), .C2(new_n423), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT16), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n347), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n419), .B1(new_n328), .B2(G20), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n205), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n215), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n430), .B1(new_n435), .B2(new_n429), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n416), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT18), .B1(new_n413), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n428), .A2(new_n427), .ZN(new_n439));
  XNOR2_X1  g0239(.A(G58), .B(G68), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT80), .B1(new_n440), .B2(G20), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n420), .A2(G68), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n419), .B1(new_n397), .B2(new_n205), .ZN(new_n444));
  OAI211_X1 g0244(.A(KEYINPUT16), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n257), .A3(new_n436), .ZN(new_n446));
  AOI211_X1 g0246(.A(G190), .B(new_n403), .C1(new_n290), .C2(new_n411), .ZN(new_n447));
  AOI21_X1  g0247(.A(G200), .B1(new_n401), .B2(new_n404), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n415), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n415), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n401), .A2(G179), .A3(new_n404), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n363), .B2(new_n412), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n401), .A2(new_n321), .A3(new_n404), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G200), .B2(new_n412), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n438), .A2(new_n451), .A3(new_n456), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n359), .A2(new_n360), .A3(new_n365), .ZN(new_n463));
  INV_X1    g0263(.A(new_n387), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n385), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g0266(.A1(new_n325), .A2(new_n389), .A3(new_n461), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G244), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1698), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT4), .B1(new_n417), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n328), .A2(G250), .A3(G1698), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT4), .A2(G244), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n328), .A2(new_n330), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n290), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n297), .A2(G1), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n295), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G257), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT83), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n295), .A2(new_n482), .A3(new_n486), .A4(G257), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n481), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n479), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n295), .A2(new_n490), .A3(G274), .A4(new_n478), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n477), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n285), .B2(G107), .ZN(new_n495));
  XNOR2_X1  g0295(.A(G97), .B(G107), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(G20), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n258), .A2(G77), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n376), .B1(new_n433), .B2(new_n434), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n257), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n268), .A2(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n204), .A2(G33), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n347), .A2(new_n268), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(G97), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n477), .A2(new_n488), .A3(G190), .A4(new_n491), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n493), .A2(new_n501), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n492), .A2(new_n363), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n501), .A2(new_n506), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n477), .A2(new_n488), .A3(new_n314), .A4(new_n491), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n284), .A2(G303), .ZN(new_n514));
  INV_X1    g0314(.A(G264), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G1698), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G257), .B2(G1698), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n397), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n290), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n491), .C1(new_n210), .C2(new_n483), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n517), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n417), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n289), .B1(new_n523), .B2(new_n514), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n491), .B1(new_n483), .B2(new_n210), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G190), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n271), .A2(new_n209), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n256), .A2(new_n227), .B1(G20), .B2(new_n209), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n475), .B(new_n205), .C1(G33), .C2(new_n285), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT20), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  OAI221_X1 g0332(.A(new_n528), .B1(new_n504), .B2(new_n209), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n521), .A2(new_n527), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT21), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n531), .A2(new_n532), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n528), .B1(new_n504), .B2(new_n209), .ZN(new_n538));
  OAI21_X1  g0338(.A(G169), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n520), .A2(new_n533), .A3(KEYINPUT21), .A4(G169), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n526), .A2(G179), .A3(new_n533), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n535), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n205), .B1(new_n280), .B2(new_n285), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n207), .A2(new_n285), .A3(new_n376), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n262), .A2(KEYINPUT19), .A3(new_n285), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n390), .A2(new_n392), .A3(new_n205), .A4(new_n281), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n215), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n257), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n371), .A2(new_n271), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n505), .A2(G87), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n469), .A2(G1698), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G238), .B2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n397), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n290), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n208), .B1(new_n297), .B2(G1), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n297), .A2(G1), .A3(G274), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n295), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n563), .A3(G190), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT85), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n290), .B2(new_n558), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT85), .A3(G190), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n559), .A2(new_n563), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G200), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n554), .A2(new_n566), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n363), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n371), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n505), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n551), .A2(new_n552), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(new_n314), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n513), .A2(new_n543), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT22), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n205), .A2(G87), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n284), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n376), .A3(G20), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT86), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(KEYINPUT23), .B2(G107), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n205), .A2(KEYINPUT23), .A3(G107), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n555), .A2(new_n584), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(KEYINPUT86), .B1(new_n589), .B2(new_n205), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n583), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n581), .A2(new_n207), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n549), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT24), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n417), .A2(new_n205), .A3(new_n592), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n588), .A2(KEYINPUT86), .B1(new_n584), .B2(new_n376), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n585), .A2(new_n586), .B1(new_n598), .B2(G20), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n596), .A2(new_n600), .A3(new_n601), .A4(new_n583), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n257), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT25), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n268), .A2(new_n605), .A3(G107), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n268), .B2(G107), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n505), .A2(G107), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n484), .A2(G1698), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(G250), .B2(G1698), .ZN(new_n612));
  INV_X1    g0412(.A(G294), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n397), .A2(new_n612), .B1(new_n280), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n290), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n295), .A2(new_n482), .A3(G264), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n491), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n363), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n615), .A2(new_n314), .A3(new_n491), .A4(new_n616), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n620), .A3(KEYINPUT87), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  INV_X1    g0422(.A(new_n609), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n603), .B2(new_n257), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n618), .A2(new_n619), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n483), .ZN(new_n627));
  AOI22_X1  g0427(.A1(G264), .A2(new_n627), .B1(new_n614), .B2(new_n290), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(G190), .A3(new_n491), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n617), .A2(G200), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n621), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n580), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n468), .A2(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n365), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n324), .A2(new_n382), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n451), .B(new_n459), .C1(new_n319), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n438), .A3(new_n456), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(new_n361), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n550), .A2(new_n257), .B1(new_n271), .B2(new_n371), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n570), .A2(new_n640), .A3(new_n553), .A4(new_n564), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n578), .ZN(new_n642));
  OR3_X1    g0442(.A1(new_n512), .A2(new_n642), .A3(KEYINPUT26), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n492), .A2(new_n363), .B1(new_n501), .B2(new_n506), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n571), .A3(new_n511), .A4(new_n578), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n578), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n513), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n641), .A2(new_n578), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n631), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n610), .A2(new_n620), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n624), .A2(new_n625), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT88), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n649), .A2(new_n651), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n639), .B1(new_n468), .B2(new_n661), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G343), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n653), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n610), .A2(new_n669), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n621), .A2(new_n626), .A3(new_n671), .A4(new_n631), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n656), .A2(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n657), .A2(new_n668), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n670), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n534), .A2(new_n668), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n657), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n543), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(KEYINPUT89), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n684), .B2(G330), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n672), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT90), .B1(new_n672), .B2(new_n673), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n686), .A2(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n681), .A2(new_n691), .ZN(G399));
  OR3_X1    g0492(.A1(new_n231), .A2(KEYINPUT91), .A3(G41), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT91), .B1(new_n231), .B2(G41), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n546), .A2(G116), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n204), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n226), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND3_X1  g0500(.A1(new_n580), .A2(new_n632), .A3(new_n668), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n526), .A2(new_n567), .A3(G179), .A4(new_n628), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n492), .ZN(new_n705));
  INV_X1    g0505(.A(new_n492), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n520), .A2(new_n314), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n628), .A2(new_n567), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT30), .A4(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n526), .A2(new_n567), .A3(G179), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n617), .A3(new_n492), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT92), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n669), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n712), .A2(KEYINPUT92), .A3(KEYINPUT31), .A4(new_n669), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(G330), .B1(new_n702), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n578), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n644), .A2(new_n511), .A3(new_n578), .A4(new_n641), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT26), .ZN(new_n725));
  OR3_X1    g0525(.A1(new_n579), .A2(new_n512), .A3(KEYINPUT26), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n621), .A2(new_n652), .A3(new_n626), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n650), .A2(new_n508), .A3(new_n631), .A4(new_n512), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n725), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n729), .A2(KEYINPUT93), .A3(new_n668), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT93), .B1(new_n729), .B2(new_n668), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT29), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n660), .A2(new_n668), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n722), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n700), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n686), .A2(new_n688), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n205), .A2(G13), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n204), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n738), .B1(G330), .B2(new_n684), .C1(new_n696), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n696), .A2(new_n742), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n231), .A2(new_n284), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G355), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G116), .B2(new_n232), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n251), .A2(G45), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n417), .A2(new_n231), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n297), .B2(new_n226), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n227), .B1(G20), .B2(new_n363), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n744), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n205), .A2(G179), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G159), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n205), .A2(new_n314), .ZN(new_n767));
  INV_X1    g0567(.A(G200), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n767), .A2(G190), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n321), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n328), .B1(new_n213), .B2(new_n769), .C1(new_n772), .C2(new_n260), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n767), .A2(new_n762), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT96), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(KEYINPUT96), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n766), .B(new_n773), .C1(G77), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT97), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n761), .A2(new_n321), .A3(G200), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT98), .Z(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G107), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n321), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n205), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n770), .A2(G190), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G97), .A2(new_n792), .B1(new_n793), .B2(G68), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n779), .A2(new_n786), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n793), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n798), .B1(new_n769), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT100), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n771), .A2(G326), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n328), .B1(new_n764), .B2(G329), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n613), .C2(new_n791), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G311), .B2(new_n778), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n785), .A2(G303), .B1(new_n788), .B2(G283), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n801), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n796), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n760), .B1(new_n808), .B2(new_n757), .ZN(new_n809));
  INV_X1    g0609(.A(new_n756), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n684), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n743), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  INV_X1    g0613(.A(KEYINPUT105), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n382), .B(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n815), .A2(new_n384), .ZN(new_n816));
  AND4_X1   g0616(.A1(new_n649), .A2(new_n651), .A3(new_n655), .A4(new_n658), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n668), .C1(new_n817), .C2(new_n647), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n669), .B1(new_n648), .B2(new_n659), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n815), .B(new_n384), .C1(new_n373), .C2(new_n668), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n382), .A2(new_n668), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n744), .B1(new_n823), .B2(new_n721), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n721), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n757), .A2(new_n754), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n744), .B1(G77), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT102), .Z(new_n829));
  INV_X1    g0629(.A(new_n788), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(new_n207), .B1(new_n376), .B2(new_n784), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n284), .B1(new_n763), .B2(new_n832), .C1(new_n769), .C2(new_n613), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n778), .B2(G116), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G97), .A2(new_n792), .B1(new_n771), .B2(G303), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n797), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT103), .ZN(new_n839));
  INV_X1    g0639(.A(new_n769), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n797), .B2(new_n342), .C1(new_n842), .C2(new_n772), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G159), .B2(new_n778), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT34), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n788), .A2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n417), .B1(new_n848), .B2(new_n763), .C1(new_n213), .C2(new_n791), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n785), .B2(G50), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n829), .B1(new_n852), .B2(new_n757), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT104), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n755), .B2(new_n822), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n825), .A2(new_n855), .ZN(G384));
  OAI21_X1  g0656(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT35), .ZN(new_n858));
  OAI211_X1 g0658(.A(G116), .B(new_n228), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  XOR2_X1   g0660(.A(KEYINPUT106), .B(KEYINPUT36), .Z(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n226), .B(G77), .C1(new_n213), .C2(new_n215), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n260), .A2(G68), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n204), .B(G13), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n277), .A2(new_n668), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n319), .B2(new_n324), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n315), .A2(new_n309), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n318), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n276), .ZN(new_n872));
  INV_X1    g0672(.A(new_n324), .ZN(new_n873));
  INV_X1    g0673(.A(new_n867), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n718), .A2(new_n713), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n701), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n822), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n443), .A2(new_n444), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n430), .B1(new_n880), .B2(new_n429), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n416), .B1(new_n881), .B2(new_n432), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n449), .B1(new_n666), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n413), .A2(new_n882), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n452), .A2(new_n455), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n452), .A2(new_n667), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n449), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n882), .A2(new_n666), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n460), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT107), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n896), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  INV_X1    g0701(.A(new_n879), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT109), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n886), .A2(new_n887), .A3(new_n449), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  INV_X1    g0705(.A(new_n887), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n889), .A2(new_n905), .B1(new_n460), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n889), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n460), .A2(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(KEYINPUT109), .A3(new_n894), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n896), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n467), .A2(new_n878), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n901), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n917), .B1(new_n901), .B2(new_n916), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(G330), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n871), .A2(new_n276), .A3(new_n668), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT108), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n319), .A2(new_n923), .A3(new_n668), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n889), .A2(new_n885), .B1(new_n460), .B2(new_n891), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT39), .B1(new_n926), .B2(KEYINPUT38), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT109), .B1(new_n911), .B2(new_n894), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n903), .B(KEYINPUT38), .C1(new_n909), .C2(new_n910), .ZN(new_n929));
  OAI211_X1 g0729(.A(KEYINPUT110), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n895), .B2(new_n896), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT110), .B1(new_n913), .B2(new_n927), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n925), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n898), .A2(new_n899), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n815), .A2(new_n669), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n818), .A2(new_n939), .B1(new_n868), .B2(new_n875), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n438), .A2(new_n456), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n937), .A2(new_n940), .B1(new_n941), .B2(new_n666), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n732), .A2(new_n467), .A3(new_n735), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n639), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n943), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n920), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n204), .B2(new_n740), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n920), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n866), .B1(new_n948), .B2(new_n949), .ZN(G367));
  NAND2_X1  g0750(.A1(new_n510), .A2(new_n669), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n649), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n644), .A2(new_n511), .A3(new_n669), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n691), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n554), .A2(new_n668), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n578), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n650), .B2(new_n957), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT111), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n679), .B1(new_n676), .B2(new_n677), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n954), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n621), .A2(new_n626), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n649), .A2(new_n966), .A3(new_n951), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n669), .B1(new_n967), .B2(new_n512), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n964), .B2(KEYINPUT42), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n962), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n960), .A2(new_n961), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n965), .A2(new_n969), .A3(new_n961), .A4(new_n960), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n956), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n956), .A3(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT112), .B(KEYINPUT41), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n695), .B(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n685), .B(KEYINPUT89), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n680), .B1(new_n689), .B2(new_n690), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n982), .B1(new_n984), .B2(new_n983), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n736), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT114), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n691), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n670), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n983), .A2(new_n991), .A3(new_n954), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n983), .A2(KEYINPUT45), .A3(new_n991), .A4(new_n954), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n681), .B2(new_n954), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n955), .B(new_n999), .C1(new_n963), .C2(new_n670), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n691), .A2(new_n989), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n996), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n988), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n732), .A2(new_n735), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n721), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n981), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n978), .B1(new_n1010), .B2(new_n741), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n246), .A2(new_n750), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n758), .B1(new_n232), .B2(new_n371), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n744), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n284), .B1(new_n764), .B2(G137), .ZN(new_n1015));
  INV_X1    g0815(.A(G159), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n263), .B2(new_n787), .C1(new_n797), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G50), .B2(new_n778), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n213), .B2(new_n784), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G143), .A2(new_n771), .B1(new_n840), .B2(G150), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n215), .B2(new_n791), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT115), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n784), .A2(new_n209), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT46), .ZN(new_n1024));
  INV_X1    g0824(.A(G317), .ZN(new_n1025));
  INV_X1    g0825(.A(G303), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n397), .B1(new_n763), .B2(new_n1025), .C1(new_n769), .C2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n778), .B2(G283), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G107), .A2(new_n792), .B1(new_n793), .B2(G294), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n787), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n771), .A2(G311), .B1(new_n1030), .B2(G97), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1019), .A2(new_n1022), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1014), .B1(new_n1034), .B2(new_n757), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n960), .A2(new_n756), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1011), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n987), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n678), .A2(new_n810), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1016), .A2(new_n772), .B1(new_n797), .B2(new_n341), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT116), .B(G150), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n769), .A2(new_n260), .B1(new_n763), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n397), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n574), .A2(new_n792), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n785), .A2(G77), .B1(new_n788), .B2(G97), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n778), .A2(G68), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n417), .B1(G326), .B2(new_n764), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n784), .A2(new_n613), .B1(new_n836), .B2(new_n791), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G311), .A2(new_n793), .B1(new_n840), .B2(G317), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n778), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1052), .B1(new_n799), .B2(new_n772), .C1(new_n1053), .C2(new_n1026), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1050), .B1(new_n209), .B2(new_n787), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n757), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n369), .B2(new_n260), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n341), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n297), .B1(new_n215), .B2(new_n263), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n697), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n242), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n750), .B1(new_n1068), .B2(new_n297), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n746), .A2(new_n697), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n232), .A2(G107), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n758), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1062), .A2(new_n744), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1040), .A2(new_n741), .B1(new_n1041), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1040), .A2(new_n1009), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n696), .A3(new_n988), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(new_n988), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n996), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1003), .B1(new_n996), .B2(new_n1001), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1005), .A2(new_n988), .A3(new_n1006), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n696), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n742), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n758), .B1(new_n285), .B2(new_n232), .C1(new_n751), .C2(new_n254), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n744), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT51), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n772), .A2(new_n342), .B1(new_n1016), .B2(new_n769), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1089), .A2(new_n1090), .B1(new_n785), .B2(G68), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n1089), .B2(new_n1090), .C1(new_n207), .C2(new_n830), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n397), .B1(new_n764), .B2(G143), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G77), .A2(new_n792), .B1(new_n793), .B2(G50), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n1053), .C2(new_n341), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n772), .A2(new_n1025), .B1(new_n832), .B2(new_n769), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT52), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1096), .A2(new_n1097), .B1(new_n788), .B2(G107), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n1097), .B2(new_n1096), .C1(new_n836), .C2(new_n784), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n284), .B1(new_n763), .B2(new_n799), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G303), .B2(new_n793), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n209), .B2(new_n791), .C1(new_n1053), .C2(new_n613), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1092), .A2(new_n1095), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1088), .B1(new_n1103), .B2(new_n757), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n954), .B2(new_n810), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1085), .A2(new_n1086), .A3(new_n1105), .ZN(G390));
  INV_X1    g0906(.A(G330), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n877), .B2(new_n701), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n876), .A2(new_n1108), .A3(new_n822), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n818), .A2(new_n939), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n925), .B1(new_n1111), .B2(new_n876), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n934), .A2(new_n935), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n874), .B1(new_n872), .B2(new_n873), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n867), .B(new_n324), .C1(new_n871), .C2(new_n276), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n822), .B1(new_n730), .B2(new_n731), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n939), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n925), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n914), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1110), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n731), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n729), .A2(KEYINPUT93), .A3(new_n668), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n938), .B1(new_n1125), .B2(new_n822), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1119), .B(new_n914), .C1(new_n1126), .C2(new_n1116), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n896), .A2(new_n931), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n908), .B2(new_n912), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n932), .B1(new_n1129), .B2(KEYINPUT110), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n913), .A2(new_n927), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT110), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n938), .B1(new_n819), .B2(new_n816), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1119), .B1(new_n1134), .B2(new_n1116), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1130), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n722), .A2(new_n822), .A3(new_n876), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1127), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1122), .A2(new_n1138), .A3(new_n742), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n934), .A2(new_n755), .A3(new_n935), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G107), .A2(new_n793), .B1(new_n771), .B2(G283), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1053), .B2(new_n285), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT118), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n791), .A2(new_n263), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n284), .B1(new_n763), .B2(new_n613), .C1(new_n769), .C2(new_n209), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n785), .C2(G87), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n847), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT119), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n784), .A2(new_n1043), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G159), .A2(new_n792), .B1(new_n793), .B2(G137), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n771), .A2(G128), .B1(new_n1030), .B2(G50), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n284), .B1(new_n764), .B2(G125), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n848), .B2(new_n769), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT54), .B(G143), .Z(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT117), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n778), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1159), .A2(KEYINPUT120), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n757), .B1(new_n1159), .B2(KEYINPUT120), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n744), .B1(new_n369), .B2(new_n827), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1140), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1139), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1122), .A2(new_n1138), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n467), .A2(new_n1108), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n944), .A2(new_n639), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n822), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1116), .B1(new_n721), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1109), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1111), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1108), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1116), .B1(new_n1172), .B2(new_n1168), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1126), .A2(new_n1173), .A3(new_n1137), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1167), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n695), .B1(new_n1165), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1122), .A2(new_n1138), .A3(new_n1175), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1164), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G378));
  NAND2_X1  g0980(.A1(new_n348), .A2(new_n667), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n463), .B(new_n1181), .Z(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT121), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1119), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n899), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n940), .B1(new_n1188), .B2(new_n897), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n941), .A2(new_n666), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n936), .A2(new_n942), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n915), .B(G330), .C1(new_n900), .C2(KEYINPUT40), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1192), .A2(new_n1196), .A3(new_n1194), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n742), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n744), .B1(G50), .B2(new_n827), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n787), .A2(new_n213), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G116), .B2(new_n771), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n285), .B2(new_n797), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G77), .B2(new_n785), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n778), .A2(new_n574), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n296), .B1(new_n763), .B2(new_n836), .C1(new_n769), .C2(new_n376), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n417), .B(new_n1207), .C1(G68), .C2(new_n792), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n296), .B1(new_n397), .B2(new_n280), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1209), .A2(new_n1210), .B1(new_n260), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n785), .A2(new_n1156), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n778), .A2(G137), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G125), .A2(new_n771), .B1(new_n840), .B2(G128), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G150), .A2(new_n792), .B1(new_n793), .B2(G132), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1030), .A2(G159), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1212), .B1(new_n1210), .B2(new_n1209), .C1(new_n1218), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1201), .B1(new_n1223), .B2(new_n757), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1184), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n755), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1200), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1167), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1178), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1229), .A2(KEYINPUT57), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n696), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1192), .A2(new_n1196), .A3(new_n1194), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1196), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1229), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1227), .B1(new_n1231), .B2(new_n1235), .ZN(G375));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1239), .B2(new_n741), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(KEYINPUT123), .A3(new_n742), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n744), .B1(G68), .B2(new_n827), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1046), .B1(new_n836), .B2(new_n769), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT124), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n284), .B1(new_n763), .B2(new_n1026), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G294), .B2(new_n771), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n209), .B2(new_n797), .C1(new_n1053), .C2(new_n376), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n830), .A2(new_n263), .B1(new_n784), .B2(new_n285), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT125), .ZN(new_n1250));
  INV_X1    g1050(.A(G128), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n417), .B1(new_n1251), .B2(new_n763), .C1(new_n842), .C2(new_n769), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n778), .B2(G150), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1156), .A2(new_n793), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n791), .A2(new_n260), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1202), .B(new_n1255), .C1(G132), .C2(new_n771), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n785), .A2(G159), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1259), .A2(KEYINPUT126), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n757), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1259), .B2(KEYINPUT126), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1242), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n755), .B2(new_n876), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1240), .A2(new_n1241), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1238), .A2(new_n1228), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n980), .B(KEYINPUT122), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1176), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(G381));
  NOR4_X1   g1071(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1272));
  INV_X1    g1072(.A(G390), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1038), .A3(new_n1273), .A4(new_n1179), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(G375), .ZN(G407));
  INV_X1    g1075(.A(G343), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1179), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(G375), .C2(new_n1277), .ZN(G409));
  NOR2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n812), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n977), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(new_n975), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n980), .B1(new_n1083), .B2(new_n736), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(new_n742), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1037), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1286), .A2(new_n1287), .A3(G390), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1282), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1273), .B1(new_n1011), .B2(new_n1037), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1287), .A3(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1281), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G378), .B(new_n1227), .C1(new_n1231), .C2(new_n1235), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1234), .A2(new_n1229), .A3(new_n1269), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1200), .A2(new_n1226), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1179), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1276), .A2(G213), .ZN(new_n1301));
  INV_X1    g1101(.A(G384), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1171), .A2(new_n1174), .A3(new_n1167), .A4(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n696), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1268), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1306), .B2(new_n1265), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1306), .A2(new_n1265), .A3(new_n1302), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .A4(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1295), .A2(new_n1298), .B1(G213), .B2(new_n1276), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1276), .A2(G213), .A3(G2897), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1316));
  OR3_X1    g1116(.A1(new_n1306), .A2(new_n1265), .A3(new_n1302), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1307), .A3(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1311), .B(new_n1312), .C1(new_n1313), .C2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1300), .B1(new_n1313), .B2(new_n1310), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1294), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT63), .B1(new_n1313), .B2(new_n1319), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1313), .A2(new_n1310), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1290), .A2(new_n1312), .A3(new_n1293), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1326), .B(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1310), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1322), .A2(new_n1330), .ZN(G405));
  INV_X1    g1131(.A(new_n1310), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1179), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1295), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1332), .B1(new_n1333), .B2(new_n1295), .ZN(new_n1336));
  OR3_X1    g1136(.A1(new_n1335), .A2(new_n1336), .A3(new_n1294), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1294), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


