//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n190), .A2(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT65), .B1(new_n188), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n190), .A3(G146), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n193), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n207), .A3(new_n211), .A4(new_n208), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n202), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n204), .A2(G137), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n206), .A2(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(G131), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n195), .A2(new_n197), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n189), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n189), .A2(new_n191), .A3(new_n224), .A4(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n217), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n227), .B2(G119), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G116), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(G119), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n235));
  INV_X1    g049(.A(G113), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(KEYINPUT2), .B2(G113), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n237), .A2(new_n239), .B1(KEYINPUT2), .B2(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n239), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT2), .A2(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT68), .A3(new_n233), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n213), .A2(new_n226), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n193), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n219), .B2(new_n200), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n210), .A2(new_n212), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n212), .A2(new_n216), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n225), .B1(new_n198), .B2(new_n221), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n251), .A2(new_n254), .B1(new_n241), .B2(new_n245), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT28), .B1(new_n247), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n258), .B(KEYINPUT71), .Z(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n259), .B(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n249), .A2(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n264));
  INV_X1    g078(.A(new_n246), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT28), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n256), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n271));
  OAI21_X1  g085(.A(KEYINPUT66), .B1(new_n264), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n273));
  INV_X1    g087(.A(new_n271), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n273), .B(new_n274), .C1(new_n213), .C2(new_n226), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n264), .A2(KEYINPUT30), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n272), .A2(new_n275), .A3(new_n246), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n264), .A2(new_n265), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n263), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n270), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n246), .B1(new_n213), .B2(new_n226), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n278), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n266), .B1(new_n282), .B2(KEYINPUT28), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT29), .B1(new_n283), .B2(new_n263), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n278), .ZN(new_n285));
  INV_X1    g099(.A(new_n263), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n287), .A3(KEYINPUT72), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT73), .B(G902), .Z(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n268), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n280), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G472), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n277), .A2(new_n263), .A3(new_n278), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n277), .A2(new_n299), .A3(new_n263), .A4(new_n278), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n256), .A2(new_n267), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n286), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(G472), .A2(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n307), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n293), .A2(KEYINPUT74), .A3(G472), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n296), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n289), .B2(G234), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n220), .A2(KEYINPUT23), .A3(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n230), .A2(G128), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n230), .A2(G128), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(KEYINPUT23), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT24), .B(G110), .Z(new_n319));
  XNOR2_X1  g133(.A(G119), .B(G128), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n318), .A2(G110), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT75), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT16), .B1(new_n323), .B2(G125), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n188), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n188), .B1(new_n326), .B2(new_n328), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n321), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  OAI22_X1  g147(.A1(new_n318), .A2(G110), .B1(new_n319), .B2(new_n320), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n323), .A2(G125), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n337), .A3(new_n188), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT76), .ZN(new_n339));
  XNOR2_X1  g153(.A(G125), .B(G140), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n188), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n334), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G221), .A3(G234), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n347), .A2(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(KEYINPUT77), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n348), .B2(new_n349), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n345), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n332), .A2(new_n344), .A3(new_n353), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n289), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n289), .A4(new_n356), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n314), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n356), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n353), .B1(new_n332), .B2(new_n344), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n313), .A2(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n355), .A2(new_n356), .A3(new_n366), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n361), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n311), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G952), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G953), .ZN(new_n374));
  NAND2_X1  g188(.A1(G234), .A2(G237), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n290), .A2(G953), .A3(new_n375), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT21), .B(G898), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G128), .B(G143), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n190), .A2(G128), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n382), .B(G134), .C1(KEYINPUT13), .C2(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(G116), .B(G122), .Z(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G107), .ZN(new_n386));
  XNOR2_X1  g200(.A(G116), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n381), .A2(new_n204), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n381), .B(new_n204), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n227), .A2(KEYINPUT14), .A3(G122), .ZN(new_n394));
  OAI211_X1 g208(.A(G107), .B(new_n394), .C1(new_n385), .C2(KEYINPUT14), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT9), .B(G234), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n398), .A2(new_n312), .A3(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n396), .A3(new_n399), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n289), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT93), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT15), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(new_n408), .A3(new_n289), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n404), .A2(new_n407), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n415));
  AOI21_X1  g229(.A(G143), .B1(new_n257), .B2(G214), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT18), .B(G131), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n324), .A2(G146), .A3(new_n325), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n341), .B1(new_n340), .B2(new_n188), .ZN(new_n419));
  AND4_X1   g233(.A1(new_n341), .A2(new_n335), .A3(new_n337), .A4(new_n188), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT90), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n415), .A2(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT18), .A2(G131), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G237), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n346), .A3(G214), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n190), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n422), .A2(new_n428), .A3(new_n429), .A4(new_n424), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n417), .B(new_n421), .C1(new_n425), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G113), .B(G122), .ZN(new_n432));
  INV_X1    g246(.A(G104), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n415), .B2(new_n416), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n428), .A2(new_n211), .A3(new_n429), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(KEYINPUT17), .B(G131), .C1(new_n415), .C2(new_n416), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n438), .A2(new_n329), .A3(new_n333), .A4(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n431), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n324), .A2(KEYINPUT19), .A3(new_n325), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n335), .A2(new_n337), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n442), .B1(new_n446), .B2(G146), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n435), .A2(new_n437), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n443), .A2(new_n445), .A3(KEYINPUT91), .A4(new_n188), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n333), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n434), .B1(new_n431), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n414), .B1(new_n441), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT20), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(new_n414), .C1(new_n441), .C2(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G902), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n434), .B1(new_n431), .B2(new_n440), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n441), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G475), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n456), .A2(KEYINPUT92), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT92), .B1(new_n456), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n380), .B(new_n413), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n253), .A2(new_n336), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n336), .B2(new_n202), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n346), .A2(G224), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G122), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n388), .A2(KEYINPUT80), .A3(G104), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n388), .A3(KEYINPUT80), .A4(G104), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n433), .A2(G107), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G101), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT81), .B(G101), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n474), .A2(new_n480), .A3(new_n476), .A4(new_n477), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n472), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G101), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n473), .A2(KEYINPUT3), .B1(new_n433), .B2(G107), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n476), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n246), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n246), .C1(new_n482), .C2(new_n486), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n244), .A2(new_n233), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT87), .B(KEYINPUT5), .Z(new_n492));
  NOR2_X1   g306(.A1(new_n227), .A2(G119), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n236), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n233), .A2(new_n492), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n477), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n433), .A2(G107), .ZN(new_n498));
  OAI21_X1  g312(.A(G101), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n481), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n488), .A2(new_n490), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n471), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n488), .A2(KEYINPUT88), .A3(new_n490), .A4(new_n504), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n488), .A2(new_n490), .A3(new_n504), .A4(new_n471), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT6), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n490), .A2(new_n504), .ZN(new_n511));
  INV_X1    g325(.A(new_n481), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT4), .B1(new_n512), .B2(new_n485), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n479), .A2(new_n472), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n489), .B1(new_n515), .B2(new_n246), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n506), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n471), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n517), .A2(KEYINPUT6), .A3(new_n508), .A4(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n470), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G210), .B1(G237), .B2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n468), .B(new_n523), .Z(new_n524));
  XNOR2_X1  g338(.A(new_n471), .B(KEYINPUT8), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n228), .A2(new_n231), .A3(KEYINPUT5), .A4(new_n232), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n491), .B1(new_n494), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n527), .B2(new_n500), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n496), .B2(new_n500), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n530), .B2(new_n509), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n521), .A2(new_n522), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n522), .ZN(new_n533));
  INV_X1    g347(.A(new_n470), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n517), .A2(new_n508), .A3(new_n518), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n537), .B2(new_n519), .ZN(new_n538));
  INV_X1    g352(.A(new_n531), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n540), .A3(KEYINPUT89), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n542), .B(new_n533), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  OAI21_X1  g357(.A(G221), .B1(new_n398), .B2(G902), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT79), .Z(new_n545));
  INV_X1    g359(.A(new_n225), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT82), .B1(new_n194), .B2(new_n224), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT82), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(G128), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n189), .A2(new_n191), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n500), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n253), .B1(new_n481), .B2(new_n499), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n250), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT12), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n249), .B1(new_n482), .B2(new_n486), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n502), .A2(KEYINPUT10), .A3(new_n253), .A4(new_n503), .ZN(new_n558));
  INV_X1    g372(.A(new_n250), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT10), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n552), .B2(new_n500), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n481), .A2(new_n499), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n549), .A2(G128), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n548), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n551), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n225), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n500), .A2(new_n223), .A3(new_n225), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n250), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G140), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n346), .A2(G227), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n556), .A2(new_n562), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n250), .A2(KEYINPUT84), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT10), .B1(new_n563), .B2(new_n567), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n515), .B2(new_n249), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n582), .B2(new_n558), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n557), .A2(new_n558), .A3(new_n561), .A4(new_n580), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n575), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n571), .B1(new_n570), .B2(new_n250), .ZN(new_n587));
  AOI211_X1 g401(.A(KEYINPUT12), .B(new_n559), .C1(new_n568), .C2(new_n569), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n589), .A2(KEYINPUT85), .A3(new_n576), .A4(new_n562), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n289), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n556), .A2(new_n562), .A3(new_n572), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n575), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n596));
  INV_X1    g410(.A(new_n580), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n576), .A3(new_n584), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(G469), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(G469), .A2(G902), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n545), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n466), .A2(new_n541), .A3(new_n543), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n372), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(new_n480), .ZN(G3));
  AOI21_X1  g420(.A(new_n465), .B1(new_n532), .B2(new_n540), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n431), .A2(new_n434), .A3(new_n440), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n431), .A2(new_n450), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n434), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n454), .B1(new_n610), .B2(new_n414), .ZN(new_n611));
  INV_X1    g425(.A(new_n455), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n460), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT92), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n453), .A2(new_n455), .B1(G475), .B2(new_n459), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT92), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n403), .A2(KEYINPUT33), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n403), .A2(KEYINPUT33), .ZN(new_n620));
  OAI211_X1 g434(.A(G478), .B(new_n289), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n607), .A2(new_n624), .A3(new_n380), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n593), .A2(new_n602), .ZN(new_n626));
  INV_X1    g440(.A(new_n545), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n297), .A2(KEYINPUT31), .B1(new_n301), .B2(new_n286), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n290), .B1(new_n629), .B2(new_n300), .ZN(new_n630));
  INV_X1    g444(.A(G472), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n305), .B(new_n371), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n625), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND2_X1  g452(.A1(new_n607), .A2(new_n380), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n412), .A2(new_n616), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n634), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT35), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT95), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND4_X1  g458(.A1(new_n618), .A2(new_n464), .A3(new_n380), .A4(new_n413), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n628), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n359), .A2(new_n360), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n313), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n345), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n366), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n305), .B(new_n652), .C1(new_n630), .C2(new_n631), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n646), .A2(new_n543), .A3(new_n654), .A4(new_n541), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n376), .B1(new_n377), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n412), .A2(new_n616), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n628), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n311), .A2(new_n662), .A3(new_n607), .A4(new_n652), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NAND3_X1  g478(.A1(new_n615), .A2(new_n617), .A3(new_n412), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n465), .A3(new_n652), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT96), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n659), .B(KEYINPUT39), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n603), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n286), .B1(new_n277), .B2(new_n278), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n457), .B1(new_n282), .B2(new_n263), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n309), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n541), .A2(new_n543), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT38), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n190), .ZN(G45));
  NAND2_X1  g494(.A1(new_n621), .A2(new_n622), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n615), .A2(new_n617), .A3(new_n681), .A4(new_n660), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n628), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n311), .A2(new_n683), .A3(new_n607), .A4(new_n652), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  OR2_X1    g499(.A1(new_n592), .A2(KEYINPUT97), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n591), .A2(new_n289), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n686), .B1(new_n591), .B2(new_n289), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n687), .A2(new_n688), .A3(new_n545), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n311), .A2(new_n371), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n625), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT41), .B(G113), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  INV_X1    g507(.A(new_n371), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n640), .A2(new_n694), .A3(new_n379), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n311), .A2(new_n607), .A3(new_n689), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT98), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  INV_X1    g512(.A(new_n652), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n463), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n311), .A2(new_n607), .A3(new_n689), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NOR4_X1   g516(.A1(new_n665), .A2(new_n687), .A3(new_n688), .A4(new_n545), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n367), .A2(new_n369), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT99), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n648), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT99), .B1(new_n361), .B2(new_n370), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n708), .B(new_n305), .C1(new_n631), .C2(new_n630), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n703), .A2(new_n607), .A3(new_n710), .A4(new_n380), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n532), .A2(new_n540), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n689), .A3(new_n464), .ZN(new_n715));
  INV_X1    g529(.A(new_n682), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n654), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n653), .A2(new_n682), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n607), .A2(new_n719), .A3(KEYINPUT100), .A4(new_n689), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  XOR2_X1   g536(.A(new_n601), .B(KEYINPUT101), .Z(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n595), .B2(new_n599), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n599), .A2(new_n725), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n724), .B1(new_n728), .B2(G469), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n545), .B1(new_n729), .B2(new_n593), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n676), .A2(new_n464), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n311), .A2(new_n716), .A3(new_n708), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT42), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n293), .A2(KEYINPUT74), .A3(G472), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT74), .B1(new_n293), .B2(G472), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n694), .B1(new_n736), .B2(new_n309), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n465), .B1(new_n541), .B2(new_n543), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n738), .A3(new_n730), .A4(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT103), .B(G131), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G33));
  INV_X1    g557(.A(new_n661), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n737), .A2(new_n744), .A3(new_n738), .A4(new_n730), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NAND2_X1  g560(.A1(new_n595), .A2(new_n599), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n592), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n726), .A2(new_n727), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(new_n748), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT104), .B(new_n749), .C1(new_n750), .C2(new_n748), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n724), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n593), .B1(new_n755), .B2(KEYINPUT46), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n757), .B(new_n724), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n627), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n668), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n618), .A2(new_n681), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n305), .B1(new_n630), .B2(new_n631), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT43), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n652), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n738), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n761), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n206), .ZN(G39));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n759), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT47), .B(new_n627), .C1(new_n756), .C2(new_n758), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n676), .A2(new_n464), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n780), .A2(new_n371), .A3(new_n311), .A4(new_n682), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NAND2_X1  g597(.A1(new_n373), .A2(new_n346), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n309), .A2(new_n371), .A3(new_n376), .A4(new_n673), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n681), .B1(new_n615), .B2(new_n617), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n689), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT108), .B1(new_n738), .B2(new_n689), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n766), .A2(new_n376), .A3(new_n768), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n789), .B2(new_n790), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  INV_X1    g612(.A(new_n689), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n780), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n689), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(KEYINPUT109), .A3(new_n794), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n653), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n785), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n795), .A2(new_n796), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT109), .B1(new_n802), .B2(new_n794), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n654), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n791), .B(KEYINPUT110), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT112), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n766), .A2(new_n376), .A3(new_n710), .A4(new_n768), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n689), .A2(new_n465), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n677), .A3(KEYINPUT50), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT50), .B1(new_n813), .B2(new_n677), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n687), .A2(new_n688), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT106), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n777), .B(new_n778), .C1(new_n627), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n811), .A2(new_n780), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n805), .A2(new_n810), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n802), .A2(new_n624), .A3(new_n787), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n374), .C1(new_n715), .C2(new_n811), .ZN(new_n825));
  INV_X1    g639(.A(new_n708), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n736), .B2(new_n309), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n806), .B2(new_n807), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT48), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT48), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n830), .B(new_n827), .C1(new_n806), .C2(new_n807), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n465), .B(new_n665), .C1(new_n540), .C2(new_n532), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n652), .A2(new_n659), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT107), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n674), .A3(new_n730), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n721), .A2(new_n663), .A3(new_n684), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n663), .A2(new_n684), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n721), .A4(new_n836), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n701), .B(new_n655), .C1(new_n690), .C2(new_n625), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n413), .B1(new_n461), .B2(new_n462), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n615), .A2(new_n617), .A3(new_n623), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n379), .A2(new_n465), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n633), .A2(new_n848), .A3(new_n543), .A4(new_n541), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(new_n711), .C1(new_n372), .C2(new_n604), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n697), .A2(new_n844), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n413), .A2(new_n652), .A3(new_n616), .A4(new_n660), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n628), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n676), .A2(new_n311), .A3(new_n464), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n676), .A2(new_n464), .A3(new_n719), .A4(new_n730), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(new_n733), .A3(new_n740), .A4(new_n745), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n842), .A2(new_n860), .A3(KEYINPUT53), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n838), .A2(new_n841), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n843), .A2(new_n850), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n731), .A2(new_n372), .A3(new_n661), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n857), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n741), .A2(new_n864), .A3(new_n866), .A4(new_n697), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT54), .B1(new_n861), .B2(new_n868), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n823), .B(new_n832), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n814), .A2(new_n815), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n808), .A2(new_n809), .A3(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n873), .A2(KEYINPUT111), .B1(new_n820), .B2(new_n821), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n808), .A2(new_n809), .A3(new_n875), .A4(new_n872), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT51), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n784), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  OR4_X1    g692(.A1(new_n545), .A2(new_n762), .A3(new_n465), .A4(new_n826), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n674), .B(new_n879), .C1(new_n819), .C2(KEYINPUT49), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n880), .B(new_n677), .C1(KEYINPUT49), .C2(new_n819), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(KEYINPUT113), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(G75));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n842), .B2(new_n860), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n863), .A2(new_n867), .A3(new_n862), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n289), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n533), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n510), .A2(new_n520), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n534), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n521), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(KEYINPUT56), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n891), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n891), .B2(new_n892), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n373), .A2(G953), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT115), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(G51));
  NOR2_X1   g718(.A1(new_n869), .A2(new_n870), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n723), .B(KEYINPUT57), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(KEYINPUT116), .A3(new_n906), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n591), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n890), .A2(new_n753), .A3(new_n754), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(G54));
  NAND2_X1  g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT117), .Z(new_n915));
  AND2_X1   g729(.A1(new_n890), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n610), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n610), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n903), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n619), .A2(new_n620), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT118), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n902), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n922), .B2(new_n925), .ZN(G63));
  NAND2_X1  g741(.A1(new_n861), .A2(new_n868), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT119), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n933), .B(new_n930), .C1(new_n861), .C2(new_n868), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n650), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n931), .B1(new_n887), .B2(new_n888), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n928), .A2(KEYINPUT119), .A3(new_n931), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n364), .B(KEYINPUT120), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n935), .A2(new_n940), .A3(new_n902), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  INV_X1    g756(.A(new_n650), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n937), .B2(new_n938), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n944), .B2(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT61), .B1(new_n935), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n935), .A2(new_n940), .A3(new_n902), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(G66));
  INV_X1    g765(.A(G224), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n378), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT123), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n852), .B(KEYINPUT122), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n346), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n893), .B1(G898), .B2(new_n346), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n956), .B(new_n959), .ZN(G69));
  NOR2_X1   g774(.A1(new_n628), .A2(new_n760), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n737), .A2(new_n845), .A3(new_n961), .A4(new_n846), .ZN(new_n962));
  OAI22_X1  g776(.A1(new_n761), .A2(new_n773), .B1(new_n780), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n779), .B2(new_n781), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n839), .A2(new_n721), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n679), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  AOI21_X1  g781(.A(G953), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(new_n446), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n968), .A2(KEYINPUT126), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT126), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  NAND2_X1  g786(.A1(G900), .A2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n761), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n827), .A2(new_n833), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n774), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n965), .A2(new_n865), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n741), .A3(new_n782), .A4(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n970), .B(new_n973), .C1(new_n978), .C2(G953), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n971), .A2(new_n972), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n346), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n971), .A2(new_n983), .A3(new_n972), .A4(new_n979), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n978), .B2(new_n955), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n285), .A2(new_n263), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT127), .Z(new_n990));
  AND2_X1   g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n964), .A2(new_n967), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n987), .B1(new_n992), .B2(new_n955), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n671), .ZN(new_n994));
  INV_X1    g808(.A(new_n987), .ZN(new_n995));
  NOR4_X1   g809(.A1(new_n889), .A2(new_n671), .A3(new_n995), .A4(new_n989), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n991), .A2(new_n994), .A3(new_n903), .A4(new_n996), .ZN(G57));
endmodule


