

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763;

  XNOR2_X1 U369 ( .A(n459), .B(n569), .ZN(n611) );
  XNOR2_X2 U370 ( .A(n377), .B(KEYINPUT70), .ZN(n477) );
  XNOR2_X2 U371 ( .A(KEYINPUT69), .B(G131), .ZN(n377) );
  AND2_X1 U372 ( .A1(n615), .A2(n347), .ZN(n717) );
  NAND2_X1 U373 ( .A1(n407), .A2(n404), .ZN(n600) );
  AND2_X1 U374 ( .A1(n682), .A2(n374), .ZN(n684) );
  NOR2_X1 U375 ( .A1(n661), .A2(n660), .ZN(n665) );
  AND2_X1 U376 ( .A1(n685), .A2(n709), .ZN(n563) );
  AND2_X1 U377 ( .A1(n642), .A2(n350), .ZN(n460) );
  BUF_X1 U378 ( .A(n642), .Z(n347) );
  XNOR2_X1 U379 ( .A(n395), .B(n349), .ZN(n598) );
  AND2_X1 U380 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U381 ( .A(KEYINPUT44), .ZN(n366) );
  XNOR2_X1 U382 ( .A(n600), .B(KEYINPUT1), .ZN(n642) );
  XNOR2_X1 U383 ( .A(G143), .B(G128), .ZN(n467) );
  NAND2_X2 U384 ( .A1(n383), .A2(n381), .ZN(n628) );
  AND2_X1 U385 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X1 U386 ( .A(n457), .B(n421), .ZN(n676) );
  XNOR2_X1 U387 ( .A(G119), .B(G113), .ZN(n453) );
  XNOR2_X1 U388 ( .A(n588), .B(KEYINPUT79), .ZN(n589) );
  XNOR2_X1 U389 ( .A(n380), .B(n379), .ZN(n378) );
  OR2_X1 U390 ( .A1(n632), .A2(KEYINPUT47), .ZN(n616) );
  AND2_X1 U391 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U392 ( .A1(n392), .A2(n391), .ZN(n390) );
  NOR2_X1 U393 ( .A1(n393), .A2(n717), .ZN(n392) );
  INV_X1 U394 ( .A(n394), .ZN(n393) );
  AND2_X1 U395 ( .A1(n516), .A2(n515), .ZN(n517) );
  AND2_X1 U396 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U397 ( .A(KEYINPUT96), .B(KEYINPUT17), .ZN(n492) );
  XNOR2_X1 U398 ( .A(n376), .B(n495), .ZN(n750) );
  XNOR2_X1 U399 ( .A(n477), .B(G134), .ZN(n376) );
  XNOR2_X1 U400 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n534) );
  XNOR2_X1 U401 ( .A(n483), .B(n361), .ZN(n485) );
  XNOR2_X1 U402 ( .A(n484), .B(n362), .ZN(n361) );
  XNOR2_X1 U403 ( .A(n502), .B(n744), .ZN(n720) );
  NAND2_X1 U404 ( .A1(n628), .A2(n643), .ZN(n613) );
  OR2_X1 U405 ( .A1(n676), .A2(n405), .ZN(n404) );
  NAND2_X1 U406 ( .A1(n406), .A2(n504), .ZN(n405) );
  OR2_X2 U407 ( .A1(n566), .A2(n556), .ZN(n396) );
  AND2_X2 U408 ( .A1(n675), .A2(n674), .ZN(n730) );
  NAND2_X1 U409 ( .A1(n372), .A2(n370), .ZN(n369) );
  NOR2_X1 U410 ( .A1(n371), .A2(n736), .ZN(n370) );
  NAND2_X1 U411 ( .A1(n730), .A2(n358), .ZN(n372) );
  NOR2_X1 U412 ( .A1(n357), .A2(G475), .ZN(n371) );
  NAND2_X1 U413 ( .A1(n627), .A2(n626), .ZN(n394) );
  AND2_X1 U414 ( .A1(n638), .A2(n713), .ZN(n632) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n476) );
  XNOR2_X1 U416 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U417 ( .A(n750), .B(G146), .ZN(n457) );
  XNOR2_X1 U418 ( .A(n402), .B(n401), .ZN(n464) );
  INV_X1 U419 ( .A(KEYINPUT8), .ZN(n401) );
  XNOR2_X1 U420 ( .A(G143), .B(G104), .ZN(n484) );
  INV_X1 U421 ( .A(G140), .ZN(n362) );
  XNOR2_X1 U422 ( .A(G113), .B(G122), .ZN(n481) );
  XOR2_X1 U423 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n482) );
  XNOR2_X1 U424 ( .A(KEYINPUT18), .B(KEYINPUT83), .ZN(n489) );
  XNOR2_X1 U425 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n375) );
  NAND2_X1 U426 ( .A1(n651), .A2(n650), .ZN(n663) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n661) );
  INV_X1 U428 ( .A(KEYINPUT45), .ZN(n363) );
  NAND2_X1 U429 ( .A1(n598), .A2(n643), .ZN(n380) );
  INV_X1 U430 ( .A(KEYINPUT30), .ZN(n379) );
  OR2_X2 U431 ( .A1(n692), .A2(G902), .ZN(n395) );
  NAND2_X1 U432 ( .A1(n423), .A2(G902), .ZN(n408) );
  XNOR2_X1 U433 ( .A(G104), .B(G107), .ZN(n419) );
  INV_X1 U434 ( .A(G107), .ZN(n468) );
  BUF_X1 U435 ( .A(n663), .Z(n755) );
  XNOR2_X1 U436 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U437 ( .A(n705), .B(n360), .ZN(n638) );
  INV_X1 U438 ( .A(KEYINPUT101), .ZN(n360) );
  XNOR2_X1 U439 ( .A(n613), .B(KEYINPUT19), .ZN(n618) );
  XNOR2_X1 U440 ( .A(KEYINPUT16), .B(G122), .ZN(n500) );
  NAND2_X1 U441 ( .A1(n730), .A2(G469), .ZN(n680) );
  XNOR2_X1 U442 ( .A(n592), .B(KEYINPUT40), .ZN(n690) );
  XNOR2_X1 U443 ( .A(n367), .B(n559), .ZN(n685) );
  NOR2_X1 U444 ( .A1(n629), .A2(n648), .ZN(n630) );
  NOR2_X1 U445 ( .A1(n373), .A2(n369), .ZN(n729) );
  NOR2_X1 U446 ( .A1(n730), .A2(n357), .ZN(n373) );
  AND2_X1 U447 ( .A1(n596), .A2(n354), .ZN(n348) );
  XOR2_X1 U448 ( .A(n560), .B(KEYINPUT102), .Z(n349) );
  XNOR2_X1 U449 ( .A(n467), .B(n375), .ZN(n495) );
  AND2_X1 U450 ( .A1(n596), .A2(n594), .ZN(n350) );
  XNOR2_X1 U451 ( .A(n397), .B(KEYINPUT0), .ZN(n566) );
  XOR2_X1 U452 ( .A(n607), .B(KEYINPUT46), .Z(n351) );
  AND2_X1 U453 ( .A1(n550), .A2(n549), .ZN(n352) );
  AND2_X1 U454 ( .A1(n546), .A2(n583), .ZN(n353) );
  NOR2_X1 U455 ( .A1(n593), .A2(n403), .ZN(n354) );
  AND2_X1 U456 ( .A1(n577), .A2(n701), .ZN(n355) );
  XOR2_X1 U457 ( .A(KEYINPUT94), .B(KEYINPUT39), .Z(n356) );
  XOR2_X1 U458 ( .A(n727), .B(n726), .Z(n357) );
  AND2_X1 U459 ( .A1(n357), .A2(G475), .ZN(n358) );
  INV_X1 U460 ( .A(n736), .ZN(n374) );
  XNOR2_X1 U461 ( .A(n359), .B(n637), .ZN(n651) );
  NAND2_X1 U462 ( .A1(n636), .A2(n351), .ZN(n359) );
  NAND2_X1 U463 ( .A1(n526), .A2(n550), .ZN(n705) );
  XNOR2_X1 U464 ( .A(n565), .B(n366), .ZN(n365) );
  NAND2_X1 U465 ( .A1(n365), .A2(n355), .ZN(n364) );
  NAND2_X1 U466 ( .A1(n575), .A2(n558), .ZN(n367) );
  XNOR2_X2 U467 ( .A(n396), .B(n557), .ZN(n575) );
  NAND2_X1 U468 ( .A1(n368), .A2(n394), .ZN(n389) );
  AND2_X1 U469 ( .A1(n368), .A2(KEYINPUT72), .ZN(n391) );
  XNOR2_X1 U470 ( .A(n634), .B(KEYINPUT87), .ZN(n368) );
  NAND2_X1 U471 ( .A1(n589), .A2(n378), .ZN(n629) );
  NAND2_X1 U472 ( .A1(n720), .A2(n506), .ZN(n385) );
  OR2_X1 U473 ( .A1(n720), .A2(n382), .ZN(n381) );
  OR2_X1 U474 ( .A1(n506), .A2(n667), .ZN(n382) );
  NAND2_X1 U475 ( .A1(n506), .A2(n667), .ZN(n384) );
  NAND2_X1 U476 ( .A1(n390), .A2(n386), .ZN(n636) );
  NAND2_X1 U477 ( .A1(n717), .A2(n635), .ZN(n387) );
  NAND2_X1 U478 ( .A1(n389), .A2(n635), .ZN(n388) );
  XNOR2_X2 U479 ( .A(n395), .B(G472), .ZN(n569) );
  NAND2_X1 U480 ( .A1(n618), .A2(n353), .ZN(n397) );
  NAND2_X1 U481 ( .A1(n400), .A2(n398), .ZN(n592) );
  INV_X1 U482 ( .A(n713), .ZN(n398) );
  NAND2_X1 U483 ( .A1(n400), .A2(n399), .ZN(n640) );
  INV_X1 U484 ( .A(n638), .ZN(n399) );
  XNOR2_X1 U485 ( .A(n591), .B(n356), .ZN(n400) );
  NAND2_X1 U486 ( .A1(n756), .A2(G234), .ZN(n402) );
  INV_X4 U487 ( .A(G953), .ZN(n756) );
  NAND2_X1 U488 ( .A1(n600), .A2(n350), .ZN(n587) );
  NAND2_X1 U489 ( .A1(n600), .A2(n348), .ZN(n588) );
  INV_X1 U490 ( .A(n594), .ZN(n403) );
  XNOR2_X2 U491 ( .A(n439), .B(n438), .ZN(n596) );
  INV_X1 U492 ( .A(n423), .ZN(n406) );
  NAND2_X1 U493 ( .A1(n676), .A2(n423), .ZN(n409) );
  XNOR2_X2 U494 ( .A(n410), .B(KEYINPUT35), .ZN(n761) );
  NAND2_X1 U495 ( .A1(n411), .A2(n352), .ZN(n410) );
  XNOR2_X1 U496 ( .A(n412), .B(n548), .ZN(n411) );
  NAND2_X1 U497 ( .A1(n414), .A2(n413), .ZN(n412) );
  INV_X1 U498 ( .A(n566), .ZN(n413) );
  INV_X1 U499 ( .A(n547), .ZN(n414) );
  NOR2_X2 U500 ( .A1(n695), .A2(n736), .ZN(n697) );
  NOR2_X2 U501 ( .A1(n723), .A2(n736), .ZN(n725) );
  NOR2_X1 U502 ( .A1(n713), .A2(n609), .ZN(n610) );
  XNOR2_X1 U503 ( .A(n680), .B(n679), .ZN(n682) );
  XNOR2_X1 U504 ( .A(n663), .B(n662), .ZN(n664) );
  AND2_X1 U505 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U506 ( .A1(n620), .A2(n624), .ZN(n621) );
  XNOR2_X1 U507 ( .A(n518), .B(KEYINPUT51), .ZN(n519) );
  INV_X1 U508 ( .A(KEYINPUT72), .ZN(n635) );
  INV_X1 U509 ( .A(KEYINPUT77), .ZN(n449) );
  INV_X1 U510 ( .A(KEYINPUT78), .ZN(n662) );
  INV_X1 U511 ( .A(n608), .ZN(n609) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n420), .B(n497), .ZN(n421) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT103), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U517 ( .A(G472), .ZN(n560) );
  XNOR2_X1 U518 ( .A(n471), .B(n470), .ZN(n473) );
  INV_X1 U519 ( .A(KEYINPUT125), .ZN(n731) );
  XNOR2_X1 U520 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U521 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U522 ( .A(n659), .B(n658), .ZN(G75) );
  XNOR2_X1 U523 ( .A(KEYINPUT71), .B(G140), .ZN(n415) );
  XNOR2_X1 U524 ( .A(n415), .B(G137), .ZN(n424) );
  NAND2_X1 U525 ( .A1(G227), .A2(n756), .ZN(n416) );
  XOR2_X1 U526 ( .A(n416), .B(KEYINPUT82), .Z(n417) );
  XNOR2_X1 U527 ( .A(n424), .B(n417), .ZN(n420) );
  INV_X1 U528 ( .A(G110), .ZN(n418) );
  XNOR2_X1 U529 ( .A(n419), .B(n418), .ZN(n742) );
  XNOR2_X1 U530 ( .A(KEYINPUT67), .B(G101), .ZN(n450) );
  XNOR2_X1 U531 ( .A(n742), .B(n450), .ZN(n497) );
  INV_X1 U532 ( .A(KEYINPUT73), .ZN(n422) );
  XNOR2_X1 U533 ( .A(n422), .B(G469), .ZN(n423) );
  XNOR2_X2 U534 ( .A(G146), .B(G125), .ZN(n490) );
  XNOR2_X1 U535 ( .A(n490), .B(KEYINPUT10), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(n424), .ZN(n749) );
  XOR2_X1 U537 ( .A(KEYINPUT23), .B(G110), .Z(n426) );
  NAND2_X1 U538 ( .A1(n464), .A2(G221), .ZN(n425) );
  XNOR2_X1 U539 ( .A(n426), .B(n425), .ZN(n430) );
  XNOR2_X1 U540 ( .A(G119), .B(G128), .ZN(n427) );
  XNOR2_X1 U541 ( .A(KEYINPUT81), .B(n427), .ZN(n428) );
  XNOR2_X1 U542 ( .A(n428), .B(KEYINPUT24), .ZN(n429) );
  XNOR2_X1 U543 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U544 ( .A(n749), .B(n431), .ZN(n699) );
  INV_X1 U545 ( .A(G902), .ZN(n504) );
  NAND2_X1 U546 ( .A1(n699), .A2(n504), .ZN(n439) );
  INV_X1 U547 ( .A(KEYINPUT15), .ZN(n432) );
  XNOR2_X1 U548 ( .A(n432), .B(G902), .ZN(n667) );
  INV_X1 U549 ( .A(n667), .ZN(n660) );
  NAND2_X1 U550 ( .A1(n660), .A2(G234), .ZN(n434) );
  XOR2_X1 U551 ( .A(KEYINPUT20), .B(KEYINPUT99), .Z(n433) );
  XNOR2_X1 U552 ( .A(n434), .B(n433), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n440), .A2(G217), .ZN(n437) );
  INV_X1 U554 ( .A(KEYINPUT80), .ZN(n435) );
  XNOR2_X1 U555 ( .A(n435), .B(KEYINPUT25), .ZN(n436) );
  XNOR2_X1 U556 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U557 ( .A1(n440), .A2(G221), .ZN(n442) );
  INV_X1 U558 ( .A(KEYINPUT21), .ZN(n441) );
  XNOR2_X1 U559 ( .A(n442), .B(n441), .ZN(n594) );
  INV_X1 U560 ( .A(KEYINPUT6), .ZN(n459) );
  INV_X1 U561 ( .A(KEYINPUT5), .ZN(n443) );
  NAND2_X1 U562 ( .A1(G137), .A2(n443), .ZN(n446) );
  INV_X1 U563 ( .A(G137), .ZN(n444) );
  NAND2_X1 U564 ( .A1(n444), .A2(KEYINPUT5), .ZN(n445) );
  NAND2_X1 U565 ( .A1(n446), .A2(n445), .ZN(n448) );
  NAND2_X1 U566 ( .A1(n476), .A2(G210), .ZN(n447) );
  XNOR2_X1 U567 ( .A(n448), .B(n447), .ZN(n452) );
  XNOR2_X1 U568 ( .A(n453), .B(KEYINPUT3), .ZN(n455) );
  XNOR2_X1 U569 ( .A(G116), .B(KEYINPUT74), .ZN(n454) );
  XNOR2_X1 U570 ( .A(n455), .B(n454), .ZN(n501) );
  XOR2_X1 U571 ( .A(n456), .B(n501), .Z(n458) );
  XNOR2_X1 U572 ( .A(n458), .B(n457), .ZN(n692) );
  NAND2_X1 U573 ( .A1(n460), .A2(n611), .ZN(n463) );
  XOR2_X1 U574 ( .A(KEYINPUT33), .B(KEYINPUT95), .Z(n461) );
  XNOR2_X1 U575 ( .A(n463), .B(n462), .ZN(n547) );
  BUF_X1 U576 ( .A(n547), .Z(n530) );
  NAND2_X1 U577 ( .A1(n464), .A2(G217), .ZN(n466) );
  XOR2_X1 U578 ( .A(G134), .B(KEYINPUT7), .Z(n465) );
  XNOR2_X1 U579 ( .A(n466), .B(n465), .ZN(n471) );
  XOR2_X1 U580 ( .A(n467), .B(G116), .Z(n469) );
  XOR2_X1 U581 ( .A(G122), .B(KEYINPUT9), .Z(n472) );
  XNOR2_X1 U582 ( .A(n473), .B(n472), .ZN(n732) );
  NOR2_X1 U583 ( .A1(n732), .A2(G902), .ZN(n475) );
  XOR2_X1 U584 ( .A(KEYINPUT100), .B(G478), .Z(n474) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n550) );
  AND2_X1 U586 ( .A1(n476), .A2(G214), .ZN(n478) );
  XNOR2_X1 U587 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U588 ( .A(n480), .B(n479), .ZN(n486) );
  XNOR2_X1 U589 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U590 ( .A(n486), .B(n485), .Z(n727) );
  NOR2_X1 U591 ( .A1(G902), .A2(n727), .ZN(n488) );
  XNOR2_X1 U592 ( .A(KEYINPUT13), .B(G475), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n549) );
  OR2_X1 U594 ( .A1(n550), .A2(n549), .ZN(n554) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n494) );
  NAND2_X1 U596 ( .A1(n756), .A2(G224), .ZN(n491) );
  XNOR2_X1 U597 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n496) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n499) );
  INV_X1 U600 ( .A(n497), .ZN(n498) );
  XNOR2_X1 U601 ( .A(n499), .B(n498), .ZN(n502) );
  XNOR2_X1 U602 ( .A(n501), .B(n500), .ZN(n744) );
  INV_X1 U603 ( .A(G237), .ZN(n503) );
  NAND2_X1 U604 ( .A1(n504), .A2(n503), .ZN(n507) );
  NAND2_X1 U605 ( .A1(n507), .A2(G210), .ZN(n505) );
  XNOR2_X1 U606 ( .A(n505), .B(KEYINPUT85), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n628), .B(KEYINPUT38), .ZN(n590) );
  INV_X1 U608 ( .A(n590), .ZN(n523) );
  NAND2_X1 U609 ( .A1(n507), .A2(G214), .ZN(n643) );
  NAND2_X1 U610 ( .A1(n523), .A2(n643), .ZN(n527) );
  NOR2_X1 U611 ( .A1(n554), .A2(n527), .ZN(n508) );
  XNOR2_X1 U612 ( .A(KEYINPUT41), .B(n508), .ZN(n602) );
  NOR2_X1 U613 ( .A1(n530), .A2(n602), .ZN(n541) );
  NAND2_X1 U614 ( .A1(n569), .A2(n350), .ZN(n509) );
  INV_X1 U615 ( .A(n347), .ZN(n573) );
  NOR2_X1 U616 ( .A1(n509), .A2(n573), .ZN(n567) );
  OR2_X1 U617 ( .A1(n347), .A2(n350), .ZN(n510) );
  XNOR2_X1 U618 ( .A(n510), .B(KEYINPUT50), .ZN(n516) );
  NOR2_X1 U619 ( .A1(n596), .A2(n594), .ZN(n511) );
  XOR2_X1 U620 ( .A(KEYINPUT115), .B(n511), .Z(n512) );
  XNOR2_X1 U621 ( .A(KEYINPUT49), .B(n512), .ZN(n514) );
  INV_X1 U622 ( .A(n569), .ZN(n513) );
  NOR2_X1 U623 ( .A1(n567), .A2(n517), .ZN(n520) );
  INV_X1 U624 ( .A(KEYINPUT116), .ZN(n518) );
  NOR2_X1 U625 ( .A1(n602), .A2(n521), .ZN(n522) );
  XOR2_X1 U626 ( .A(KEYINPUT117), .B(n522), .Z(n533) );
  NOR2_X1 U627 ( .A1(n523), .A2(n643), .ZN(n524) );
  NOR2_X1 U628 ( .A1(n554), .A2(n524), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n525), .B(KEYINPUT118), .ZN(n529) );
  INV_X1 U630 ( .A(n549), .ZN(n526) );
  OR2_X1 U631 ( .A1(n550), .A2(n526), .ZN(n713) );
  NOR2_X1 U632 ( .A1(n527), .A2(n632), .ZN(n528) );
  NOR2_X1 U633 ( .A1(n529), .A2(n528), .ZN(n531) );
  NOR2_X1 U634 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U635 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U636 ( .A1(n536), .A2(G952), .ZN(n539) );
  NAND2_X1 U637 ( .A1(G237), .A2(G234), .ZN(n537) );
  XNOR2_X1 U638 ( .A(n537), .B(KEYINPUT14), .ZN(n583) );
  INV_X1 U639 ( .A(n583), .ZN(n538) );
  NOR2_X1 U640 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U641 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U642 ( .A(n542), .B(KEYINPUT120), .ZN(n543) );
  NAND2_X1 U643 ( .A1(n543), .A2(n756), .ZN(n656) );
  NOR2_X1 U644 ( .A1(G898), .A2(n756), .ZN(n544) );
  XNOR2_X1 U645 ( .A(KEYINPUT98), .B(n544), .ZN(n745) );
  NAND2_X1 U646 ( .A1(n745), .A2(G902), .ZN(n545) );
  NAND2_X1 U647 ( .A1(n756), .A2(G952), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n545), .A2(n581), .ZN(n546) );
  INV_X1 U649 ( .A(KEYINPUT34), .ZN(n548) );
  INV_X1 U650 ( .A(n761), .ZN(n564) );
  XNOR2_X1 U651 ( .A(n611), .B(KEYINPUT84), .ZN(n553) );
  INV_X1 U652 ( .A(n596), .ZN(n551) );
  NAND2_X1 U653 ( .A1(n347), .A2(n551), .ZN(n552) );
  NOR2_X1 U654 ( .A1(n553), .A2(n552), .ZN(n558) );
  INV_X1 U655 ( .A(n554), .ZN(n555) );
  NAND2_X1 U656 ( .A1(n555), .A2(n594), .ZN(n556) );
  XNOR2_X1 U657 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n557) );
  XNOR2_X1 U658 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n559) );
  OR2_X1 U659 ( .A1(n347), .A2(n596), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n598), .A2(n561), .ZN(n562) );
  NAND2_X1 U661 ( .A1(n562), .A2(n575), .ZN(n709) );
  NAND2_X1 U662 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U663 ( .A1(n567), .A2(n413), .ZN(n568) );
  XOR2_X1 U664 ( .A(KEYINPUT31), .B(n568), .Z(n715) );
  NOR2_X1 U665 ( .A1(n569), .A2(n587), .ZN(n570) );
  NAND2_X1 U666 ( .A1(n413), .A2(n570), .ZN(n706) );
  NAND2_X1 U667 ( .A1(n715), .A2(n706), .ZN(n572) );
  INV_X1 U668 ( .A(n632), .ZN(n571) );
  NAND2_X1 U669 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U670 ( .A1(n573), .A2(n596), .ZN(n574) );
  NOR2_X1 U671 ( .A1(n611), .A2(n574), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n701) );
  INV_X1 U673 ( .A(n661), .ZN(n737) );
  NAND2_X1 U674 ( .A1(G902), .A2(n583), .ZN(n578) );
  NOR2_X1 U675 ( .A1(G900), .A2(n578), .ZN(n579) );
  NAND2_X1 U676 ( .A1(G953), .A2(n579), .ZN(n580) );
  XOR2_X1 U677 ( .A(KEYINPUT104), .B(n580), .Z(n585) );
  INV_X1 U678 ( .A(n581), .ZN(n582) );
  AND2_X1 U679 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U680 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U681 ( .A(n586), .B(KEYINPUT86), .ZN(n593) );
  NOR2_X1 U682 ( .A1(n629), .A2(n590), .ZN(n591) );
  INV_X1 U683 ( .A(n593), .ZN(n595) );
  NAND2_X1 U684 ( .A1(n595), .A2(n594), .ZN(n597) );
  NOR2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n608) );
  AND2_X1 U686 ( .A1(n598), .A2(n608), .ZN(n599) );
  XNOR2_X1 U687 ( .A(KEYINPUT28), .B(n599), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n601), .A2(n600), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n602), .A2(n617), .ZN(n605) );
  INV_X1 U690 ( .A(KEYINPUT109), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n603), .B(KEYINPUT42), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n605), .B(n604), .ZN(n763) );
  INV_X1 U693 ( .A(n763), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n690), .A2(n606), .ZN(n607) );
  XNOR2_X1 U695 ( .A(KEYINPUT105), .B(n612), .ZN(n641) );
  NOR2_X1 U696 ( .A1(n641), .A2(n613), .ZN(n614) );
  XNOR2_X1 U697 ( .A(n614), .B(KEYINPUT36), .ZN(n615) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT76), .ZN(n622) );
  INV_X1 U699 ( .A(n617), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n623) );
  INV_X1 U701 ( .A(n623), .ZN(n620) );
  INV_X1 U702 ( .A(KEYINPUT89), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n627) );
  XOR2_X1 U704 ( .A(n624), .B(KEYINPUT47), .Z(n625) );
  NAND2_X1 U705 ( .A1(n623), .A2(n625), .ZN(n626) );
  INV_X1 U706 ( .A(n628), .ZN(n648) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT108), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n631), .A2(n352), .ZN(n689) );
  NAND2_X1 U709 ( .A1(n632), .A2(KEYINPUT47), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n689), .A2(n633), .ZN(n634) );
  XNOR2_X1 U711 ( .A(KEYINPUT93), .B(KEYINPUT48), .ZN(n637) );
  INV_X1 U712 ( .A(KEYINPUT110), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n762) );
  XOR2_X1 U714 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n646) );
  NOR2_X1 U715 ( .A1(n347), .A2(n641), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT43), .ZN(n649) );
  AND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n687) );
  NOR2_X1 U720 ( .A1(n762), .A2(n687), .ZN(n650) );
  INV_X1 U721 ( .A(n755), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n737), .A2(n652), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n653), .A2(KEYINPUT88), .ZN(n654) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n672) );
  XNOR2_X1 U725 ( .A(n654), .B(n672), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n659) );
  INV_X1 U727 ( .A(KEYINPUT53), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT121), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U730 ( .A(n666), .B(KEYINPUT90), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n667), .B(KEYINPUT91), .ZN(n668) );
  NOR2_X1 U732 ( .A1(n668), .A2(n672), .ZN(n669) );
  XNOR2_X1 U733 ( .A(n669), .B(KEYINPUT65), .ZN(n670) );
  NAND2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U735 ( .A1(n755), .A2(n672), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n737), .A2(n673), .ZN(n674) );
  XNOR2_X1 U737 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n678) );
  XNOR2_X1 U738 ( .A(n676), .B(KEYINPUT57), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n678), .B(n677), .ZN(n679) );
  INV_X1 U740 ( .A(G952), .ZN(n681) );
  AND2_X1 U741 ( .A1(n681), .A2(G953), .ZN(n736) );
  INV_X1 U742 ( .A(KEYINPUT123), .ZN(n683) );
  XNOR2_X1 U743 ( .A(n684), .B(n683), .ZN(G54) );
  XNOR2_X1 U744 ( .A(n685), .B(G119), .ZN(G21) );
  XNOR2_X1 U745 ( .A(G140), .B(KEYINPUT114), .ZN(n686) );
  XOR2_X1 U746 ( .A(n687), .B(n686), .Z(G42) );
  XOR2_X1 U747 ( .A(G143), .B(KEYINPUT113), .Z(n688) );
  XNOR2_X1 U748 ( .A(n689), .B(n688), .ZN(G45) );
  XNOR2_X1 U749 ( .A(n690), .B(G131), .ZN(G33) );
  NAND2_X1 U750 ( .A1(n730), .A2(G472), .ZN(n694) );
  XOR2_X1 U751 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n691) );
  XNOR2_X1 U752 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U753 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U754 ( .A(KEYINPUT97), .B(KEYINPUT63), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n697), .B(n696), .ZN(G57) );
  NAND2_X1 U756 ( .A1(n730), .A2(G217), .ZN(n698) );
  XOR2_X1 U757 ( .A(n699), .B(n698), .Z(n700) );
  NOR2_X1 U758 ( .A1(n700), .A2(n736), .ZN(G66) );
  XNOR2_X1 U759 ( .A(G101), .B(n701), .ZN(G3) );
  NOR2_X1 U760 ( .A1(n706), .A2(n713), .ZN(n702) );
  XOR2_X1 U761 ( .A(G104), .B(n702), .Z(G6) );
  XOR2_X1 U762 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n704) );
  XNOR2_X1 U763 ( .A(G107), .B(KEYINPUT112), .ZN(n703) );
  XNOR2_X1 U764 ( .A(n704), .B(n703), .ZN(n708) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U766 ( .A(n708), .B(n707), .Z(G9) );
  XNOR2_X1 U767 ( .A(G110), .B(n709), .ZN(G12) );
  NOR2_X1 U768 ( .A1(n623), .A2(n705), .ZN(n711) );
  XNOR2_X1 U769 ( .A(G128), .B(KEYINPUT29), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(G30) );
  NOR2_X1 U771 ( .A1(n623), .A2(n713), .ZN(n712) );
  XOR2_X1 U772 ( .A(G146), .B(n712), .Z(G48) );
  NOR2_X1 U773 ( .A1(n713), .A2(n715), .ZN(n714) );
  XOR2_X1 U774 ( .A(G113), .B(n714), .Z(G15) );
  NOR2_X1 U775 ( .A1(n705), .A2(n715), .ZN(n716) );
  XOR2_X1 U776 ( .A(G116), .B(n716), .Z(G18) );
  XNOR2_X1 U777 ( .A(G125), .B(n717), .ZN(n718) );
  XNOR2_X1 U778 ( .A(n718), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U779 ( .A1(n730), .A2(G210), .ZN(n722) );
  XOR2_X1 U780 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n719) );
  XNOR2_X1 U781 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U783 ( .A(KEYINPUT92), .B(KEYINPUT56), .ZN(n724) );
  XNOR2_X1 U784 ( .A(n725), .B(n724), .ZN(G51) );
  XOR2_X1 U785 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n726) );
  XNOR2_X1 U786 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n728) );
  XNOR2_X1 U787 ( .A(n729), .B(n728), .ZN(G60) );
  NAND2_X1 U788 ( .A1(n730), .A2(G478), .ZN(n734) );
  NOR2_X1 U789 ( .A1(n736), .A2(n735), .ZN(G63) );
  NAND2_X1 U790 ( .A1(n737), .A2(n756), .ZN(n741) );
  NAND2_X1 U791 ( .A1(G953), .A2(G224), .ZN(n738) );
  XNOR2_X1 U792 ( .A(KEYINPUT61), .B(n738), .ZN(n739) );
  NAND2_X1 U793 ( .A1(n739), .A2(G898), .ZN(n740) );
  NAND2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n748) );
  XOR2_X1 U795 ( .A(G101), .B(n742), .Z(n743) );
  XNOR2_X1 U796 ( .A(n744), .B(n743), .ZN(n746) );
  NOR2_X1 U797 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(G69) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(n754) );
  XOR2_X1 U800 ( .A(G227), .B(n754), .Z(n751) );
  NAND2_X1 U801 ( .A1(n751), .A2(G900), .ZN(n752) );
  XOR2_X1 U802 ( .A(KEYINPUT126), .B(n752), .Z(n753) );
  NAND2_X1 U803 ( .A1(G953), .A2(n753), .ZN(n759) );
  XNOR2_X1 U804 ( .A(n755), .B(n754), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n760), .B(KEYINPUT127), .ZN(G72) );
  XOR2_X1 U808 ( .A(n761), .B(G122), .Z(G24) );
  XOR2_X1 U809 ( .A(G134), .B(n762), .Z(G36) );
  XOR2_X1 U810 ( .A(n763), .B(G137), .Z(G39) );
endmodule

