//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT79), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n192), .B(G119), .C1(KEYINPUT77), .C2(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n195), .B2(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n199), .A2(G110), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(KEYINPUT78), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(KEYINPUT78), .ZN(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT76), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n201), .B(new_n202), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(G125), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(G146), .B(new_n209), .C1(new_n213), .C2(new_n207), .ZN(new_n214));
  INV_X1    g028(.A(new_n213), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n205), .A2(new_n203), .B1(G110), .B2(new_n199), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n209), .B1(new_n213), .B2(new_n207), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n214), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n218), .A2(KEYINPUT80), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT80), .B1(new_n218), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n191), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(new_n191), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT25), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(G234), .B2(new_n229), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G902), .ZN(new_n237));
  XOR2_X1   g051(.A(new_n237), .B(KEYINPUT81), .Z(new_n238));
  AND2_X1   g052(.A1(new_n227), .A2(new_n228), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n234), .A2(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(G134), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G137), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT66), .B(new_n244), .C1(new_n245), .C2(G137), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n243), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT67), .B(G137), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT11), .A2(G134), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G137), .ZN(new_n258));
  AND4_X1   g072(.A1(new_n252), .A2(new_n256), .A3(new_n258), .A4(new_n254), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n250), .B(new_n251), .C1(new_n255), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n263), .A3(G143), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n221), .A2(G143), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n192), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n261), .A2(new_n263), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n253), .A2(G134), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n245), .A2(G137), .ZN(new_n276));
  OAI21_X1  g090(.A(G131), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n260), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n271), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(new_n216), .B2(G143), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n265), .B1(new_n216), .B2(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n283), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n256), .A2(new_n258), .A3(new_n254), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n256), .A2(new_n258), .A3(new_n254), .A4(new_n252), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n293), .A2(new_n251), .A3(new_n250), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n251), .B1(new_n293), .B2(new_n250), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n260), .A2(new_n274), .A3(KEYINPUT71), .A4(new_n277), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n280), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n195), .A2(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(KEYINPUT2), .A2(G113), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g119(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n302), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n308), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n280), .A2(new_n296), .A3(new_n310), .A4(new_n297), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n310), .A3(new_n278), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n187), .A3(G210), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT27), .Z(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G101), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n313), .A2(new_n319), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n280), .A2(new_n296), .A3(KEYINPUT30), .A4(new_n297), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n286), .A2(new_n288), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n255), .A2(new_n259), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n248), .A2(new_n249), .ZN(new_n333));
  INV_X1    g147(.A(new_n243), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G131), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n331), .B1(new_n336), .B2(new_n260), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n260), .A2(new_n274), .A3(new_n277), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n339), .A3(new_n308), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n340), .A2(new_n324), .A3(new_n311), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n310), .B1(new_n296), .B2(new_n278), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n316), .B2(new_n314), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n296), .A2(new_n297), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n344), .A2(KEYINPUT28), .A3(new_n310), .A4(new_n280), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n324), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n325), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n313), .A2(new_n319), .A3(new_n348), .A4(new_n326), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n328), .A2(new_n347), .A3(new_n229), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G472), .ZN(new_n351));
  INV_X1    g165(.A(new_n324), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n340), .A2(new_n352), .A3(new_n311), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT31), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n314), .A2(new_n316), .ZN(new_n358));
  INV_X1    g172(.A(new_n342), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n311), .A2(new_n316), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n324), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n340), .A2(new_n352), .A3(new_n311), .A4(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT32), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT32), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n351), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n350), .B2(G472), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT75), .A3(new_n368), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n241), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n274), .A2(new_n211), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n211), .B2(new_n331), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT86), .B(G224), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n187), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT7), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n378), .B(new_n381), .Z(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n383), .A2(KEYINPUT3), .A3(G107), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT82), .B(G104), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(G113), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n300), .A2(KEYINPUT5), .A3(new_n301), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n307), .B2(new_n302), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n394), .B1(new_n399), .B2(KEYINPUT88), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(KEYINPUT88), .B2(new_n399), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G122), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n402), .B(KEYINPUT8), .Z(new_n403));
  NOR2_X1   g217(.A1(new_n302), .A2(new_n307), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(KEYINPUT85), .A3(new_n396), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n403), .B1(new_n408), .B2(new_n394), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n382), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G101), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n414), .A3(G101), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n415), .A2(KEYINPUT83), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(KEYINPUT83), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n308), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n394), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n406), .A2(new_n419), .A3(new_n407), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n420), .A3(new_n402), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n410), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n420), .ZN(new_n423));
  INV_X1    g237(.A(new_n402), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT6), .A3(new_n421), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n380), .B(KEYINPUT87), .Z(new_n427));
  XNOR2_X1  g241(.A(new_n378), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n429), .A3(new_n424), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n422), .A2(new_n431), .A3(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(KEYINPUT89), .A3(new_n436), .ZN(new_n437));
  OR3_X1    g251(.A1(new_n432), .A2(KEYINPUT89), .A3(new_n434), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(new_n383), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n213), .B(KEYINPUT91), .Z(new_n443));
  OAI21_X1  g257(.A(new_n217), .B1(new_n443), .B2(new_n221), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n320), .A2(new_n187), .A3(G214), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n270), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n320), .A2(new_n187), .A3(G143), .A4(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n251), .B1(new_n446), .B2(new_n447), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT92), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT17), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n223), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n448), .B(G131), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n457), .A2(new_n458), .B1(KEYINPUT17), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n456), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n455), .B1(new_n452), .B2(KEYINPUT17), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n222), .B(new_n214), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT93), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n442), .B(new_n451), .C1(new_n460), .C2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n215), .A2(KEYINPUT19), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n443), .B2(KEYINPUT19), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n214), .B(new_n459), .C1(new_n467), .C2(new_n272), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n451), .ZN(new_n469));
  INV_X1    g283(.A(new_n442), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G475), .A2(G902), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(KEYINPUT20), .B2(new_n474), .ZN(new_n478));
  INV_X1    g292(.A(new_n465), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n459), .A2(KEYINPUT17), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n463), .B2(KEYINPUT93), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n457), .A2(new_n458), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n442), .B1(new_n483), .B2(new_n451), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n229), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G475), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G952), .ZN(new_n489));
  AOI211_X1 g303(.A(G953), .B(new_n489), .C1(G234), .C2(G237), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n229), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT21), .B(G898), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT98), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT94), .B(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G116), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT95), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT95), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n499), .A3(G116), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n299), .A2(G122), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT14), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(KEYINPUT97), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n502), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n498), .A2(new_n500), .B1(KEYINPUT14), .B2(new_n502), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT97), .ZN(new_n510));
  OAI21_X1  g324(.A(G107), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n500), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n499), .B1(new_n496), .B2(G116), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n391), .B(new_n502), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n501), .A2(KEYINPUT96), .A3(new_n391), .A4(new_n502), .ZN(new_n517));
  XNOR2_X1  g331(.A(G128), .B(G143), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n245), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n501), .A2(new_n502), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G107), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n270), .A2(G128), .ZN(new_n524));
  OAI21_X1  g338(.A(G134), .B1(new_n524), .B2(KEYINPUT13), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n518), .B2(KEYINPUT13), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n245), .B2(new_n518), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n511), .A2(new_n520), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT9), .B(G234), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n529), .A2(new_n235), .A3(G953), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n495), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n527), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n509), .A2(KEYINPUT97), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n509), .A2(KEYINPUT97), .B1(new_n506), .B2(new_n505), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n391), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n530), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(KEYINPUT98), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n528), .A2(new_n530), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n229), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n229), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(KEYINPUT99), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT99), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n541), .A2(new_n229), .A3(new_n546), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n541), .B2(new_n229), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n488), .A2(new_n494), .A3(new_n548), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G469), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G140), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n187), .A2(G227), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n192), .B1(new_n281), .B2(KEYINPUT1), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n268), .B1(new_n287), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n390), .A3(new_n393), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n289), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n419), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n294), .A2(new_n295), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n566), .A2(new_n567), .A3(new_n570), .A4(new_n568), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n558), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n274), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n394), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n564), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n571), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n562), .A2(new_n563), .B1(new_n575), .B2(new_n394), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT12), .B1(new_n580), .B2(new_n570), .ZN(new_n581));
  AND4_X1   g395(.A1(new_n573), .A2(new_n579), .A3(new_n558), .A4(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n554), .B(new_n229), .C1(new_n574), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n554), .A2(new_n229), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n573), .A2(new_n581), .A3(new_n579), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n557), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n572), .A2(new_n573), .A3(new_n558), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(G469), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n583), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G221), .B1(new_n529), .B2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n440), .A2(new_n553), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n376), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND2_X1  g409(.A1(new_n366), .A2(new_n229), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n366), .A2(new_n367), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n241), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n435), .A2(KEYINPUT100), .A3(new_n436), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n422), .A2(new_n431), .A3(new_n602), .A4(new_n433), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n603), .A2(new_n439), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n541), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n537), .A2(new_n538), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n540), .A3(KEYINPUT33), .ZN(new_n610));
  AND4_X1   g424(.A1(G478), .A2(new_n608), .A3(new_n229), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(G478), .B1(new_n541), .B2(new_n229), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n494), .B(new_n487), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n552), .A2(new_n548), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n472), .A2(new_n475), .A3(new_n473), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n477), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(new_n486), .A3(new_n494), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n617), .B2(new_n621), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n606), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NAND2_X1  g440(.A1(new_n218), .A2(new_n224), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n234), .A2(new_n236), .B1(new_n238), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n599), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n593), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n601), .A2(new_n604), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n373), .B2(new_n375), .ZN(new_n636));
  INV_X1    g450(.A(new_n592), .ZN(new_n637));
  INV_X1    g451(.A(new_n630), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n475), .B1(new_n472), .B2(new_n473), .ZN(new_n639));
  INV_X1    g453(.A(new_n473), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n476), .B(new_n640), .C1(new_n465), .C2(new_n471), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n490), .ZN(new_n643));
  INV_X1    g457(.A(new_n491), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(G900), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT102), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n451), .B1(new_n460), .B2(new_n464), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n470), .ZN(new_n649));
  AOI21_X1  g463(.A(G902), .B1(new_n649), .B2(new_n465), .ZN(new_n650));
  INV_X1    g464(.A(G475), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n617), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XOR2_X1   g470(.A(new_n646), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n637), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n437), .A2(new_n438), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n229), .B1(new_n312), .B2(new_n352), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n324), .B1(new_n340), .B2(new_n311), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n370), .A2(new_n368), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n617), .A2(new_n487), .ZN(new_n668));
  INV_X1    g482(.A(new_n439), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n638), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n660), .A2(new_n663), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n270), .ZN(G45));
  OAI211_X1 g486(.A(new_n487), .B(new_n647), .C1(new_n611), .C2(new_n612), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT105), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n635), .B(new_n630), .C1(new_n373), .C2(new_n375), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n637), .A4(new_n674), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(new_n229), .B1(new_n574), .B2(new_n582), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n683), .A2(new_n591), .A3(new_n583), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n605), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n613), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n376), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n376), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT41), .B(G113), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT107), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n691), .B(new_n693), .ZN(G15));
  INV_X1    g508(.A(new_n684), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n622), .A2(new_n695), .A3(new_n623), .A4(new_n241), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n636), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  AND4_X1   g512(.A1(KEYINPUT75), .A2(new_n351), .A3(new_n368), .A4(new_n370), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT75), .B1(new_n374), .B2(new_n368), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n605), .B(new_n638), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n701), .A2(new_n553), .A3(new_n695), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NOR4_X1   g517(.A1(new_n695), .A2(new_n668), .A3(new_n635), .A4(new_n493), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n352), .B1(new_n313), .B2(new_n319), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n357), .A2(new_n365), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n367), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n597), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n241), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  INV_X1    g525(.A(new_n685), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n630), .A2(new_n708), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n674), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(new_n591), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n583), .A2(new_n585), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n587), .A2(new_n588), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT108), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT108), .B1(new_n586), .B2(new_n557), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(G469), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n716), .B1(new_n718), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n669), .B1(new_n437), .B2(new_n438), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n376), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(new_n725), .A3(new_n674), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n368), .A2(KEYINPUT109), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n374), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n368), .A2(KEYINPUT109), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n240), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT42), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n251), .ZN(G33));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n376), .A3(new_n654), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  NOR2_X1   g552(.A1(new_n611), .A2(new_n612), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n487), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT43), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n599), .A3(new_n638), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n725), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n587), .B2(new_n588), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n721), .B1(new_n719), .B2(KEYINPUT108), .ZN(new_n748));
  AOI211_X1 g562(.A(new_n554), .B(new_n747), .C1(new_n748), .C2(KEYINPUT45), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(new_n584), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n583), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n716), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n657), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n242), .ZN(G39));
  XNOR2_X1  g572(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n673), .A2(new_n240), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n373), .A3(new_n375), .A4(new_n725), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  AND2_X1   g581(.A1(new_n683), .A2(new_n583), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT49), .Z(new_n769));
  NAND4_X1  g583(.A1(new_n740), .A2(new_n240), .A3(new_n439), .A4(new_n591), .ZN(new_n770));
  OR4_X1    g584(.A1(new_n663), .A2(new_n769), .A3(new_n667), .A4(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n741), .A2(new_n490), .A3(new_n709), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n663), .A2(new_n439), .A3(new_n695), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT50), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n725), .A2(new_n684), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(KEYINPUT121), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(KEYINPUT121), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n643), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n241), .A2(new_n667), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n781), .A2(new_n487), .A3(new_n612), .A4(new_n611), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n741), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n630), .A3(new_n708), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n775), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n768), .A2(new_n716), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n725), .B(new_n772), .C1(new_n762), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT51), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n783), .A2(new_n733), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT48), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n489), .B(G953), .C1(new_n772), .C2(new_n712), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n487), .B1(new_n611), .B2(new_n612), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n792), .B2(new_n781), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT51), .B1(new_n785), .B2(new_n787), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT122), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n594), .A2(new_n632), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n440), .A2(new_n800), .A3(new_n613), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n440), .B2(new_n613), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n545), .A2(new_n547), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n488), .A2(new_n494), .A3(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n801), .B(new_n802), .C1(new_n440), .C2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n799), .B1(new_n600), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n725), .A2(new_n638), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n646), .B1(new_n485), .B2(G475), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n545), .A2(new_n620), .A3(new_n808), .A4(new_n547), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n653), .A2(new_n811), .A3(new_n545), .A4(new_n547), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n810), .A2(new_n812), .A3(new_n591), .A4(new_n590), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n373), .B2(new_n375), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n554), .B(new_n721), .C1(new_n719), .C2(KEYINPUT108), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n591), .B1(new_n815), .B2(new_n717), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n708), .A3(new_n673), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n807), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n818), .A2(new_n819), .A3(new_n737), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n818), .B2(new_n737), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n806), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n735), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n696), .A2(new_n636), .B1(new_n709), .B2(new_n704), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n691), .A2(new_n824), .A3(new_n702), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n655), .A2(new_n714), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n679), .B2(new_n676), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n630), .A2(new_n647), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n816), .A2(new_n830), .A3(KEYINPUT115), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n816), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n668), .A2(new_n635), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n667), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n655), .A2(new_n714), .ZN(new_n836));
  AND4_X1   g650(.A1(KEYINPUT52), .A2(new_n680), .A3(new_n836), .A4(new_n834), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n823), .B(new_n827), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n701), .A2(new_n592), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n678), .B1(new_n841), .B2(new_n674), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n675), .A2(KEYINPUT105), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n836), .B(new_n834), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n822), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n848), .A2(new_n849), .A3(new_n827), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n826), .B(new_n822), .C1(new_n846), .C2(new_n847), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n849), .B1(new_n854), .B2(new_n851), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT118), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(KEYINPUT54), .C1(new_n853), .C2(new_n855), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n823), .B1(new_n835), .B2(new_n837), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n825), .A2(new_n702), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n691), .A4(new_n824), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n826), .A2(KEYINPUT119), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT53), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n839), .B1(new_n827), .B2(new_n862), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n848), .A3(new_n868), .A4(new_n864), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n838), .A2(new_n850), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n866), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n857), .A2(new_n859), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n798), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n771), .B1(new_n874), .B2(new_n875), .ZN(G75));
  NAND3_X1  g690(.A1(new_n866), .A2(new_n869), .A3(new_n870), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G210), .A3(G902), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n428), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n879), .A3(new_n428), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n426), .A2(new_n430), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT123), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT55), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n889), .A3(new_n883), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n187), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(G51));
  NAND2_X1  g707(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n872), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n584), .B(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n574), .B2(new_n582), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n877), .A2(G902), .A3(new_n749), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n891), .B1(new_n898), .B2(new_n899), .ZN(G54));
  NAND4_X1  g714(.A1(new_n877), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n901));
  INV_X1    g715(.A(new_n472), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n891), .ZN(G60));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n608), .A2(new_n610), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n873), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n908), .A2(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n891), .B1(new_n895), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n859), .A2(new_n872), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT117), .B1(new_n838), .B2(new_n850), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n852), .A3(new_n840), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n858), .B1(new_n918), .B2(KEYINPUT54), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n910), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n907), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT124), .A3(new_n913), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n915), .A2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  NAND3_X1  g739(.A1(new_n877), .A2(new_n629), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n877), .A2(new_n925), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n892), .B(new_n926), .C1(new_n927), .C2(new_n239), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT61), .Z(G66));
  INV_X1    g743(.A(new_n492), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n187), .B1(new_n930), .B2(new_n379), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n861), .A2(new_n691), .A3(new_n806), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n187), .ZN(new_n933));
  INV_X1    g747(.A(G898), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n886), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  NAND2_X1  g750(.A1(new_n329), .A2(new_n339), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n467), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(G900), .B(G953), .C1(new_n940), .C2(G227), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(G227), .B2(new_n940), .ZN(new_n942));
  OR4_X1    g756(.A1(new_n635), .A2(new_n756), .A3(new_n668), .A4(new_n733), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(new_n824), .A3(new_n737), .A4(new_n766), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n829), .B1(new_n746), .B2(new_n756), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT127), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(G953), .B1(new_n949), .B2(new_n940), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n671), .B1(new_n951), .B2(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n829), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n488), .A2(new_n803), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n658), .B1(new_n792), .B2(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n957), .A2(new_n376), .A3(new_n725), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n757), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n955), .A2(new_n766), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n939), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n942), .B1(new_n950), .B2(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n960), .B2(new_n932), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n891), .B1(new_n965), .B2(new_n665), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n932), .B(new_n944), .C1(new_n947), .C2(new_n948), .ZN(new_n967));
  INV_X1    g781(.A(new_n964), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n341), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n341), .A2(new_n665), .A3(new_n968), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n918), .B2(new_n971), .ZN(G57));
endmodule


