

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(n718), .B(n717), .ZN(n535) );
  INV_X1 U554 ( .A(n712), .ZN(n719) );
  NOR2_X1 U555 ( .A1(n605), .A2(n604), .ZN(n961) );
  INV_X1 U556 ( .A(KEYINPUT97), .ZN(n530) );
  NOR2_X1 U557 ( .A1(n899), .A2(n534), .ZN(n533) );
  INV_X1 U558 ( .A(KEYINPUT27), .ZN(n705) );
  INV_X1 U559 ( .A(n904), .ZN(n539) );
  NAND2_X1 U560 ( .A1(n522), .A2(KEYINPUT33), .ZN(n538) );
  XNOR2_X1 U561 ( .A(n705), .B(KEYINPUT93), .ZN(n706) );
  AND2_X1 U562 ( .A1(n773), .A2(n538), .ZN(n537) );
  NOR2_X1 U563 ( .A1(n655), .A2(n570), .ZN(n668) );
  NAND2_X1 U564 ( .A1(n543), .A2(n526), .ZN(n525) );
  INV_X1 U565 ( .A(G2105), .ZN(n526) );
  XNOR2_X1 U566 ( .A(KEYINPUT76), .B(KEYINPUT13), .ZN(n602) );
  AND2_X1 U567 ( .A1(n961), .A2(n528), .ZN(n521) );
  NOR2_X1 U568 ( .A1(n768), .A2(n539), .ZN(n522) );
  NOR2_X2 U569 ( .A1(n543), .A2(G2105), .ZN(n551) );
  OR2_X1 U570 ( .A1(n777), .A2(n776), .ZN(n523) );
  AND2_X1 U571 ( .A1(n901), .A2(n821), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n1003), .A2(G137), .ZN(n548) );
  XNOR2_X2 U573 ( .A(n525), .B(KEYINPUT17), .ZN(n1003) );
  NAND2_X1 U574 ( .A1(G160), .A2(G40), .ZN(n779) );
  NAND2_X1 U575 ( .A1(G160), .A2(n527), .ZN(n712) );
  AND2_X1 U576 ( .A1(n780), .A2(G40), .ZN(n527) );
  XNOR2_X2 U577 ( .A(n557), .B(n556), .ZN(G160) );
  INV_X1 U578 ( .A(n899), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n532), .A2(n529), .ZN(n723) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n535), .A2(n521), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n535), .A2(n961), .ZN(n724) );
  NAND2_X1 U583 ( .A1(n535), .A2(n533), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n961), .A2(KEYINPUT97), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n536), .A2(n537), .ZN(n774) );
  NAND2_X1 U586 ( .A1(n766), .A2(n522), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n774), .B(KEYINPUT101), .ZN(n778) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(n552), .Z(n540) );
  INV_X1 U589 ( .A(KEYINPUT96), .ZN(n717) );
  XNOR2_X1 U590 ( .A(n707), .B(n706), .ZN(n710) );
  INV_X1 U591 ( .A(KEYINPUT29), .ZN(n733) );
  NOR2_X1 U592 ( .A1(G164), .A2(G1384), .ZN(n780) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n655) );
  NOR2_X1 U594 ( .A1(n524), .A2(n807), .ZN(n808) );
  XNOR2_X1 U595 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U596 ( .A1(G138), .A2(n1003), .ZN(n542) );
  INV_X1 U597 ( .A(G2104), .ZN(n543) );
  NAND2_X1 U598 ( .A1(G102), .A2(n551), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n547) );
  AND2_X1 U600 ( .A1(G2104), .A2(G2105), .ZN(n999) );
  NAND2_X1 U601 ( .A1(G114), .A2(n999), .ZN(n545) );
  AND2_X1 U602 ( .A1(n543), .A2(G2105), .ZN(n1000) );
  NAND2_X1 U603 ( .A1(G126), .A2(n1000), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U606 ( .A1(n999), .A2(G113), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n550), .B(KEYINPUT67), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G101), .A2(n551), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G125), .A2(n1000), .ZN(n553) );
  AND2_X1 U611 ( .A1(n540), .A2(n553), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U613 ( .A(KEYINPUT66), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n1000), .A2(G123), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT18), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G135), .A2(n1003), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U618 ( .A(KEYINPUT82), .B(n561), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G111), .A2(n999), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G99), .A2(n551), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT83), .B(n566), .ZN(n998) );
  XNOR2_X1 U624 ( .A(G2096), .B(n998), .ZN(n567) );
  OR2_X1 U625 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U626 ( .A(G69), .ZN(G235) );
  INV_X1 U627 ( .A(G651), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G75), .A2(n668), .ZN(n569) );
  NOR2_X1 U629 ( .A1(G651), .A2(G543), .ZN(n669) );
  NAND2_X1 U630 ( .A1(G88), .A2(n669), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n576) );
  NOR2_X1 U632 ( .A1(G543), .A2(n570), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT1), .B(n571), .Z(n672) );
  NAND2_X1 U634 ( .A1(G62), .A2(n672), .ZN(n574) );
  NOR2_X1 U635 ( .A1(G651), .A2(n655), .ZN(n572) );
  XOR2_X2 U636 ( .A(KEYINPUT65), .B(n572), .Z(n673) );
  NAND2_X1 U637 ( .A1(G50), .A2(n673), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(G166) );
  NAND2_X1 U640 ( .A1(n669), .A2(G89), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT4), .B(n577), .Z(n580) );
  NAND2_X1 U642 ( .A1(n668), .A2(G76), .ZN(n578) );
  XOR2_X1 U643 ( .A(n578), .B(KEYINPUT78), .Z(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT79), .B(n581), .Z(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT5), .B(n582), .Z(n589) );
  NAND2_X1 U647 ( .A1(n672), .A2(G63), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT80), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G51), .A2(n673), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT6), .B(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(KEYINPUT81), .B(n587), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(KEYINPUT7), .B(n590), .ZN(G168) );
  NAND2_X1 U655 ( .A1(G94), .A2(G452), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n592), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n828) );
  NAND2_X1 U660 ( .A1(n828), .A2(G567), .ZN(n593) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  NAND2_X1 U662 ( .A1(n672), .A2(G56), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n594), .B(KEYINPUT14), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G43), .A2(n673), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT77), .B(n595), .Z(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n605) );
  NAND2_X1 U667 ( .A1(n668), .A2(G68), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT75), .B(n598), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n669), .A2(G81), .ZN(n599) );
  XOR2_X1 U670 ( .A(n599), .B(KEYINPUT12), .Z(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n961), .A2(G860), .ZN(G153) );
  NAND2_X1 U673 ( .A1(G77), .A2(n668), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G90), .A2(n669), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n608), .B(KEYINPUT9), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G52), .A2(n673), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U679 ( .A1(G64), .A2(n672), .ZN(n611) );
  XNOR2_X1 U680 ( .A(KEYINPUT71), .B(n611), .ZN(n612) );
  NOR2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U682 ( .A(KEYINPUT72), .B(n614), .ZN(G171) );
  INV_X1 U683 ( .A(G171), .ZN(G301) );
  NAND2_X1 U684 ( .A1(G301), .A2(G868), .ZN(n623) );
  NAND2_X1 U685 ( .A1(G79), .A2(n668), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G92), .A2(n669), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G66), .A2(n672), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G54), .A2(n673), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT15), .ZN(n899) );
  INV_X1 U693 ( .A(G868), .ZN(n682) );
  NAND2_X1 U694 ( .A1(n899), .A2(n682), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(G284) );
  XOR2_X1 U696 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U697 ( .A1(G78), .A2(n668), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G91), .A2(n669), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U700 ( .A(KEYINPUT74), .B(n626), .Z(n630) );
  NAND2_X1 U701 ( .A1(G65), .A2(n672), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G53), .A2(n673), .ZN(n627) );
  AND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(G299) );
  NOR2_X1 U705 ( .A1(G286), .A2(n682), .ZN(n632) );
  NOR2_X1 U706 ( .A1(G868), .A2(G299), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(G297) );
  INV_X1 U708 ( .A(G860), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n633), .A2(G559), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n634), .A2(n528), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U712 ( .A1(n528), .A2(G868), .ZN(n636) );
  NOR2_X1 U713 ( .A1(G559), .A2(n636), .ZN(n638) );
  AND2_X1 U714 ( .A1(n682), .A2(n961), .ZN(n637) );
  NOR2_X1 U715 ( .A1(n638), .A2(n637), .ZN(G282) );
  NAND2_X1 U716 ( .A1(G85), .A2(n669), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT68), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G72), .A2(n668), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G60), .A2(n672), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G47), .A2(n673), .ZN(n642) );
  XNOR2_X1 U722 ( .A(KEYINPUT69), .B(n642), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U725 ( .A(KEYINPUT70), .B(n647), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G48), .A2(n673), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G86), .A2(n669), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G73), .A2(n668), .ZN(n650) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n672), .A2(G61), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U734 ( .A1(G87), .A2(n655), .ZN(n657) );
  NAND2_X1 U735 ( .A1(G74), .A2(G651), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U737 ( .A1(n672), .A2(n658), .ZN(n661) );
  NAND2_X1 U738 ( .A1(G49), .A2(n673), .ZN(n659) );
  XOR2_X1 U739 ( .A(KEYINPUT85), .B(n659), .Z(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(G288) );
  NAND2_X1 U741 ( .A1(n528), .A2(G559), .ZN(n962) );
  XOR2_X1 U742 ( .A(KEYINPUT87), .B(n962), .Z(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n663) );
  XNOR2_X1 U744 ( .A(G166), .B(n961), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U746 ( .A(G290), .B(n664), .ZN(n666) );
  INV_X1 U747 ( .A(G299), .ZN(n728) );
  XNOR2_X1 U748 ( .A(G305), .B(n728), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n667), .B(G288), .ZN(n679) );
  NAND2_X1 U751 ( .A1(G80), .A2(n668), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G93), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G67), .A2(n672), .ZN(n675) );
  NAND2_X1 U755 ( .A1(G55), .A2(n673), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U758 ( .A(n678), .B(KEYINPUT84), .Z(n965) );
  XOR2_X1 U759 ( .A(n679), .B(n965), .Z(n1024) );
  XNOR2_X1 U760 ( .A(n680), .B(n1024), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n681), .A2(G868), .ZN(n684) );
  NAND2_X1 U762 ( .A1(n682), .A2(n965), .ZN(n683) );
  NAND2_X1 U763 ( .A1(n684), .A2(n683), .ZN(G295) );
  NAND2_X1 U764 ( .A1(G2084), .A2(G2078), .ZN(n685) );
  XOR2_X1 U765 ( .A(KEYINPUT20), .B(n685), .Z(n686) );
  NAND2_X1 U766 ( .A1(G2090), .A2(n686), .ZN(n687) );
  XNOR2_X1 U767 ( .A(KEYINPUT21), .B(n687), .ZN(n688) );
  NAND2_X1 U768 ( .A1(n688), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n689), .ZN(G158) );
  XNOR2_X1 U770 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U771 ( .A1(G120), .A2(G57), .ZN(n690) );
  NOR2_X1 U772 ( .A1(G235), .A2(n690), .ZN(n691) );
  XNOR2_X1 U773 ( .A(KEYINPUT90), .B(n691), .ZN(n692) );
  NAND2_X1 U774 ( .A1(n692), .A2(G108), .ZN(n966) );
  NAND2_X1 U775 ( .A1(n966), .A2(G567), .ZN(n698) );
  XOR2_X1 U776 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n694) );
  NAND2_X1 U777 ( .A1(G132), .A2(G82), .ZN(n693) );
  XNOR2_X1 U778 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U779 ( .A1(n695), .A2(G218), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G96), .A2(n696), .ZN(n967) );
  NAND2_X1 U781 ( .A1(n967), .A2(G2106), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n698), .A2(n697), .ZN(n1035) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n699) );
  XOR2_X1 U784 ( .A(KEYINPUT91), .B(n699), .Z(n700) );
  NOR2_X1 U785 ( .A1(n1035), .A2(n700), .ZN(n832) );
  NAND2_X1 U786 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U787 ( .A(G166), .ZN(G303) );
  INV_X1 U788 ( .A(G1961), .ZN(n927) );
  NAND2_X1 U789 ( .A1(n712), .A2(n927), .ZN(n704) );
  XNOR2_X1 U790 ( .A(G2078), .B(KEYINPUT25), .ZN(n702) );
  XNOR2_X1 U791 ( .A(n702), .B(KEYINPUT92), .ZN(n883) );
  NAND2_X1 U792 ( .A1(n719), .A2(n883), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n740) );
  NAND2_X1 U794 ( .A1(n740), .A2(G171), .ZN(n736) );
  NAND2_X1 U795 ( .A1(G2072), .A2(n719), .ZN(n707) );
  XOR2_X1 U796 ( .A(G1956), .B(KEYINPUT94), .Z(n932) );
  NOR2_X1 U797 ( .A1(n719), .A2(n932), .ZN(n708) );
  XOR2_X1 U798 ( .A(KEYINPUT95), .B(n708), .Z(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n727) );
  NOR2_X1 U800 ( .A1(n728), .A2(n727), .ZN(n711) );
  XOR2_X1 U801 ( .A(n711), .B(KEYINPUT28), .Z(n732) );
  INV_X1 U802 ( .A(G1996), .ZN(n875) );
  NOR2_X1 U803 ( .A1(n712), .A2(n875), .ZN(n714) );
  XOR2_X1 U804 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n713) );
  XNOR2_X1 U805 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n712), .A2(G1341), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U808 ( .A1(G2067), .A2(n712), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n719), .A2(G1348), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U812 ( .A1(n899), .A2(n724), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n734) );
  XNOR2_X1 U817 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U818 ( .A1(n736), .A2(n735), .ZN(n745) );
  NAND2_X1 U819 ( .A1(G8), .A2(n712), .ZN(n777) );
  NOR2_X1 U820 ( .A1(G1966), .A2(n777), .ZN(n756) );
  NOR2_X1 U821 ( .A1(G2084), .A2(n712), .ZN(n757) );
  NOR2_X1 U822 ( .A1(n756), .A2(n757), .ZN(n737) );
  NAND2_X1 U823 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U824 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U825 ( .A1(G168), .A2(n739), .ZN(n742) );
  NOR2_X1 U826 ( .A1(n740), .A2(G171), .ZN(n741) );
  NOR2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U828 ( .A(KEYINPUT31), .B(n743), .Z(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n754) );
  NAND2_X1 U830 ( .A1(n754), .A2(G286), .ZN(n751) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n777), .ZN(n746) );
  XNOR2_X1 U832 ( .A(KEYINPUT99), .B(n746), .ZN(n749) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n712), .ZN(n747) );
  NOR2_X1 U834 ( .A1(G166), .A2(n747), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U838 ( .A(n753), .B(KEYINPUT32), .ZN(n761) );
  XOR2_X1 U839 ( .A(n754), .B(KEYINPUT98), .Z(n755) );
  NOR2_X1 U840 ( .A1(n756), .A2(n755), .ZN(n759) );
  NAND2_X1 U841 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U842 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U843 ( .A1(n761), .A2(n760), .ZN(n770) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n912) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n918) );
  NOR2_X1 U846 ( .A1(n912), .A2(n918), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n770), .A2(n762), .ZN(n763) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n913) );
  NAND2_X1 U849 ( .A1(n763), .A2(n913), .ZN(n764) );
  XNOR2_X1 U850 ( .A(n764), .B(KEYINPUT100), .ZN(n765) );
  NOR2_X1 U851 ( .A1(n765), .A2(n777), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n912), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U853 ( .A1(n777), .A2(n767), .ZN(n768) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n904) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G8), .A2(n769), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n772), .A2(n777), .ZN(n773) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U860 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  NAND2_X1 U861 ( .A1(n778), .A2(n523), .ZN(n809) );
  XNOR2_X1 U862 ( .A(G1986), .B(G290), .ZN(n901) );
  NOR2_X1 U863 ( .A1(n780), .A2(n779), .ZN(n821) );
  NAND2_X1 U864 ( .A1(G141), .A2(n1003), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G129), .A2(n1000), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n551), .A2(G105), .ZN(n783) );
  XOR2_X1 U868 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U870 ( .A1(n999), .A2(G117), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n1019) );
  AND2_X1 U872 ( .A1(n1019), .A2(G1996), .ZN(n795) );
  NAND2_X1 U873 ( .A1(G131), .A2(n1003), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G95), .A2(n551), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G107), .A2(n999), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G119), .A2(n1000), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n1014) );
  INV_X1 U880 ( .A(G1991), .ZN(n877) );
  NOR2_X1 U881 ( .A1(n1014), .A2(n877), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n855) );
  INV_X1 U883 ( .A(n821), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n855), .A2(n796), .ZN(n813) );
  INV_X1 U885 ( .A(n813), .ZN(n806) );
  NAND2_X1 U886 ( .A1(G140), .A2(n1003), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G104), .A2(n551), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n799), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G116), .A2(n999), .ZN(n801) );
  NAND2_X1 U891 ( .A1(G128), .A2(n1000), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n802), .Z(n803) );
  NOR2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n805), .ZN(n996) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U897 ( .A1(n996), .A2(n819), .ZN(n854) );
  NAND2_X1 U898 ( .A1(n821), .A2(n854), .ZN(n818) );
  NAND2_X1 U899 ( .A1(n806), .A2(n818), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n825) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n1019), .ZN(n861) );
  AND2_X1 U902 ( .A1(n877), .A2(n1014), .ZN(n857) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n810) );
  XNOR2_X1 U904 ( .A(KEYINPUT102), .B(n810), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n857), .A2(n811), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U907 ( .A1(n861), .A2(n814), .ZN(n815) );
  XOR2_X1 U908 ( .A(n815), .B(KEYINPUT39), .Z(n816) );
  XNOR2_X1 U909 ( .A(KEYINPUT103), .B(n816), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n996), .A2(n819), .ZN(n852) );
  NAND2_X1 U912 ( .A1(n820), .A2(n852), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U914 ( .A(KEYINPUT104), .B(n823), .ZN(n824) );
  NAND2_X1 U915 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n826) );
  XNOR2_X1 U917 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U918 ( .A1(n828), .A2(G2106), .ZN(n829) );
  XOR2_X1 U919 ( .A(KEYINPUT107), .B(n829), .Z(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U921 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U924 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  NAND2_X1 U926 ( .A1(G124), .A2(n1000), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT44), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n999), .A2(G112), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n839) );
  NAND2_X1 U930 ( .A1(G136), .A2(n1003), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G100), .A2(n551), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G162) );
  XOR2_X1 U934 ( .A(G164), .B(G2078), .Z(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT116), .B(n840), .ZN(n850) );
  NAND2_X1 U936 ( .A1(G139), .A2(n1003), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G103), .A2(n551), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n848) );
  NAND2_X1 U939 ( .A1(G115), .A2(n999), .ZN(n844) );
  NAND2_X1 U940 ( .A1(G127), .A2(n1000), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(KEYINPUT47), .B(n845), .Z(n846) );
  XNOR2_X1 U943 ( .A(KEYINPUT112), .B(n846), .ZN(n847) );
  NOR2_X1 U944 ( .A1(n848), .A2(n847), .ZN(n1013) );
  XOR2_X1 U945 ( .A(G2072), .B(n1013), .Z(n849) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT50), .B(n851), .Z(n869) );
  INV_X1 U948 ( .A(n852), .ZN(n853) );
  NOR2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U950 ( .A1(n855), .A2(n998), .ZN(n856) );
  NOR2_X1 U951 ( .A1(n857), .A2(n856), .ZN(n858) );
  NAND2_X1 U952 ( .A1(n859), .A2(n858), .ZN(n866) );
  XNOR2_X1 U953 ( .A(G2084), .B(G160), .ZN(n864) );
  XOR2_X1 U954 ( .A(G2090), .B(G162), .Z(n860) );
  NOR2_X1 U955 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U956 ( .A(KEYINPUT51), .B(n862), .Z(n863) );
  NAND2_X1 U957 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U958 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U959 ( .A(KEYINPUT115), .B(n867), .ZN(n868) );
  NOR2_X1 U960 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U961 ( .A(KEYINPUT52), .B(n870), .ZN(n871) );
  XNOR2_X1 U962 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n894) );
  NAND2_X1 U963 ( .A1(n871), .A2(n894), .ZN(n872) );
  NAND2_X1 U964 ( .A1(n872), .A2(G29), .ZN(n959) );
  XNOR2_X1 U965 ( .A(G2090), .B(G35), .ZN(n889) );
  XNOR2_X1 U966 ( .A(G2067), .B(G26), .ZN(n874) );
  XNOR2_X1 U967 ( .A(G33), .B(G2072), .ZN(n873) );
  NOR2_X1 U968 ( .A1(n874), .A2(n873), .ZN(n882) );
  XNOR2_X1 U969 ( .A(G32), .B(n875), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n876), .A2(G28), .ZN(n880) );
  XOR2_X1 U971 ( .A(KEYINPUT118), .B(n877), .Z(n878) );
  XNOR2_X1 U972 ( .A(G25), .B(n878), .ZN(n879) );
  NOR2_X1 U973 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U974 ( .A1(n882), .A2(n881), .ZN(n885) );
  XOR2_X1 U975 ( .A(G27), .B(n883), .Z(n884) );
  NOR2_X1 U976 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U977 ( .A(KEYINPUT53), .B(n886), .Z(n887) );
  XNOR2_X1 U978 ( .A(n887), .B(KEYINPUT119), .ZN(n888) );
  NOR2_X1 U979 ( .A1(n889), .A2(n888), .ZN(n892) );
  XOR2_X1 U980 ( .A(G2084), .B(KEYINPUT54), .Z(n890) );
  XNOR2_X1 U981 ( .A(G34), .B(n890), .ZN(n891) );
  NAND2_X1 U982 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U983 ( .A(n894), .B(n893), .ZN(n896) );
  INV_X1 U984 ( .A(G29), .ZN(n895) );
  NAND2_X1 U985 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U986 ( .A1(G11), .A2(n897), .ZN(n957) );
  XNOR2_X1 U987 ( .A(G16), .B(KEYINPUT56), .ZN(n926) );
  XOR2_X1 U988 ( .A(G1348), .B(KEYINPUT120), .Z(n898) );
  XNOR2_X1 U989 ( .A(n899), .B(n898), .ZN(n903) );
  XNOR2_X1 U990 ( .A(G1956), .B(G299), .ZN(n900) );
  NOR2_X1 U991 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U992 ( .A1(n903), .A2(n902), .ZN(n908) );
  XNOR2_X1 U993 ( .A(G1966), .B(G168), .ZN(n905) );
  NAND2_X1 U994 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U995 ( .A(KEYINPUT57), .B(n906), .Z(n907) );
  NOR2_X1 U996 ( .A1(n908), .A2(n907), .ZN(n924) );
  XNOR2_X1 U997 ( .A(G171), .B(G1961), .ZN(n911) );
  XOR2_X1 U998 ( .A(n961), .B(G1341), .Z(n909) );
  XNOR2_X1 U999 ( .A(KEYINPUT123), .B(n909), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(n911), .A2(n910), .ZN(n922) );
  INV_X1 U1001 ( .A(n912), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1003 ( .A(n915), .B(KEYINPUT121), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(G1971), .A2(G303), .ZN(n916) );
  NAND2_X1 U1005 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1006 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1007 ( .A(KEYINPUT122), .B(n920), .Z(n921) );
  NOR2_X1 U1008 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1009 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1010 ( .A1(n926), .A2(n925), .ZN(n955) );
  INV_X1 U1011 ( .A(G16), .ZN(n953) );
  XNOR2_X1 U1012 ( .A(n927), .B(G5), .ZN(n949) );
  XOR2_X1 U1013 ( .A(G1966), .B(G21), .Z(n940) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G19), .ZN(n928) );
  XNOR2_X1 U1015 ( .A(n928), .B(KEYINPUT124), .ZN(n930) );
  XNOR2_X1 U1016 ( .A(G6), .B(G1981), .ZN(n929) );
  NOR2_X1 U1017 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1018 ( .A(KEYINPUT125), .B(n931), .Z(n934) );
  XNOR2_X1 U1019 ( .A(n932), .B(G20), .ZN(n933) );
  NAND2_X1 U1020 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1021 ( .A(KEYINPUT59), .B(G1348), .Z(n935) );
  XNOR2_X1 U1022 ( .A(G4), .B(n935), .ZN(n936) );
  NOR2_X1 U1023 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1024 ( .A(KEYINPUT60), .B(n938), .ZN(n939) );
  NAND2_X1 U1025 ( .A1(n940), .A2(n939), .ZN(n947) );
  XNOR2_X1 U1026 ( .A(G1971), .B(G22), .ZN(n942) );
  XNOR2_X1 U1027 ( .A(G23), .B(G1976), .ZN(n941) );
  NOR2_X1 U1028 ( .A1(n942), .A2(n941), .ZN(n944) );
  XOR2_X1 U1029 ( .A(G1986), .B(G24), .Z(n943) );
  NAND2_X1 U1030 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1031 ( .A(KEYINPUT58), .B(n945), .ZN(n946) );
  NOR2_X1 U1032 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1033 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1034 ( .A(n950), .B(KEYINPUT61), .ZN(n951) );
  XOR2_X1 U1035 ( .A(KEYINPUT126), .B(n951), .Z(n952) );
  NAND2_X1 U1036 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1037 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1038 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1039 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1040 ( .A(KEYINPUT62), .B(n960), .Z(G311) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  XOR2_X1 U1042 ( .A(n962), .B(n961), .Z(n963) );
  NOR2_X1 U1043 ( .A1(G860), .A2(n963), .ZN(n964) );
  XOR2_X1 U1044 ( .A(n965), .B(n964), .Z(G145) );
  INV_X1 U1045 ( .A(G132), .ZN(G219) );
  INV_X1 U1046 ( .A(G108), .ZN(G238) );
  INV_X1 U1047 ( .A(G96), .ZN(G221) );
  INV_X1 U1048 ( .A(G82), .ZN(G220) );
  INV_X1 U1049 ( .A(G57), .ZN(G237) );
  NOR2_X1 U1050 ( .A1(n967), .A2(n966), .ZN(G325) );
  INV_X1 U1051 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1052 ( .A(G2678), .B(G2067), .Z(n969) );
  XNOR2_X1 U1053 ( .A(G2084), .B(G2078), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1055 ( .A(n970), .B(KEYINPUT109), .Z(n972) );
  XNOR2_X1 U1056 ( .A(G2072), .B(KEYINPUT42), .ZN(n971) );
  XNOR2_X1 U1057 ( .A(n972), .B(n971), .ZN(n976) );
  XOR2_X1 U1058 ( .A(G2100), .B(G2096), .Z(n974) );
  XNOR2_X1 U1059 ( .A(G2090), .B(KEYINPUT43), .ZN(n973) );
  XNOR2_X1 U1060 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1061 ( .A(n976), .B(n975), .Z(G227) );
  XOR2_X1 U1062 ( .A(G1986), .B(G1956), .Z(n978) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G1966), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1065 ( .A(n979), .B(KEYINPUT41), .Z(n981) );
  XNOR2_X1 U1066 ( .A(G1961), .B(G1976), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(n981), .B(n980), .ZN(n985) );
  XOR2_X1 U1068 ( .A(G2474), .B(G1991), .Z(n983) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G1971), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(n983), .B(n982), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(n985), .B(n984), .ZN(G229) );
  XNOR2_X1 U1072 ( .A(G1341), .B(G2454), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(n986), .B(G2430), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(n987), .B(G1348), .ZN(n993) );
  XOR2_X1 U1075 ( .A(G2443), .B(G2427), .Z(n989) );
  XNOR2_X1 U1076 ( .A(G2438), .B(G2446), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n989), .B(n988), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G2451), .B(G2435), .Z(n990) );
  XNOR2_X1 U1079 ( .A(n991), .B(n990), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(n993), .B(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n994), .A2(G14), .ZN(n995) );
  XOR2_X1 U1082 ( .A(KEYINPUT106), .B(n995), .Z(G401) );
  XOR2_X1 U1083 ( .A(G160), .B(n996), .Z(n997) );
  XNOR2_X1 U1084 ( .A(n998), .B(n997), .ZN(n1022) );
  NAND2_X1 U1085 ( .A1(G118), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1086 ( .A1(G130), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(G142), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(n1004), .B(KEYINPUT110), .ZN(n1006) );
  NAND2_X1 U1090 ( .A1(G106), .A2(n551), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(KEYINPUT45), .B(n1007), .Z(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1018) );
  XOR2_X1 U1094 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1011) );
  XNOR2_X1 U1095 ( .A(G164), .B(KEYINPUT111), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(n1012), .B(G162), .Z(n1016) );
  XNOR2_X1 U1098 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NOR2_X1 U1103 ( .A1(G37), .A2(n1023), .ZN(G395) );
  XOR2_X1 U1104 ( .A(KEYINPUT113), .B(n1024), .Z(n1026) );
  XNOR2_X1 U1105 ( .A(n528), .B(G286), .ZN(n1025) );
  XNOR2_X1 U1106 ( .A(n1026), .B(n1025), .ZN(n1027) );
  XNOR2_X1 U1107 ( .A(G301), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1108 ( .A1(G37), .A2(n1028), .ZN(G397) );
  NOR2_X1 U1109 ( .A1(G227), .A2(G229), .ZN(n1030) );
  XNOR2_X1 U1110 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n1029) );
  XNOR2_X1 U1111 ( .A(n1030), .B(n1029), .ZN(n1032) );
  OR2_X1 U1112 ( .A1(n1035), .A2(G401), .ZN(n1031) );
  NOR2_X1 U1113 ( .A1(n1032), .A2(n1031), .ZN(n1034) );
  NOR2_X1 U1114 ( .A1(G395), .A2(G397), .ZN(n1033) );
  NAND2_X1 U1115 ( .A1(n1034), .A2(n1033), .ZN(G225) );
  INV_X1 U1116 ( .A(G225), .ZN(G308) );
  INV_X1 U1117 ( .A(n1035), .ZN(G319) );
endmodule

