//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT66), .B(G77), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G87), .A2(G250), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n212), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT68), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n212), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n229), .B(new_n235), .C1(new_n223), .C2(new_n224), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n226), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT70), .B(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G274), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n259), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n269), .B1(new_n270), .B2(new_n272), .C1(new_n214), .C2(new_n271), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n258), .B(new_n261), .C1(new_n273), .C2(new_n259), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n277), .A2(new_n232), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n233), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  INV_X1    g0081(.A(G1), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G13), .A3(G20), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT8), .B(G58), .Z(new_n284));
  NAND2_X1  g0084(.A1(new_n233), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n233), .A2(new_n262), .A3(KEYINPUT71), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT71), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G20), .B2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n284), .A2(new_n286), .B1(new_n290), .B2(G150), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n201), .A2(new_n203), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n281), .B1(G50), .B2(new_n283), .C1(new_n294), .C2(new_n278), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n274), .B2(G169), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n276), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT72), .B1(new_n274), .B2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n274), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n295), .B(KEYINPUT9), .Z(new_n301));
  OR3_X1    g0101(.A1(new_n300), .A2(KEYINPUT10), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n300), .B2(new_n301), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT16), .ZN(new_n305));
  INV_X1    g0105(.A(G68), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT75), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT75), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(new_n264), .A3(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n309), .A3(new_n263), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n311), .B1(new_n271), .B2(G20), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n306), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(G58), .B(G68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G20), .ZN(new_n317));
  INV_X1    g0117(.A(new_n290), .ZN(new_n318));
  INV_X1    g0118(.A(G159), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n305), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n278), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n263), .A2(new_n265), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT7), .B1(new_n323), .B2(new_n233), .ZN(new_n324));
  AOI211_X1 g0124(.A(new_n311), .B(G20), .C1(new_n263), .C2(new_n265), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n290), .A2(G159), .B1(new_n316), .B2(G20), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(KEYINPUT16), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n321), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n279), .A2(new_n284), .ZN(new_n330));
  INV_X1    g0130(.A(new_n284), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n283), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n263), .A2(new_n265), .A3(G226), .A4(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G87), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n335), .B(new_n336), .C1(new_n267), .C2(new_n270), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n259), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n259), .A2(new_n257), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n258), .B1(new_n339), .B2(G232), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G169), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(G179), .A3(new_n340), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT18), .B1(new_n334), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT76), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n323), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n306), .B1(new_n314), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n320), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n278), .B1(new_n351), .B2(KEYINPUT16), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n321), .B1(new_n330), .B2(new_n332), .ZN(new_n353));
  INV_X1    g0153(.A(new_n344), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT76), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n344), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n341), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n299), .B1(new_n338), .B2(new_n340), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n333), .A3(new_n329), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT17), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n353), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n347), .A2(new_n358), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G50), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n318), .A2(new_n370), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n285), .A2(new_n202), .B1(new_n233), .B2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n322), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT73), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n322), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT11), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(KEYINPUT11), .A3(new_n376), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n283), .A2(G68), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT74), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(KEYINPUT74), .A3(new_n382), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n385), .A2(new_n386), .B1(G68), .B2(new_n280), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n379), .A2(new_n380), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n263), .A2(new_n265), .A3(G232), .A4(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n267), .C2(new_n260), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n259), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n258), .B1(new_n339), .B2(G238), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(G179), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G169), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n395), .B2(new_n397), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n397), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n401), .B(G169), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n388), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n259), .A2(new_n257), .A3(new_n215), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n268), .A2(G232), .ZN(new_n409));
  INV_X1    g0209(.A(G238), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n409), .B1(new_n207), .B2(new_n271), .C1(new_n410), .C2(new_n272), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n258), .B(new_n408), .C1(new_n411), .C2(new_n259), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n412), .A2(new_n275), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT15), .B(G87), .Z(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n286), .B1(new_n213), .B2(G20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n284), .A2(new_n290), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n278), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n279), .A2(new_n202), .B1(new_n213), .B2(new_n283), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n412), .B2(G169), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n380), .A2(new_n387), .ZN(new_n424));
  OAI21_X1  g0224(.A(G200), .B1(new_n403), .B2(new_n404), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n395), .A2(G190), .A3(new_n397), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n424), .A2(new_n379), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n420), .B1(new_n412), .B2(G190), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n299), .B2(new_n412), .ZN(new_n429));
  AND4_X1   g0229(.A1(new_n407), .A2(new_n423), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n304), .A2(new_n369), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n207), .B1(new_n313), .B2(new_n314), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n290), .A2(G77), .ZN(new_n434));
  AND2_X1   g0234(.A1(G97), .A2(G107), .ZN(new_n435));
  NOR2_X1   g0235(.A1(G97), .A2(G107), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n435), .A2(new_n436), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G97), .A2(G107), .ZN(new_n438));
  NOR2_X1   g0238(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n208), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n434), .B1(new_n442), .B2(new_n233), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n322), .B1(new_n433), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n283), .A2(G97), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT78), .B1(new_n262), .B2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n282), .A3(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n278), .A2(new_n283), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n445), .B1(new_n450), .B2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT80), .B1(new_n453), .B2(KEYINPUT79), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT80), .ZN(new_n456));
  OAI21_X1  g0256(.A(G244), .B1(new_n456), .B2(KEYINPUT4), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n267), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n215), .B1(KEYINPUT80), .B2(new_n453), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n271), .A2(new_n459), .A3(new_n266), .A4(new_n454), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n259), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n256), .A2(G1), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n232), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(G257), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G274), .A3(new_n465), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n452), .B1(G200), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n464), .B2(new_n478), .ZN(new_n482));
  AOI211_X1 g0282(.A(KEYINPUT81), .B(new_n477), .C1(new_n463), .C2(new_n259), .ZN(new_n483));
  OAI21_X1  g0283(.A(G190), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n482), .A2(new_n483), .A3(G169), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n477), .B1(new_n463), .B2(new_n259), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n275), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n452), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n481), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n399), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n452), .A2(new_n489), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT82), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n485), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(new_n266), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n263), .A2(new_n265), .A3(G264), .A4(G1698), .ZN(new_n499));
  INV_X1    g0299(.A(G303), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n271), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n259), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n282), .A2(G45), .A3(G274), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n473), .B2(new_n474), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n475), .A2(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G270), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n448), .A2(new_n283), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(G116), .A3(new_n278), .A4(new_n446), .ZN(new_n509));
  INV_X1    g0309(.A(new_n283), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n277), .A2(new_n232), .B1(G20), .B2(new_n511), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n461), .B(new_n233), .C1(G33), .C2(new_n206), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n509), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n507), .A2(G169), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n502), .A2(new_n506), .A3(G190), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n468), .A2(G270), .A3(new_n471), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n476), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n259), .B2(new_n501), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n521), .B(new_n522), .C1(new_n525), .C2(new_n299), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT21), .A4(G169), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(G179), .A3(new_n517), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n520), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n233), .B1(new_n390), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n436), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n263), .A2(new_n265), .A3(new_n233), .A4(G68), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n530), .B1(new_n285), .B2(new_n206), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n322), .ZN(new_n538));
  INV_X1    g0338(.A(new_n414), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n510), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n446), .A2(new_n448), .A3(new_n283), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G87), .A3(new_n278), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n263), .A2(new_n265), .A3(G238), .A4(new_n266), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n259), .ZN(new_n549));
  OAI21_X1  g0349(.A(G250), .B1(new_n256), .B2(G1), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n503), .B1(new_n259), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n548), .B2(new_n259), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n544), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n399), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n449), .B2(new_n539), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n541), .A2(KEYINPUT83), .A3(new_n278), .A4(new_n414), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n560), .A2(new_n538), .A3(new_n540), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n275), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n529), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n450), .A2(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n283), .A2(G107), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n271), .A2(new_n233), .A3(G87), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n233), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n286), .A2(G116), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n323), .A2(G20), .A3(new_n532), .ZN(new_n578));
  XOR2_X1   g0378(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n579));
  OAI211_X1 g0379(.A(new_n573), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n278), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n570), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n468), .A2(G264), .A3(new_n471), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n263), .A2(new_n265), .A3(G250), .A4(new_n266), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT85), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n271), .A2(new_n589), .A3(G250), .A4(new_n266), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n586), .B1(new_n593), .B2(new_n259), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n399), .B1(new_n594), .B2(new_n476), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n476), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(new_n275), .ZN(new_n598));
  AOI211_X1 g0398(.A(KEYINPUT86), .B(new_n399), .C1(new_n594), .C2(new_n476), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n585), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(G200), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n594), .A2(G190), .A3(new_n476), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n584), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n566), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n432), .A2(new_n497), .A3(new_n604), .ZN(G372));
  AND2_X1   g0405(.A1(new_n422), .A2(new_n427), .ZN(new_n606));
  INV_X1    g0406(.A(new_n407), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n367), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n355), .A2(new_n357), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n610), .A2(KEYINPUT90), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n302), .A2(new_n303), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(KEYINPUT90), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n297), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n487), .B1(new_n486), .B2(new_n490), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT82), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(new_n617), .B1(new_n484), .B2(new_n480), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n520), .A2(new_n527), .A3(new_n528), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT89), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n520), .A2(new_n621), .A3(new_n527), .A4(new_n528), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n600), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n603), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n543), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n538), .A2(KEYINPUT87), .A3(new_n540), .A4(new_n542), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n627), .A2(new_n554), .A3(new_n556), .A4(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n629), .B2(new_n564), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n564), .A3(new_n625), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n618), .A2(new_n623), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n564), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n494), .A2(new_n495), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n631), .B2(new_n632), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n616), .A2(new_n617), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n640), .B2(new_n565), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n634), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n431), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n615), .A2(new_n643), .ZN(G369));
  INV_X1    g0444(.A(KEYINPUT91), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n233), .A2(G13), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n282), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n529), .A2(new_n645), .B1(new_n517), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n645), .B2(new_n529), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n620), .A2(new_n622), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n517), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n600), .A2(new_n603), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n585), .A2(new_n652), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n600), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n652), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n652), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n619), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT92), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n652), .B(KEYINPUT93), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n665), .A2(new_n670), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n227), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n533), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n230), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n482), .A2(new_n483), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n490), .B1(new_n682), .B2(new_n399), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n629), .A2(new_n564), .A3(new_n625), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n630), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT26), .ZN(new_n686));
  INV_X1    g0486(.A(new_n565), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n616), .A2(new_n617), .A3(new_n638), .A4(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n686), .A2(new_n564), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n618), .B(new_n633), .C1(new_n663), .C2(new_n619), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n652), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n594), .A2(new_n525), .A3(G179), .A4(new_n555), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n682), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n555), .A2(new_n502), .A3(new_n506), .A4(G179), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n593), .A2(new_n259), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n697), .A2(new_n698), .A3(new_n586), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n699), .B(KEYINPUT30), .C1(new_n482), .C2(new_n483), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n525), .A2(G179), .A3(new_n555), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n479), .A3(new_n597), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT94), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n696), .A2(new_n700), .A3(KEYINPUT94), .A4(new_n702), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n652), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n618), .A2(new_n660), .A3(new_n566), .A4(new_n672), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n642), .A2(new_n692), .A3(new_n672), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n693), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n681), .B1(new_n716), .B2(G1), .ZN(G364));
  AOI21_X1  g0517(.A(new_n282), .B1(new_n646), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n676), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n659), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n657), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n271), .A2(new_n227), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n210), .A2(new_n725), .B1(G116), .B2(new_n227), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n250), .A2(G45), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n675), .A2(new_n271), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n256), .B2(new_n231), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n232), .B1(G20), .B2(new_n399), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n720), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n233), .B1(new_n739), .B2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(G58), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n233), .A2(new_n359), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n275), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n271), .B1(new_n740), .B2(new_n206), .C1(new_n741), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n275), .A2(new_n299), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n233), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n743), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G50), .A2(new_n748), .B1(new_n751), .B2(new_n213), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n746), .A2(new_n749), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n306), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n299), .A2(G179), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT97), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n742), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n745), .B(new_n754), .C1(G87), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n749), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G107), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n749), .A2(new_n739), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n759), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  INV_X1    g0570(.A(G329), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n744), .A2(new_n770), .B1(new_n764), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n323), .B1(new_n740), .B2(new_n773), .C1(new_n747), .C2(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n772), .B(new_n775), .C1(G311), .C2(new_n751), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n753), .B1(new_n778), .B2(G317), .ZN(new_n779));
  INV_X1    g0579(.A(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n758), .A2(G303), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n776), .B(new_n782), .C1(new_n783), .C2(new_n761), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n738), .B1(new_n785), .B2(new_n735), .ZN(new_n786));
  INV_X1    g0586(.A(new_n734), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n657), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n722), .A2(new_n723), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n724), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  INV_X1    g0591(.A(new_n735), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n762), .A2(G87), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n323), .B1(new_n740), .B2(new_n206), .C1(new_n747), .C2(new_n500), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n750), .A2(new_n511), .B1(new_n764), .B2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n783), .A2(new_n753), .B1(new_n744), .B2(new_n773), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n793), .B(new_n798), .C1(new_n207), .C2(new_n757), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n762), .A2(G68), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n750), .A2(new_n319), .ZN(new_n801));
  INV_X1    g0601(.A(G143), .ZN(new_n802));
  INV_X1    g0602(.A(G150), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n744), .B1(new_n753), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(G137), .C2(new_n748), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n271), .B1(new_n740), .B2(new_n741), .C1(new_n808), .C2(new_n764), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n758), .B2(G50), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n800), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n792), .B1(new_n799), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n792), .A2(new_n733), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n720), .B1(new_n813), .B2(G77), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n413), .A2(new_n421), .A3(new_n652), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n420), .A2(new_n652), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n429), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n817), .B2(new_n423), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n812), .B(new_n814), .C1(new_n819), .C2(new_n732), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT100), .Z(new_n821));
  NAND2_X1  g0621(.A1(new_n642), .A2(new_n672), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n819), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n642), .A2(new_n672), .A3(new_n818), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n822), .A2(KEYINPUT101), .A3(new_n819), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n713), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(KEYINPUT102), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n720), .B(new_n829), .C1(new_n713), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(KEYINPUT102), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n821), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G384));
  INV_X1    g0634(.A(KEYINPUT35), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n442), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n442), .A2(new_n835), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(G116), .A3(new_n234), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT36), .Z(new_n839));
  OAI211_X1 g0639(.A(new_n213), .B(new_n231), .C1(new_n741), .C2(new_n306), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n201), .A2(G68), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n282), .B(G13), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n388), .A2(new_n652), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n427), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n407), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(KEYINPUT103), .B(new_n388), .C1(new_n402), .C2(new_n406), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n407), .A2(new_n667), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n818), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n667), .B1(new_n703), .B2(new_n704), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n709), .A2(new_n854), .A3(new_n710), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n305), .B1(new_n350), .B2(new_n320), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(KEYINPUT104), .A3(new_n322), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n328), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT104), .B1(new_n856), .B2(new_n322), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n333), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT105), .ZN(new_n861));
  INV_X1    g0661(.A(new_n650), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n333), .C1(new_n858), .C2(new_n859), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n368), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n354), .A2(new_n650), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n353), .B2(new_n362), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n650), .B1(new_n329), .B2(new_n333), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n334), .A2(new_n344), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n363), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n869), .A2(new_n871), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n867), .B2(new_n876), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n852), .B(new_n855), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT31), .B1(new_n853), .B2(new_n706), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n497), .A2(new_n604), .A3(new_n671), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n851), .B1(new_n885), .B2(new_n854), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT106), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n872), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n875), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n873), .B1(new_n367), .B2(new_n609), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n881), .B1(new_n877), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n886), .A2(KEYINPUT107), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT107), .B1(new_n886), .B2(new_n893), .ZN(new_n895));
  OAI211_X1 g0695(.A(G330), .B(new_n882), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n855), .A2(G330), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n431), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n609), .A2(KEYINPUT76), .B1(new_n364), .B2(new_n366), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n865), .B1(new_n901), .B2(new_n358), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n869), .A2(new_n871), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n875), .A2(new_n870), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n887), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n877), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT40), .B1(new_n886), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n877), .A2(new_n892), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n909), .A2(KEYINPUT40), .A3(new_n852), .A4(new_n855), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT107), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n886), .A2(KEYINPUT107), .A3(new_n893), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n431), .A3(new_n855), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n900), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n693), .A2(new_n714), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n431), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n615), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n916), .B(new_n919), .Z(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT39), .B1(new_n878), .B2(new_n879), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n877), .A2(new_n922), .A3(new_n892), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n847), .A2(new_n667), .A3(new_n848), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n849), .A2(new_n850), .ZN(new_n927));
  INV_X1    g0727(.A(new_n815), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n825), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n907), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n355), .A2(new_n357), .A3(new_n650), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n282), .B2(new_n646), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n920), .A2(new_n932), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n843), .B1(new_n934), .B2(new_n935), .ZN(G367));
  INV_X1    g0736(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n627), .A2(new_n628), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n652), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n684), .B2(new_n630), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n635), .A2(new_n938), .A3(new_n652), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n671), .A2(new_n452), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n618), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n683), .A2(new_n671), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(KEYINPUT109), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT109), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n949), .B2(new_n950), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n952), .A2(new_n600), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n671), .B1(new_n956), .B2(new_n640), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n951), .A2(new_n665), .A3(new_n670), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT42), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n937), .B(new_n947), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n959), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n952), .A2(new_n954), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n663), .B1(new_n616), .B2(new_n617), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n962), .B1(new_n964), .B2(new_n671), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n937), .B1(new_n965), .B2(new_n947), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n957), .A2(new_n959), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT110), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n946), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT110), .B1(new_n965), .B2(new_n945), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n963), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n967), .A2(new_n972), .B1(new_n666), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n947), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT111), .B1(new_n968), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n960), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n973), .A2(new_n666), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n977), .A2(new_n978), .A3(new_n970), .A4(new_n971), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n673), .B2(new_n951), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n660), .A2(new_n661), .B1(new_n663), .B2(new_n652), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n982), .A2(new_n669), .B1(new_n600), .B2(new_n671), .ZN(new_n983));
  INV_X1    g0783(.A(new_n951), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n983), .B2(new_n984), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n986), .A2(new_n666), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n666), .B1(new_n986), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n665), .A2(new_n670), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n982), .A2(new_n669), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT112), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT112), .B1(new_n994), .B2(new_n995), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n658), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n658), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n715), .B1(new_n993), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n676), .B(KEYINPUT41), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n718), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n974), .A2(new_n979), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n753), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n201), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1008), .A2(G159), .B1(new_n751), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1011), .A2(KEYINPUT114), .B1(new_n758), .B2(G58), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n760), .A2(new_n214), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n323), .B(new_n1013), .C1(G137), .C2(new_n765), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(KEYINPUT114), .C2(new_n1011), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n747), .A2(new_n802), .B1(new_n744), .B2(new_n803), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n740), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(G68), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n757), .A2(new_n511), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT46), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n323), .B1(new_n740), .B2(new_n207), .C1(new_n783), .C2(new_n750), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n773), .A2(new_n753), .B1(new_n744), .B2(new_n500), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n747), .A2(new_n795), .B1(new_n764), .B2(new_n780), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n206), .B2(new_n760), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1015), .A2(new_n1019), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT47), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n735), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n245), .A2(new_n729), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n736), .B1(new_n227), .B2(new_n539), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n720), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT115), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n942), .B2(new_n787), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1007), .A2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n720), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n725), .A2(new_n678), .B1(G107), .B2(new_n227), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT116), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n242), .A2(new_n256), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n331), .B2(G50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n678), .A3(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n331), .A2(new_n1042), .A3(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n728), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1038), .B1(new_n1048), .B2(new_n736), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n748), .A2(G322), .B1(new_n751), .B2(G303), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n795), .B2(new_n753), .C1(new_n780), .C2(new_n744), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT48), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n783), .B2(new_n740), .C1(new_n773), .C2(new_n757), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n323), .B1(new_n774), .B2(new_n764), .C1(new_n760), .C2(new_n511), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n762), .A2(G97), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n757), .A2(new_n214), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n271), .B1(new_n747), .B2(new_n319), .C1(new_n539), .C2(new_n740), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n750), .A2(new_n306), .B1(new_n764), .B2(new_n803), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n331), .A2(new_n753), .B1(new_n370), .B2(new_n744), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1055), .A2(new_n1057), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1049), .B1(new_n665), .B2(new_n787), .C1(new_n1064), .C2(new_n792), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n676), .B1(new_n1002), .B2(new_n715), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1003), .A2(new_n716), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1065), .B1(new_n718), .B2(new_n1002), .C1(new_n1066), .C2(new_n1067), .ZN(G393));
  NOR2_X1   g0868(.A1(new_n1002), .A2(new_n715), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n677), .B1(new_n993), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n993), .B2(new_n1069), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n993), .A2(new_n719), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n253), .A2(new_n729), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n737), .B1(G97), .B2(new_n675), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1038), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1008), .A2(G303), .B1(new_n765), .B2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n323), .C1(new_n773), .C2(new_n750), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT52), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n747), .A2(new_n780), .B1(new_n744), .B2(new_n795), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n758), .A2(G283), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1078), .B(new_n1082), .C1(G116), .C2(new_n1017), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT51), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n747), .A2(new_n803), .B1(new_n744), .B2(new_n319), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n758), .A2(G68), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n740), .A2(new_n202), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n271), .B1(new_n764), .B2(new_n802), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n331), .A2(new_n750), .B1(new_n201), .B2(new_n753), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1083), .A2(new_n763), .B1(new_n793), .B2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1076), .B1(new_n792), .B2(new_n1092), .C1(new_n963), .C2(new_n787), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1071), .A2(new_n1072), .A3(new_n1093), .ZN(G390));
  OAI21_X1  g0894(.A(new_n927), .B1(new_n713), .B2(new_n819), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT119), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n897), .A2(new_n851), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT119), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n927), .C1(new_n713), .C2(new_n819), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n825), .A2(new_n928), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n927), .B1(new_n897), .B2(new_n819), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n817), .A2(new_n423), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n815), .B1(new_n691), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n852), .A2(new_n712), .A3(G330), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n615), .A2(new_n918), .A3(new_n899), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n925), .B1(new_n877), .B2(new_n892), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1106), .B2(new_n927), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n927), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n925), .B1(new_n1102), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1107), .C1(new_n1116), .C2(new_n924), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT118), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n921), .B(new_n923), .C1(new_n929), .C2(new_n925), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1097), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT118), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1122), .A3(new_n1114), .A4(new_n1107), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1112), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1108), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n1110), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1118), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1130), .A3(new_n676), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n921), .A2(new_n732), .A3(new_n923), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n720), .B1(new_n813), .B2(new_n284), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n744), .A2(new_n511), .B1(new_n764), .B2(new_n773), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n323), .B1(new_n747), .B2(new_n783), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1088), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n753), .A2(new_n207), .B1(new_n750), .B2(new_n206), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT120), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n757), .A2(new_n532), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1138), .B2(new_n1137), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n800), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT121), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n757), .A2(new_n803), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n271), .B1(new_n740), .B2(new_n319), .C1(new_n747), .C2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n750), .A2(new_n1147), .B1(new_n764), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(G137), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n808), .A2(new_n744), .B1(new_n753), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1146), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1144), .B(new_n1152), .C1(new_n201), .C2(new_n760), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1141), .A2(KEYINPUT121), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1142), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1133), .B1(new_n1155), .B2(new_n735), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1129), .A2(new_n719), .B1(new_n1132), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1131), .A2(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(new_n932), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n295), .A2(new_n862), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n302), .A2(new_n303), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n297), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n304), .A2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n896), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n914), .B2(G330), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1159), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n896), .A2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n912), .A2(new_n913), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1176), .A2(new_n1170), .A3(G330), .A4(new_n882), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n932), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1111), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT123), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT123), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1183), .A4(KEYINPUT57), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1110), .B1(new_n1129), .B2(new_n1109), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1175), .A2(new_n932), .A3(new_n1177), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n932), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1185), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1182), .A2(new_n676), .A3(new_n1184), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1171), .A2(new_n732), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n720), .B1(new_n813), .B2(new_n1009), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n744), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G97), .A2(new_n1008), .B1(new_n1194), .B2(G107), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n783), .B2(new_n764), .C1(new_n539), .C2(new_n750), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n271), .A2(G41), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n306), .B2(new_n740), .C1(new_n511), .C2(new_n747), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n760), .A2(new_n741), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1196), .A2(new_n1059), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT122), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT58), .Z(new_n1202));
  NOR2_X1   g1002(.A1(G33), .A2(G41), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1197), .A2(G50), .A3(new_n1203), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n744), .A2(new_n1145), .B1(new_n750), .B2(new_n1150), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n747), .A2(new_n1148), .B1(new_n753), .B2(new_n808), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G150), .C2(new_n1017), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n757), .B2(new_n1147), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n765), .A2(G124), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1203), .B(new_n1210), .C1(new_n760), .C2(new_n319), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1208), .B2(KEYINPUT59), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1202), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1193), .B1(new_n1214), .B2(new_n735), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1179), .A2(new_n719), .B1(new_n1192), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1191), .A2(new_n1216), .ZN(G375));
  NOR2_X1   g1017(.A1(new_n1128), .A2(new_n1005), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1127), .A2(new_n1110), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n720), .B1(new_n813), .B2(G68), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT124), .Z(new_n1222));
  OAI221_X1 g1022(.A(new_n323), .B1(new_n764), .B2(new_n500), .C1(new_n539), .C2(new_n740), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G283), .A2(new_n1194), .B1(new_n751), .B2(G107), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n511), .B2(new_n753), .C1(new_n773), .C2(new_n747), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G97), .C2(new_n758), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n762), .A2(G77), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n271), .B1(new_n753), .B2(new_n1147), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n747), .A2(new_n808), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1229), .A2(new_n1230), .B1(new_n370), .B2(new_n740), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1228), .B(new_n1231), .C1(new_n1230), .C2(new_n1229), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G137), .A2(new_n1194), .B1(new_n765), .B2(G128), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n803), .B2(new_n750), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1199), .B(new_n1234), .C1(G159), .C2(new_n758), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1226), .A2(new_n1227), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1222), .B1(new_n1236), .B2(new_n792), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n927), .B2(new_n732), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1109), .B2(new_n719), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1220), .A2(new_n1239), .ZN(G381));
  NOR2_X1   g1040(.A1(G375), .A2(G378), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G396), .A2(G384), .A3(G393), .A4(G390), .ZN(new_n1243));
  OR4_X1    g1043(.A1(G387), .A2(new_n1242), .A3(G381), .A4(new_n1243), .ZN(G407));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G343), .C2(new_n1242), .ZN(G409));
  NAND3_X1  g1045(.A1(new_n1007), .A2(new_n1036), .A3(G390), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT127), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(G393), .B(G396), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1246), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n1249), .A3(KEYINPUT127), .A4(new_n1246), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n651), .A2(G213), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1216), .A2(new_n1131), .A3(new_n1157), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1186), .A2(new_n1189), .A3(new_n1005), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G375), .B2(G378), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1219), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1127), .A2(KEYINPUT60), .A3(new_n1110), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n676), .A3(new_n1112), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1239), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n833), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G384), .A2(new_n1239), .A3(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT126), .B1(new_n1261), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1191), .B2(new_n1216), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1260), .A4(new_n1269), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1271), .A2(new_n1275), .A3(KEYINPUT62), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1267), .A2(new_n1268), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1277), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1269), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1278), .B(new_n1280), .C1(new_n1273), .C2(new_n1260), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1273), .A2(new_n1260), .A3(new_n1269), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1281), .B(new_n1282), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1256), .B1(new_n1276), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1281), .A2(new_n1288), .A3(new_n1282), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1287), .B(new_n1289), .C1(new_n1290), .C2(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(new_n1291), .ZN(G405));
  OAI21_X1  g1092(.A(new_n1256), .B1(new_n1241), .B2(new_n1273), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1241), .A2(new_n1273), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1288), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1293), .A2(new_n1269), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1269), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


