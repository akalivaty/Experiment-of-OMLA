//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n205), .A2(new_n204), .B1(new_n215), .B2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n203), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT25), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n206), .A2(new_n207), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(new_n206), .B2(new_n207), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT25), .B(new_n210), .C1(new_n212), .C2(new_n209), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n202), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n213), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n216), .A2(new_n221), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(KEYINPUT25), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n206), .A2(new_n203), .A3(new_n207), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n230), .A2(new_n208), .A3(new_n213), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n229), .B(KEYINPUT66), .C1(new_n231), .C2(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234));
  INV_X1    g033(.A(G113gat), .ZN(new_n235));
  INV_X1    g034(.A(G120gat), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT1), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT71), .B(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n237), .B1(new_n235), .B2(new_n236), .ZN(new_n242));
  INV_X1    g041(.A(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n205), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n249), .A2(KEYINPUT26), .A3(new_n209), .ZN(new_n250));
  AOI211_X1 g049(.A(new_n246), .B(new_n250), .C1(KEYINPUT26), .C2(new_n209), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n252));
  INV_X1    g051(.A(G183gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT27), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT27), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G183gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n255), .B2(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n252), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n254), .A2(new_n256), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT69), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n254), .A2(new_n256), .A3(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n252), .A2(G190gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n267), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n251), .B1(new_n263), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n233), .A2(new_n245), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n245), .B1(new_n233), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT34), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n277), .A2(KEYINPUT34), .A3(new_n278), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT72), .B1(new_n277), .B2(new_n278), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n233), .A2(new_n274), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n238), .A2(new_n240), .B1(new_n243), .B2(new_n242), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n233), .A2(new_n245), .A3(new_n274), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n278), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT32), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n285), .B2(new_n291), .ZN(new_n294));
  XOR2_X1   g093(.A(G15gat), .B(G43gat), .Z(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n288), .A2(new_n278), .A3(new_n289), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n303), .B2(new_n290), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT33), .B1(new_n303), .B2(new_n290), .ZN(new_n305));
  INV_X1    g104(.A(new_n297), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n298), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n299), .B1(new_n298), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n284), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n298), .A2(new_n283), .A3(new_n307), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT36), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n283), .B1(new_n298), .B2(new_n307), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n319));
  AOI221_X4 g118(.A(new_n300), .B1(KEYINPUT33), .B2(new_n297), .C1(new_n303), .C2(new_n290), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n284), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n307), .A3(new_n283), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT74), .A3(new_n312), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(new_n318), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G211gat), .ZN(new_n326));
  INV_X1    g125(.A(G218gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G197gat), .ZN(new_n329));
  INV_X1    g128(.A(G204gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332));
  OAI22_X1  g131(.A1(KEYINPUT22), .A2(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G148gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n339), .A2(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G141gat), .B(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G141gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n336), .B1(new_n342), .B2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G155gat), .B(G162gat), .Z(new_n350));
  AOI22_X1  g149(.A1(new_n344), .A2(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n335), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n354), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n352), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n346), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n350), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G22gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT31), .B(G50gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT81), .B1(new_n363), .B2(new_n364), .ZN(new_n373));
  INV_X1    g172(.A(new_n371), .ZN(new_n374));
  OAI21_X1  g173(.A(G22gat), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n365), .A2(new_n366), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n372), .B2(new_n375), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n335), .ZN(new_n381));
  INV_X1    g180(.A(G226gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n229), .B1(new_n231), .B2(KEYINPUT25), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n274), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n233), .A2(new_n274), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n384), .A2(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n381), .B(new_n386), .C1(new_n387), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n274), .A2(new_n385), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n387), .A2(new_n384), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n392), .B2(new_n381), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT84), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n391), .A2(new_n388), .ZN(new_n402));
  INV_X1    g201(.A(new_n384), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n381), .C1(new_n403), .C2(new_n286), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n401), .A2(new_n404), .B1(new_n405), .B2(new_n335), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n381), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n390), .B(new_n400), .C1(new_n392), .C2(new_n381), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT38), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n397), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n399), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n287), .A2(new_n351), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT4), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n287), .A2(new_n351), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(new_n353), .A3(new_n245), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n420), .A2(KEYINPUT5), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n245), .A2(new_n360), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n413), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT77), .A3(new_n416), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n432), .A3(KEYINPUT4), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n419), .A2(new_n433), .A3(new_n421), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n425), .B(new_n429), .C1(new_n431), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n430), .A2(new_n419), .A3(new_n433), .A4(new_n421), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n425), .B1(new_n437), .B2(new_n429), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n424), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(G57gat), .B(G85gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT80), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n439), .A2(new_n449), .A3(new_n444), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n443), .B(new_n424), .C1(new_n436), .C2(new_n438), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n445), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n439), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT83), .B(new_n424), .C1(new_n436), .C2(new_n438), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n412), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n393), .A2(KEYINPUT75), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n390), .B(new_n460), .C1(new_n392), .C2(new_n381), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(KEYINPUT37), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n397), .A3(new_n409), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT38), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n380), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n455), .A2(new_n456), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n420), .A2(new_n422), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n443), .B1(new_n468), .B2(KEYINPUT39), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT39), .B1(new_n428), .B2(new_n422), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n420), .B2(new_n422), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n461), .A3(new_n397), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n399), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n398), .A2(KEYINPUT30), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n466), .B(new_n474), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n439), .A2(new_n444), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n445), .A3(new_n452), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n448), .A2(new_n481), .A3(new_n450), .ZN(new_n482));
  INV_X1    g281(.A(new_n478), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n476), .A2(new_n399), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n475), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n465), .A2(new_n479), .B1(new_n485), .B2(new_n380), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n448), .A2(new_n481), .A3(new_n450), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n487), .A2(new_n477), .A3(new_n478), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n379), .A2(new_n322), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n310), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(new_n323), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n478), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n451), .A2(new_n457), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n379), .A4(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n325), .A2(new_n486), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(KEYINPUT13), .Z(new_n499));
  XOR2_X1   g298(.A(KEYINPUT85), .B(G36gat), .Z(new_n500));
  OAI21_X1  g299(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n502));
  INV_X1    g301(.A(G29gat), .ZN(new_n503));
  INV_X1    g302(.A(G36gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n500), .A2(G29gat), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G43gat), .ZN(new_n508));
  INV_X1    g307(.A(G43gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G50gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT15), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n506), .A2(new_n515), .A3(KEYINPUT87), .A4(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n519));
  OAI21_X1  g318(.A(G29gat), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n501), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n513), .ZN(new_n523));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n511), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT85), .B(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n521), .B1(new_n503), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n516), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n517), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(G1gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT16), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n533), .A2(G1gat), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n536), .A2(new_n537), .A3(G8gat), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XOR2_X1   g338(.A(G15gat), .B(G22gat), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n534), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n535), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n532), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n538), .A2(new_n543), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n547), .A2(new_n527), .B1(new_n522), .B2(new_n525), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n548), .B2(new_n517), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n499), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT90), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(new_n499), .C1(new_n545), .C2(new_n549), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n532), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(KEYINPUT17), .A3(new_n517), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n546), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n549), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n498), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n551), .A2(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT18), .A4(new_n498), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT11), .B(G169gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n561), .B(new_n571), .C1(new_n564), .C2(new_n565), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n497), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT8), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n581), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n579), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT95), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(new_n595), .B2(new_n579), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n577), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n588), .A2(new_n589), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n591), .A3(new_n579), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT96), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n555), .A2(new_n556), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT96), .B1(new_n598), .B2(new_n599), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n532), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT97), .A4(new_n605), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n608), .A2(G190gat), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(G190gat), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n327), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n259), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(G190gat), .A3(new_n609), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(G218gat), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G57gat), .B(G64gat), .Z(new_n627));
  OR2_X1    g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n627), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G57gat), .B(G64gat), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n629), .B(new_n628), .C1(new_n634), .C2(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT91), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n635), .A3(KEYINPUT91), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n626), .B1(new_n640), .B2(KEYINPUT21), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n633), .A2(new_n635), .A3(KEYINPUT91), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT91), .B1(new_n633), .B2(new_n635), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT21), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n625), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n641), .B2(new_n646), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n624), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G183gat), .B(G211gat), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n650), .ZN(new_n654));
  INV_X1    g453(.A(new_n624), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n648), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n651), .B2(new_n656), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n546), .B1(new_n644), .B2(new_n645), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT92), .B(KEYINPUT93), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n657), .B2(new_n658), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n612), .A2(new_n616), .A3(new_n617), .A4(new_n621), .ZN(new_n666));
  OAI22_X1  g465(.A1(new_n590), .A2(new_n596), .B1(new_n642), .B2(new_n643), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n598), .A2(new_n599), .A3(new_n636), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n597), .A2(new_n600), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n644), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n669), .B2(new_n679), .ZN(new_n683));
  AOI211_X1 g482(.A(KEYINPUT98), .B(KEYINPUT10), .C1(new_n667), .C2(new_n668), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n677), .B1(new_n685), .B2(new_n671), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n639), .A2(new_n638), .B1(new_n598), .B2(new_n599), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n598), .A2(new_n599), .A3(new_n636), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n679), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT98), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n669), .A2(new_n682), .A3(new_n679), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n690), .A2(new_n691), .B1(new_n678), .B2(new_n680), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n671), .B(KEYINPUT99), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n673), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n676), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n686), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n623), .A2(new_n665), .A3(new_n666), .A4(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n576), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n482), .A2(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n482), .A2(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n534), .ZN(G1324gat));
  INV_X1    g505(.A(new_n701), .ZN(new_n707));
  INV_X1    g506(.A(new_n493), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n539), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT16), .B(G8gat), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n701), .A2(new_n493), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT42), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT42), .B2(new_n711), .ZN(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n701), .B2(new_n325), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n323), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n701), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n379), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n623), .A2(new_n666), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n673), .B(new_n676), .C1(new_n692), .C2(new_n672), .ZN(new_n722));
  INV_X1    g521(.A(new_n693), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n685), .A2(new_n723), .B1(new_n672), .B2(new_n670), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n676), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n721), .A2(new_n665), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n576), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n704), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n503), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n497), .B2(new_n721), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n325), .A2(new_n486), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT73), .B1(new_n319), .B2(new_n320), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n298), .A2(new_n307), .A3(new_n299), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n283), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n379), .A2(new_n322), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n736), .A2(new_n485), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT35), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n496), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(KEYINPUT44), .A3(new_n720), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n665), .B(KEYINPUT102), .Z(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(new_n575), .A3(new_n725), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n704), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n747), .ZN(G1328gat));
  NOR2_X1   g547(.A1(new_n493), .A2(new_n500), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n727), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT103), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n727), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n500), .B1(new_n746), .B2(new_n493), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(G1329gat));
  NAND2_X1  g558(.A1(new_n576), .A2(new_n726), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n509), .B1(new_n760), .B2(new_n323), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n325), .A2(new_n509), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n746), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n766), .B(new_n761), .C1(new_n746), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1330gat));
  NOR3_X1   g567(.A1(new_n760), .A2(G50gat), .A3(new_n379), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n732), .A2(new_n742), .A3(new_n380), .A4(new_n745), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G50gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n772), .A3(KEYINPUT48), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n771), .A2(new_n774), .A3(G50gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n771), .B2(G50gat), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n775), .A2(new_n776), .A3(new_n769), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(G1331gat));
  NAND4_X1  g578(.A1(new_n721), .A2(new_n575), .A3(new_n665), .A4(new_n725), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n497), .A2(KEYINPUT106), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT106), .B1(new_n497), .B2(new_n780), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n728), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n782), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n493), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(G1333gat));
  INV_X1    g590(.A(G71gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n783), .A2(new_n792), .A3(new_n492), .ZN(new_n793));
  OAI21_X1  g592(.A(G71gat), .B1(new_n786), .B2(new_n325), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT50), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1334gat));
  NOR2_X1   g598(.A1(new_n786), .A2(new_n379), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT107), .B(G78gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1335gat));
  INV_X1    g601(.A(new_n665), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n575), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT108), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n696), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n743), .A2(new_n728), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G85gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  INV_X1    g610(.A(new_n805), .ZN(new_n812));
  AND4_X1   g611(.A1(KEYINPUT51), .A2(new_n741), .A3(new_n720), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n721), .B1(new_n733), .B2(new_n740), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n814), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n725), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n728), .A2(new_n583), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n810), .A2(new_n811), .B1(new_n816), .B2(new_n817), .ZN(G1336gat));
  NOR3_X1   g617(.A1(new_n493), .A2(G92gat), .A3(new_n696), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT110), .Z(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n813), .B2(new_n815), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n732), .A2(new_n742), .A3(new_n708), .A4(new_n806), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G92gat), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT111), .B(new_n820), .C1(new_n813), .C2(new_n815), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n819), .B1(new_n813), .B2(new_n815), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n825), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1337gat));
  INV_X1    g631(.A(new_n325), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n743), .A2(new_n833), .A3(new_n806), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G99gat), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n323), .A2(G99gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n816), .B2(new_n836), .ZN(G1338gat));
  NAND4_X1  g636(.A1(new_n732), .A2(new_n742), .A3(new_n380), .A4(new_n806), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n379), .A2(G106gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n816), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g641(.A1(new_n573), .A2(new_n574), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n697), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n681), .B(new_n693), .C1(new_n683), .C2(new_n684), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n846), .B(KEYINPUT54), .C1(new_n692), .C2(new_n672), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n685), .A2(new_n848), .A3(new_n723), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n695), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n695), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n722), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n498), .B1(new_n557), .B2(new_n558), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n545), .A2(new_n549), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n855), .A2(new_n856), .B1(new_n857), .B2(new_n499), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n570), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n574), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n852), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n720), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n861), .B2(new_n696), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n725), .A2(KEYINPUT113), .A3(new_n574), .A4(new_n860), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n851), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n843), .A2(new_n868), .A3(new_n722), .A4(new_n853), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n720), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT114), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n845), .B1(new_n874), .B2(new_n744), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n728), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n736), .A2(new_n737), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n708), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n235), .A3(new_n843), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n323), .A2(new_n380), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n493), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n575), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(KEYINPUT115), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(KEYINPUT115), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(G1340gat));
  NOR2_X1   g686(.A1(new_n696), .A2(new_n239), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G120gat), .B1(new_n883), .B2(new_n696), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1341gat));
  INV_X1    g693(.A(G127gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n895), .A3(new_n665), .ZN(new_n896));
  INV_X1    g695(.A(new_n744), .ZN(new_n897));
  OAI21_X1  g696(.A(G127gat), .B1(new_n883), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1342gat));
  NOR4_X1   g698(.A1(new_n879), .A2(G134gat), .A3(new_n708), .A4(new_n721), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT56), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n883), .B2(new_n721), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1343gat));
  OAI211_X1 g702(.A(new_n380), .B(new_n325), .C1(new_n876), .C2(KEYINPUT121), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n875), .B2(new_n728), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n575), .A2(G141gat), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR4_X1   g707(.A1(new_n904), .A2(new_n906), .A3(new_n708), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT58), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n833), .A2(new_n708), .A3(new_n704), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n720), .A2(new_n862), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n861), .A2(new_n696), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n850), .A2(new_n914), .A3(new_n851), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n850), .B2(new_n851), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n575), .A2(new_n854), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n912), .B1(new_n919), .B2(new_n720), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n844), .B1(new_n920), .B2(new_n803), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n379), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT119), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n868), .A2(KEYINPUT118), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n850), .A2(new_n914), .A3(new_n851), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n843), .A2(new_n722), .A3(new_n853), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n929), .A2(new_n930), .B1(new_n696), .B2(new_n861), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n721), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n665), .B1(new_n932), .B2(new_n912), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n926), .B(new_n923), .C1(new_n933), .C2(new_n844), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n925), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n875), .B2(new_n380), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n911), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G141gat), .B1(new_n938), .B2(new_n575), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n910), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT120), .B(new_n911), .C1(new_n935), .C2(new_n937), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n843), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n909), .B1(new_n944), .B2(G141gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT58), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(G1344gat));
  NAND2_X1  g746(.A1(new_n911), .A2(new_n725), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n698), .A2(new_n575), .A3(new_n699), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT122), .ZN(new_n950));
  INV_X1    g749(.A(new_n933), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n698), .A2(new_n952), .A3(new_n575), .A4(new_n699), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT57), .B1(new_n954), .B2(new_n380), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n875), .A2(new_n380), .A3(new_n936), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n948), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT59), .B1(new_n958), .B2(new_n347), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n942), .A2(new_n725), .A3(new_n943), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n347), .A2(KEYINPUT59), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n904), .A2(new_n708), .A3(new_n906), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n347), .A3(new_n725), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1345gat));
  NAND3_X1  g764(.A1(new_n963), .A2(new_n337), .A3(new_n665), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n942), .A2(new_n744), .A3(new_n943), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n337), .ZN(G1346gat));
  NOR2_X1   g767(.A1(new_n904), .A2(new_n906), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n969), .A2(new_n338), .A3(new_n493), .A4(new_n720), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n942), .A2(new_n720), .A3(new_n943), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n338), .ZN(G1347gat));
  NOR2_X1   g771(.A1(new_n728), .A2(new_n493), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n875), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n878), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n247), .A3(new_n843), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n843), .A3(new_n882), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT123), .B1(new_n978), .B2(G169gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n983), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1348gat));
  NAND3_X1  g784(.A1(new_n974), .A2(new_n882), .A3(new_n725), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G176gat), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n725), .A2(new_n248), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n975), .B2(new_n988), .ZN(G1349gat));
  AND3_X1   g788(.A1(new_n665), .A2(new_n265), .A3(new_n267), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n875), .A2(new_n882), .A3(new_n744), .A4(new_n973), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n253), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  AOI22_X1  g793(.A1(new_n976), .A2(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n996));
  NOR2_X1   g795(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n997));
  AND2_X1   g796(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n996), .A2(new_n999), .ZN(G1350gat));
  NAND3_X1  g799(.A1(new_n976), .A2(new_n259), .A3(new_n720), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n974), .A2(new_n882), .A3(new_n720), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G190gat), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n1003), .A2(KEYINPUT61), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1003), .A2(KEYINPUT61), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(G1351gat));
  AND2_X1   g805(.A1(new_n325), .A2(new_n973), .ZN(new_n1007));
  AND3_X1   g806(.A1(new_n1007), .A2(new_n875), .A3(new_n380), .ZN(new_n1008));
  AOI21_X1  g807(.A(G197gat), .B1(new_n1008), .B2(new_n843), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n956), .A2(KEYINPUT127), .A3(new_n957), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  INV_X1    g810(.A(new_n957), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n955), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1010), .A2(new_n1007), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n575), .A2(new_n329), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(G1352gat));
  OAI21_X1  g816(.A(G204gat), .B1(new_n1014), .B2(new_n696), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1008), .A2(new_n330), .A3(new_n725), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1020));
  OR2_X1    g819(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(G1353gat));
  NAND3_X1  g821(.A1(new_n1008), .A2(new_n326), .A3(new_n665), .ZN(new_n1023));
  OAI211_X1 g822(.A(new_n665), .B(new_n1007), .C1(new_n955), .C2(new_n1012), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1024), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  OAI21_X1  g826(.A(G218gat), .B1(new_n1014), .B2(new_n721), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1008), .A2(new_n327), .A3(new_n720), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(G1355gat));
endmodule


