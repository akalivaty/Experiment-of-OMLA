//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n472), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n487), .A2(new_n492), .A3(G138), .A4(new_n472), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(new_n472), .B2(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT5), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(new_n505), .B1(new_n501), .B2(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  INV_X1    g091(.A(new_n511), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  INV_X1    g093(.A(new_n514), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n502), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n501), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n506), .A2(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n523), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n517), .A2(G90), .B1(G52), .B2(new_n519), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n508), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n508), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT73), .B(G43), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n519), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n511), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  AOI22_X1  g128(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n508), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(G91), .B2(new_n517), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n519), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT74), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n556), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND3_X1  g140(.A1(new_n506), .A2(G87), .A3(new_n510), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n524), .A2(KEYINPUT71), .A3(new_n525), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT71), .B1(new_n524), .B2(new_n525), .ZN(new_n570));
  NOR3_X1   g145(.A1(new_n569), .A2(new_n570), .A3(G74), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n568), .B1(new_n571), .B2(new_n508), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n506), .B2(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT76), .B1(new_n576), .B2(new_n508), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n524), .A2(G61), .A3(new_n525), .ZN(new_n578));
  INV_X1    g153(.A(new_n575), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(new_n581), .A3(G651), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n524), .A2(G86), .A3(new_n525), .A4(new_n510), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n577), .A2(new_n582), .A3(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  XNOR2_X1  g165(.A(KEYINPUT78), .B(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n517), .A2(new_n591), .B1(G47), .B2(new_n519), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(G290));
  NAND3_X1  g168(.A1(G301), .A2(KEYINPUT79), .A3(G868), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n511), .A2(KEYINPUT80), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(new_n511), .B2(new_n595), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT10), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT81), .B(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n526), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT79), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(G171), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n594), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G284));
  XOR2_X1   g185(.A(new_n609), .B(KEYINPUT82), .Z(G321));
  NOR2_X1   g186(.A1(G286), .A2(new_n606), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n606), .ZN(G297));
  AOI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n606), .ZN(G280));
  INV_X1    g190(.A(new_n605), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n547), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n606), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n605), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n478), .A2(G2104), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n476), .A2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n478), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2435), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2438), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(G14), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT84), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(KEYINPUT85), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n651), .B(new_n655), .C1(new_n657), .C2(new_n654), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n654), .A3(new_n650), .ZN(new_n659));
  INV_X1    g234(.A(new_n654), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n650), .A3(new_n652), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n634), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT86), .ZN(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n672), .A2(new_n673), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n669), .A2(new_n674), .A3(new_n671), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n673), .C2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(G1986), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT22), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G24), .ZN(new_n685));
  INV_X1    g260(.A(G290), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(G1986), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(G1986), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n476), .A2(G119), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n478), .A2(G131), .ZN(new_n691));
  NOR2_X1   g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT35), .B(G1991), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n688), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G23), .B(G288), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n684), .A2(G6), .ZN(new_n702));
  INV_X1    g277(.A(G305), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n684), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n684), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n684), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT34), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n698), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(KEYINPUT87), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n698), .B(new_n712), .C1(new_n716), .C2(KEYINPUT36), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n715), .A2(new_n717), .B1(new_n716), .B2(KEYINPUT36), .ZN(new_n718));
  NAND2_X1  g293(.A1(G164), .A2(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G27), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2078), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G16), .A2(G19), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n547), .B2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n722), .B1(new_n724), .B2(G1341), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n684), .B1(new_n538), .B2(new_n539), .ZN(new_n726));
  NOR2_X1   g301(.A1(G5), .A2(G16), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n726), .A2(G1961), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(G1961), .B1(new_n726), .B2(new_n727), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G29), .A2(G32), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT26), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n487), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G2105), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n733), .B(new_n735), .C1(G129), .C2(new_n476), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT27), .B(G1996), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT91), .Z(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n744), .A2(G2090), .B1(new_n721), .B2(new_n720), .ZN(new_n745));
  AND2_X1   g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n741), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT94), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n740), .A2(new_n745), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n478), .A2(G139), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n487), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n757), .C1(new_n472), .C2(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G33), .B(new_n759), .S(G29), .Z(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G2072), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n737), .A2(new_n738), .B1(new_n741), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G168), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G16), .B2(G21), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT92), .B(G1966), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n761), .B(new_n763), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n750), .A2(new_n751), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n633), .A2(new_n741), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n730), .A2(new_n754), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n765), .A2(new_n767), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n776));
  INV_X1    g351(.A(G20), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n778), .C1(new_n613), .C2(new_n684), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n744), .A2(G2090), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT95), .Z(new_n782));
  NOR4_X1   g357(.A1(new_n772), .A2(new_n774), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n478), .A2(G140), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT88), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n476), .A2(G128), .ZN(new_n786));
  NOR2_X1   g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n472), .B2(G116), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT89), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n741), .A2(G26), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT90), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT28), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G1341), .B2(new_n724), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n783), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT31), .B(G11), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n684), .A2(G4), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n616), .B2(new_n684), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1348), .Z(new_n805));
  NAND4_X1  g380(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n783), .A2(new_n802), .A3(new_n799), .A4(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n718), .B1(new_n806), .B2(new_n808), .ZN(G311));
  INV_X1    g384(.A(new_n718), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(G150));
  XNOR2_X1  g388(.A(KEYINPUT99), .B(G860), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(new_n508), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  INV_X1    g392(.A(G55), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n511), .A2(new_n817), .B1(new_n818), .B2(new_n514), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n814), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n605), .A2(new_n617), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT39), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n816), .A2(KEYINPUT97), .A3(new_n819), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT97), .B1(new_n816), .B2(new_n819), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n826), .A2(new_n547), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n547), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n825), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n821), .B1(new_n831), .B2(new_n814), .ZN(G145));
  INV_X1    g407(.A(G37), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n626), .B(new_n694), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n478), .A2(G142), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n476), .A2(G130), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n840), .B(new_n841), .C1(G118), .C2(new_n472), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n834), .B(new_n843), .Z(new_n844));
  NOR2_X1   g419(.A1(new_n759), .A2(KEYINPUT100), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n791), .A2(G164), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n790), .A2(new_n499), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n736), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n846), .A2(new_n847), .A3(new_n845), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n846), .A2(new_n847), .ZN(new_n853));
  INV_X1    g428(.A(new_n845), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n736), .B1(new_n855), .B2(new_n848), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n844), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n844), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n850), .B1(new_n849), .B2(new_n851), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n736), .A3(new_n848), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(G160), .B(new_n633), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n482), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n857), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n857), .A2(new_n866), .A3(new_n861), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n863), .B1(new_n861), .B2(new_n866), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n833), .B(new_n865), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n857), .A2(new_n866), .A3(new_n861), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(new_n863), .C1(new_n866), .C2(new_n861), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n873), .A2(KEYINPUT104), .A3(new_n833), .A4(new_n865), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT40), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G395));
  NAND2_X1  g454(.A1(new_n613), .A2(new_n616), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n560), .A2(new_n562), .B1(new_n600), .B2(new_n604), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n829), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n826), .A2(new_n547), .A3(new_n827), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT105), .B1(new_n828), .B2(new_n829), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n621), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n621), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n888), .ZN(new_n892));
  INV_X1    g467(.A(new_n621), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n880), .A2(new_n882), .A3(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NOR2_X1   g471(.A1(G299), .A2(new_n605), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n897), .B2(new_n881), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n887), .A2(new_n888), .A3(new_n621), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G303), .B(G288), .ZN(new_n902));
  NAND2_X1  g477(.A1(G290), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n590), .A3(new_n592), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n905), .A3(new_n703), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n703), .B1(new_n903), .B2(new_n905), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(KEYINPUT106), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G305), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(KEYINPUT106), .A3(new_n906), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n891), .A2(new_n901), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n891), .A2(new_n901), .B1(new_n911), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n816), .A2(new_n819), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(G868), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n891), .A2(new_n901), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n911), .A2(new_n915), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n606), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT107), .B1(new_n928), .B2(new_n922), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n923), .ZN(G331));
  INV_X1    g506(.A(new_n909), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n538), .A2(G286), .A3(new_n539), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G286), .B1(new_n538), .B2(new_n539), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n934), .A2(new_n935), .B1(new_n828), .B2(new_n829), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n884), .A2(new_n937), .A3(new_n886), .A4(new_n933), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n899), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n938), .A2(new_n936), .B1(new_n882), .B2(new_n880), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n936), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n883), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n899), .A2(new_n936), .A3(new_n938), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n909), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n945), .A3(new_n833), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n941), .A2(new_n945), .A3(new_n948), .A4(new_n833), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(KEYINPUT44), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(G397));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n499), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n468), .A2(G40), .A3(new_n473), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n790), .B(G2067), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n736), .B(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n694), .A2(new_n696), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n694), .A2(new_n696), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G1986), .B2(G290), .ZN(new_n968));
  INV_X1    g543(.A(G1986), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n686), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n961), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n508), .B1(new_n578), .B2(new_n579), .ZN(new_n972));
  OAI21_X1  g547(.A(G1981), .B1(new_n972), .B2(new_n585), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n974));
  INV_X1    g549(.A(G1981), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n577), .A2(new_n582), .A3(new_n975), .A4(new_n586), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(G1981), .C1(new_n972), .C2(new_n585), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n497), .B1(new_n486), .B2(new_n488), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n982), .B2(new_n494), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n959), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT49), .A4(new_n978), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n981), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(G1976), .B(new_n568), .C1(new_n571), .C2(new_n508), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(new_n984), .A3(KEYINPUT109), .A4(G8), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n984), .A2(G288), .A3(G8), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n991), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT114), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n989), .B(new_n999), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G166), .A2(new_n986), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(KEYINPUT108), .A2(KEYINPUT55), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G166), .B2(new_n986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n959), .B1(new_n983), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT50), .B(G1384), .C1(new_n982), .C2(new_n494), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT112), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n956), .A2(KEYINPUT50), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n983), .A2(new_n1009), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n959), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G2090), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n983), .A2(KEYINPUT45), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n958), .A2(new_n959), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n709), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G8), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1019), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1008), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1017), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n986), .B1(new_n1028), .B2(new_n1022), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1007), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1001), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1013), .A2(new_n751), .A3(new_n959), .A4(new_n1015), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n983), .A2(KEYINPUT45), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n957), .B(G1384), .C1(new_n982), .C2(new_n494), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n960), .ZN(new_n1035));
  OAI211_X1 g610(.A(G168), .B(new_n1032), .C1(new_n1035), .C2(new_n766), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1041), .A3(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT120), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n751), .A2(new_n1027), .B1(new_n1021), .B2(new_n767), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n986), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G286), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(KEYINPUT120), .A3(KEYINPUT51), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT121), .B(G1961), .Z(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n958), .A2(new_n721), .A3(new_n959), .A4(new_n1020), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1051), .B(KEYINPUT122), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1033), .A2(new_n1034), .A3(G2078), .ZN(new_n1061));
  XOR2_X1   g636(.A(new_n473), .B(KEYINPUT123), .Z(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1053), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(G40), .A3(new_n468), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1057), .A3(new_n1051), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(G171), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(G171), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT54), .B(new_n1070), .C1(new_n1059), .C2(G171), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1031), .A2(new_n1049), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT54), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1042), .A2(KEYINPUT120), .A3(KEYINPUT51), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1043), .B2(new_n1040), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1077), .B2(new_n1047), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT124), .A3(new_n1031), .A4(new_n1071), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n605), .B(new_n1080), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1027), .A2(G1348), .B1(G2067), .B2(new_n984), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT118), .B(new_n605), .C1(new_n1082), .C2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(new_n1086), .C1(KEYINPUT60), .C2(new_n1083), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n559), .B1(KEYINPUT116), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(KEYINPUT116), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1027), .A2(G1956), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1035), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1090), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1089), .B(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1095), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(KEYINPUT61), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT58), .B(G1341), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1021), .A2(G1996), .B1(new_n985), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n547), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT59), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1087), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1091), .A2(KEYINPUT117), .A3(new_n1096), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT61), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1099), .A2(new_n1095), .B1(new_n616), .B2(new_n1082), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1106), .A2(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1074), .A2(new_n1079), .A3(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1045), .A2(new_n986), .A3(G286), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1001), .A2(new_n1026), .A3(new_n1030), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT115), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1030), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n998), .B2(new_n1000), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1026), .A4(new_n1115), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n997), .B(KEYINPUT111), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1029), .A2(new_n1007), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(new_n1115), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(new_n1126), .A3(KEYINPUT63), .A4(new_n1030), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n989), .A2(new_n992), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n976), .B1(new_n1129), .B2(G288), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1124), .A2(new_n1119), .B1(new_n1130), .B2(new_n987), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1077), .A2(new_n1132), .A3(new_n1047), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1049), .A2(KEYINPUT62), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1060), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1031), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1128), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n971), .B1(new_n1114), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n686), .A2(new_n969), .A3(new_n961), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT48), .ZN(new_n1140));
  INV_X1    g715(.A(new_n961), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n967), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n964), .A2(new_n696), .A3(new_n694), .ZN(new_n1143));
  INV_X1    g718(.A(G2067), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n790), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n962), .B2(new_n736), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT125), .Z(new_n1148));
  NOR2_X1   g723(.A1(new_n1141), .A2(G1996), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1146), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1138), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g733(.A1(G229), .A2(G401), .A3(G227), .ZN(new_n1160));
  NAND4_X1  g734(.A1(new_n950), .A2(new_n875), .A3(G319), .A4(new_n1160), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


