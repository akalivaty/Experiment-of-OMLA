//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT67), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n466), .A2(KEYINPUT3), .A3(new_n467), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n480), .A2(G137), .A3(new_n469), .A4(new_n476), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n472), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  INV_X1    g058(.A(G100), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n484), .A2(new_n469), .A3(KEYINPUT69), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n484), .B2(new_n469), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n480), .A2(new_n476), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n469), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(G2105), .ZN(new_n492));
  OAI221_X1 g067(.A(new_n487), .B1(new_n489), .B2(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT70), .ZN(G162));
  NAND2_X1  g069(.A1(new_n476), .A2(new_n477), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n469), .A3(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n469), .A2(G138), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n480), .A2(new_n476), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n480), .A2(G126), .A3(G2105), .A4(new_n476), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n469), .A2(KEYINPUT71), .A3(G114), .ZN(new_n507));
  OAI211_X1 g082(.A(G2104), .B(new_n503), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n501), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(new_n515), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(G543), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(new_n524), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n521), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n527), .B(new_n529), .C1(new_n533), .C2(KEYINPUT73), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(G651), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n521), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G90), .B1(G52), .B2(new_n528), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n518), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n521), .A2(new_n548), .B1(new_n549), .B2(new_n524), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT75), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT76), .Z(G188));
  NAND2_X1  g133(.A1(new_n521), .A2(KEYINPUT77), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n516), .A2(new_n560), .A3(new_n520), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(G91), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n516), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n516), .A2(new_n568), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n566), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  OR2_X1    g152(.A1(G166), .A2(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g153(.A1(G166), .A2(KEYINPUT79), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G303));
  OR2_X1    g155(.A1(new_n516), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(G49), .B2(new_n528), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n559), .A2(G87), .A3(new_n561), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n516), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G48), .B2(new_n528), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n559), .A2(new_n561), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n518), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n521), .A2(new_n594), .B1(new_n595), .B2(new_n524), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(new_n571), .ZN(new_n600));
  OAI21_X1  g175(.A(G66), .B1(new_n600), .B2(new_n569), .ZN(new_n601));
  INV_X1    g176(.A(G79), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n511), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n559), .A2(G92), .A3(new_n561), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G280));
  INV_X1    g190(.A(G860), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n608), .B1(G559), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(G148));
  OAI21_X1  g193(.A(KEYINPUT82), .B1(new_n551), .B2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  MUX2_X1   g197(.A(KEYINPUT82), .B(new_n619), .S(new_n622), .Z(G323));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n627));
  INV_X1    g202(.A(new_n489), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G135), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n630));
  INV_X1    g205(.A(new_n492), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G123), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n492), .A2(KEYINPUT85), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n627), .B(new_n629), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n470), .A2(new_n495), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(KEYINPUT84), .B(G2100), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT89), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n663), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n661), .B(new_n669), .C1(new_n664), .C2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n661), .A2(new_n663), .A3(new_n666), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n682), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n684), .B(new_n687), .C1(new_n679), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT91), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(G229));
  NAND3_X1  g271(.A1(new_n476), .A2(new_n477), .A3(G127), .ZN(new_n697));
  NAND2_X1  g272(.A1(G115), .A2(G2104), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n469), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n628), .A2(G139), .B1(new_n699), .B2(KEYINPUT98), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT97), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT25), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n703), .C1(KEYINPUT98), .C2(new_n699), .ZN(new_n704));
  MUX2_X1   g279(.A(G33), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(new_n442), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n628), .A2(G141), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n631), .A2(G129), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n471), .A2(G105), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n709), .A2(new_n710), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n708), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G27), .A2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G164), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n443), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n551), .B2(new_n726), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n728), .A2(G1341), .B1(G2078), .B2(new_n723), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(G1341), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n718), .B2(new_n720), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n706), .A2(new_n725), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G28), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n707), .B1(new_n733), .B2(G28), .ZN(new_n735));
  AND2_X1   g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  NOR2_X1   g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n635), .A2(new_n707), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT24), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n482), .B2(new_n707), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n740), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT99), .Z(new_n747));
  OAI21_X1  g322(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n750));
  OAI221_X1 g325(.A(G2104), .B1(G116), .B2(new_n469), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G140), .ZN(new_n752));
  INV_X1    g327(.A(G128), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n751), .B1(new_n489), .B2(new_n752), .C1(new_n753), .C2(new_n492), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n707), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n745), .A2(new_n747), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n726), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n726), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1966), .ZN(new_n764));
  NOR2_X1   g339(.A1(G5), .A2(G16), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G171), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1961), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n732), .A2(new_n761), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n609), .A2(new_n726), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G4), .B2(new_n726), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT94), .B(G1348), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n770), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n726), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G35), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G162), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT29), .ZN(new_n783));
  INV_X1    g358(.A(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n768), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT100), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n726), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n726), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1971), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n726), .A2(G6), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G305), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT32), .B(G1981), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n794), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n790), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(G16), .A2(G23), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n582), .A2(new_n583), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(G288), .A2(KEYINPUT92), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n803), .B2(new_n726), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT33), .B(G1976), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n797), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n806), .B2(new_n804), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n628), .A2(G131), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n631), .A2(G119), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n469), .A2(G107), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G25), .B(new_n816), .S(G29), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n726), .A2(G24), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n597), .B2(new_n726), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1986), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n811), .A2(KEYINPUT93), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT93), .B1(new_n811), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n810), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(new_n810), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n787), .B1(new_n828), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(new_n787), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(G150));
  AOI22_X1  g409(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n518), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n521), .A2(new_n837), .B1(new_n838), .B2(new_n524), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n616), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n609), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n551), .B(new_n840), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  OAI21_X1  g423(.A(new_n616), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n842), .B1(new_n848), .B2(new_n849), .ZN(G145));
  NOR2_X1   g425(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n716), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n754), .B(G164), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n816), .B(new_n639), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n631), .A2(G130), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n628), .A2(G142), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n855), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n854), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(G162), .B(new_n482), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n635), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n869), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g449(.A(new_n612), .B1(new_n836), .B2(new_n839), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n803), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(G166), .B(new_n597), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT42), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(KEYINPUT105), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n621), .B(new_n845), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n608), .A2(G299), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n608), .A2(G299), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT41), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n881), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n880), .A2(new_n890), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n891), .A2(new_n892), .B1(KEYINPUT105), .B2(new_n879), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n875), .B1(new_n893), .B2(new_n612), .ZN(G295));
  OAI21_X1  g469(.A(new_n875), .B1(new_n893), .B2(new_n612), .ZN(G331));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n896));
  XOR2_X1   g471(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n897));
  NOR2_X1   g472(.A1(G171), .A2(KEYINPUT108), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n845), .ZN(new_n899));
  AOI21_X1  g474(.A(G286), .B1(G171), .B2(KEYINPUT108), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n887), .A2(new_n885), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n889), .A3(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n878), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n907), .A2(new_n871), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  INV_X1    g484(.A(new_n878), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n897), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n871), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n885), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n885), .A2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n887), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n903), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n878), .B1(new_n918), .B2(new_n906), .ZN(new_n919));
  INV_X1    g494(.A(new_n897), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n913), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n896), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n908), .A2(new_n911), .A3(new_n897), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n913), .B2(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(KEYINPUT44), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n501), .B2(new_n509), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n472), .A2(new_n479), .A3(G40), .A4(new_n481), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n754), .B(new_n759), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(new_n717), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT46), .B1(new_n934), .B2(G1996), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n934), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n935), .A2(new_n934), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT110), .Z(new_n943));
  INV_X1    g518(.A(new_n934), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n716), .B(G1996), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n816), .A2(new_n819), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n754), .A2(G2067), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n934), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n816), .A2(new_n819), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n951), .B2(new_n947), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n934), .A2(G1986), .A3(G290), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT48), .Z(new_n955));
  AOI211_X1 g530(.A(new_n941), .B(new_n950), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(KEYINPUT45), .B(new_n927), .C1(new_n501), .C2(new_n509), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n930), .A2(new_n933), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n959));
  INV_X1    g534(.A(G1971), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n930), .A2(new_n933), .A3(new_n961), .A4(new_n957), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n928), .A2(KEYINPUT112), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(new_n927), .C1(new_n501), .C2(new_n509), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n933), .B1(KEYINPUT50), .B2(new_n928), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n784), .A3(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n963), .A2(KEYINPUT116), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT116), .B1(new_n963), .B2(new_n971), .ZN(new_n973));
  INV_X1    g548(.A(G8), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n578), .A2(G8), .A3(new_n579), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n976), .A2(KEYINPUT113), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT117), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n801), .A2(G1976), .A3(new_n802), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n964), .A2(new_n933), .A3(new_n966), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(G8), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT52), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n588), .B1(new_n590), .B2(new_n521), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G1981), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n588), .B(new_n989), .C1(new_n590), .C2(new_n589), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n988), .B(new_n990), .C1(KEYINPUT114), .C2(KEYINPUT49), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(G8), .A3(new_n994), .A4(new_n984), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n983), .A2(G8), .A3(new_n984), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n986), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n964), .A2(new_n1000), .A3(new_n966), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n932), .B1(new_n928), .B2(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n784), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n974), .B1(new_n963), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n999), .B1(new_n981), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n963), .A2(new_n971), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n963), .A2(KEYINPUT116), .A3(new_n971), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(G8), .A3(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT119), .B(G2084), .Z(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n967), .A2(new_n929), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(KEYINPUT118), .A3(new_n933), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT45), .B1(new_n964), .B2(new_n966), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n932), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1021), .A3(new_n957), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1024), .A2(new_n974), .A3(G286), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n982), .A2(new_n1005), .A3(new_n1013), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n981), .A2(new_n1004), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1005), .A2(KEYINPUT63), .A3(new_n1029), .A4(new_n1025), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2078), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1022), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1961), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1014), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G2078), .B1(new_n959), .B2(new_n962), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(KEYINPUT53), .ZN(new_n1039));
  OAI21_X1  g614(.A(G171), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AND4_X1   g616(.A1(new_n982), .A2(new_n1005), .A3(new_n1041), .A4(new_n1013), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G168), .A2(new_n974), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1043), .B2(KEYINPUT124), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1046), .C1(new_n1024), .C2(new_n974), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1024), .A2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n974), .B(new_n1046), .C1(new_n1024), .C2(G168), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT62), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n974), .B1(new_n1024), .B2(G168), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1046), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1048), .A4(new_n1047), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1042), .A2(new_n1051), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n981), .A2(new_n1004), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n999), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n984), .A2(G8), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n995), .A2(new_n996), .A3(new_n799), .ZN(new_n1061));
  XOR2_X1   g636(.A(new_n990), .B(KEYINPUT115), .Z(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1031), .A2(new_n1057), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n958), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1014), .A2(new_n1036), .B1(new_n1066), .B2(new_n1033), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(G301), .C1(new_n1038), .C2(KEYINPUT53), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT125), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1038), .A2(KEYINPUT53), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(G301), .A4(new_n1067), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1040), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(new_n1067), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(G171), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1035), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1039), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(G301), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1073), .A2(new_n1074), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1054), .A2(new_n1048), .A3(new_n1047), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n982), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1083), .A2(KEYINPUT126), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND3_X1  g660(.A1(new_n984), .A2(KEYINPUT121), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(G1996), .B2(new_n958), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT121), .B1(new_n984), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n551), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n551), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n566), .A2(new_n575), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(G65), .B1(new_n600), .B2(new_n569), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n518), .B1(new_n1097), .B2(new_n573), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT57), .B1(new_n1098), .B2(new_n565), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1066), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1000), .B1(new_n964), .B2(new_n966), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n778), .B1(new_n1104), .B2(new_n969), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1094), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n1105), .A3(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1093), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1100), .A2(new_n1105), .A3(KEYINPUT120), .A4(new_n1103), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT61), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT122), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1090), .A2(new_n1092), .B1(new_n1108), .B2(new_n1107), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1112), .A2(new_n1113), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(new_n1119), .C1(KEYINPUT61), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1348), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n984), .A2(G2067), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1122), .B1(new_n1126), .B2(new_n609), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1122), .A3(new_n609), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1128), .A2(new_n1129), .B1(KEYINPUT60), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1129), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(KEYINPUT60), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1127), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1117), .A2(new_n1121), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1115), .B1(new_n608), .B2(new_n1130), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1114), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1083), .A2(KEYINPUT126), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1065), .B1(new_n1084), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n597), .B(G1986), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n953), .B1(new_n934), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n956), .B1(new_n1140), .B2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g718(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1145));
  OAI211_X1 g719(.A(new_n873), .B(new_n1145), .C1(new_n912), .C2(new_n921), .ZN(G225));
  INV_X1    g720(.A(G225), .ZN(G308));
endmodule


