

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751;

  AND2_X1 U372 ( .A1(n417), .A2(n409), .ZN(n652) );
  XNOR2_X2 U373 ( .A(n432), .B(G143), .ZN(n501) );
  XNOR2_X2 U374 ( .A(G128), .B(KEYINPUT66), .ZN(n432) );
  NOR2_X1 U375 ( .A1(n746), .A2(n744), .ZN(n608) );
  XNOR2_X1 U376 ( .A(n394), .B(n393), .ZN(n750) );
  NAND2_X1 U377 ( .A1(n562), .A2(n571), .ZN(n672) );
  INV_X1 U378 ( .A(n591), .ZN(n348) );
  XNOR2_X1 U379 ( .A(n554), .B(n374), .ZN(n591) );
  INV_X1 U380 ( .A(KEYINPUT92), .ZN(n462) );
  INV_X1 U381 ( .A(KEYINPUT68), .ZN(n455) );
  XNOR2_X1 U382 ( .A(n437), .B(n364), .ZN(n370) );
  NOR2_X1 U383 ( .A1(n431), .A2(n573), .ZN(n397) );
  NOR2_X1 U384 ( .A1(n750), .A2(n655), .ZN(n564) );
  NOR2_X1 U385 ( .A1(n585), .A2(n584), .ZN(n667) );
  XNOR2_X1 U386 ( .A(n464), .B(n463), .ZN(n744) );
  AND2_X1 U387 ( .A1(n665), .A2(n674), .ZN(n378) );
  NAND2_X1 U388 ( .A1(n426), .A2(n359), .ZN(n394) );
  XNOR2_X1 U389 ( .A(n456), .B(KEYINPUT19), .ZN(n586) );
  XNOR2_X1 U390 ( .A(n615), .B(KEYINPUT38), .ZN(n459) );
  NAND2_X1 U391 ( .A1(n425), .A2(n670), .ZN(n456) );
  XNOR2_X1 U392 ( .A(n543), .B(n493), .ZN(n377) );
  XNOR2_X1 U393 ( .A(n454), .B(n735), .ZN(n543) );
  XNOR2_X1 U394 ( .A(n399), .B(n496), .ZN(n724) );
  XNOR2_X1 U395 ( .A(n501), .B(n488), .ZN(n534) );
  XNOR2_X1 U396 ( .A(n455), .B(G101), .ZN(n454) );
  XNOR2_X1 U397 ( .A(n495), .B(n494), .ZN(n399) );
  XNOR2_X1 U398 ( .A(n533), .B(G137), .ZN(n469) );
  XNOR2_X1 U399 ( .A(n467), .B(n466), .ZN(n493) );
  XNOR2_X1 U400 ( .A(n499), .B(n462), .ZN(n461) );
  XNOR2_X1 U401 ( .A(G902), .B(KEYINPUT15), .ZN(n621) );
  XNOR2_X1 U402 ( .A(G119), .B(KEYINPUT72), .ZN(n467) );
  XNOR2_X1 U403 ( .A(G116), .B(KEYINPUT3), .ZN(n466) );
  INV_X1 U404 ( .A(G953), .ZN(n446) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(G131), .Z(n533) );
  INV_X1 U406 ( .A(n585), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n588), .B(KEYINPUT1), .ZN(n559) );
  NOR2_X1 U408 ( .A1(n606), .A2(n590), .ZN(n660) );
  OR2_X1 U409 ( .A1(n606), .A2(n697), .ZN(n464) );
  BUF_X1 U410 ( .A(n665), .Z(n350) );
  XNOR2_X1 U411 ( .A(n379), .B(KEYINPUT31), .ZN(n665) );
  AND2_X2 U412 ( .A1(n424), .A2(n636), .ZN(n385) );
  BUF_X2 U413 ( .A(n566), .Z(n747) );
  AND2_X2 U414 ( .A1(n381), .A2(n355), .ZN(n390) );
  NOR2_X2 U415 ( .A1(n705), .A2(G902), .ZN(n547) );
  XNOR2_X2 U416 ( .A(n732), .B(n545), .ZN(n705) );
  XNOR2_X2 U417 ( .A(n553), .B(n535), .ZN(n732) );
  NAND2_X1 U418 ( .A1(n674), .A2(n660), .ZN(n376) );
  NOR2_X1 U419 ( .A1(n564), .A2(n555), .ZN(n556) );
  XNOR2_X1 U420 ( .A(n405), .B(n575), .ZN(n404) );
  INV_X1 U421 ( .A(G469), .ZN(n546) );
  XNOR2_X1 U422 ( .A(n377), .B(n551), .ZN(n552) );
  INV_X1 U423 ( .A(KEYINPUT6), .ZN(n391) );
  NAND2_X1 U424 ( .A1(n448), .A2(n447), .ZN(n578) );
  AND2_X1 U425 ( .A1(n452), .A2(n451), .ZN(n448) );
  NAND2_X1 U426 ( .A1(n351), .A2(n450), .ZN(n447) );
  INV_X1 U427 ( .A(KEYINPUT22), .ZN(n395) );
  INV_X1 U428 ( .A(KEYINPUT77), .ZN(n366) );
  NAND2_X1 U429 ( .A1(n370), .A2(n356), .ZN(n369) );
  NAND2_X1 U430 ( .A1(n440), .A2(n599), .ZN(n439) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n440) );
  AND2_X1 U432 ( .A1(n389), .A2(n578), .ZN(n684) );
  INV_X1 U433 ( .A(n558), .ZN(n389) );
  XNOR2_X1 U434 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U435 ( .A(n576), .B(KEYINPUT45), .ZN(n577) );
  XNOR2_X1 U436 ( .A(n401), .B(n460), .ZN(n400) );
  XNOR2_X1 U437 ( .A(n497), .B(n498), .ZN(n460) );
  XNOR2_X1 U438 ( .A(n461), .B(n500), .ZN(n401) );
  AND2_X1 U439 ( .A1(n420), .A2(n596), .ZN(n419) );
  NAND2_X1 U440 ( .A1(n557), .A2(n561), .ZN(n420) );
  XNOR2_X1 U441 ( .A(n487), .B(n486), .ZN(n518) );
  XOR2_X1 U442 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n486) );
  XNOR2_X1 U443 ( .A(n485), .B(KEYINPUT83), .ZN(n487) );
  NAND2_X1 U444 ( .A1(n446), .A2(G234), .ZN(n485) );
  INV_X1 U445 ( .A(G134), .ZN(n488) );
  XNOR2_X1 U446 ( .A(n490), .B(G116), .ZN(n442) );
  INV_X1 U447 ( .A(n718), .ZN(n413) );
  XNOR2_X1 U448 ( .A(n384), .B(n605), .ZN(n697) );
  NOR2_X1 U449 ( .A1(n675), .A2(n672), .ZN(n384) );
  NOR2_X1 U450 ( .A1(n355), .A2(n585), .ZN(n465) );
  AND2_X1 U451 ( .A1(n595), .A2(n594), .ZN(n600) );
  XNOR2_X1 U452 ( .A(n371), .B(KEYINPUT28), .ZN(n589) );
  NOR2_X1 U453 ( .A1(n348), .A2(n587), .ZN(n371) );
  AND2_X1 U454 ( .A1(n380), .A2(n348), .ZN(n417) );
  NAND2_X1 U455 ( .A1(n417), .A2(n416), .ZN(n569) );
  NOR2_X1 U456 ( .A1(n355), .A2(n458), .ZN(n457) );
  NAND2_X1 U457 ( .A1(n585), .A2(n578), .ZN(n458) );
  OR2_X2 U458 ( .A1(n652), .A2(n378), .ZN(n431) );
  OR2_X1 U459 ( .A1(n620), .A2(KEYINPUT77), .ZN(n368) );
  INV_X1 U460 ( .A(KEYINPUT47), .ZN(n375) );
  XNOR2_X1 U461 ( .A(G143), .B(G122), .ZN(n478) );
  NAND2_X1 U462 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X1 U463 ( .A(KEYINPUT73), .B(G110), .ZN(n540) );
  XNOR2_X1 U464 ( .A(G104), .B(G107), .ZN(n539) );
  XOR2_X1 U465 ( .A(KEYINPUT78), .B(KEYINPUT96), .Z(n537) );
  INV_X1 U466 ( .A(KEYINPUT95), .ZN(n535) );
  NAND2_X1 U467 ( .A1(n459), .A2(n670), .ZN(n675) );
  INV_X1 U468 ( .A(KEYINPUT76), .ZN(n382) );
  NAND2_X1 U469 ( .A1(n373), .A2(n372), .ZN(n587) );
  XNOR2_X1 U470 ( .A(n388), .B(n387), .ZN(n595) );
  INV_X1 U471 ( .A(KEYINPUT100), .ZN(n387) );
  INV_X1 U472 ( .A(n532), .ZN(n453) );
  INV_X1 U473 ( .A(G902), .ZN(n449) );
  XNOR2_X1 U474 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U475 ( .A(G119), .B(G137), .ZN(n522) );
  NAND2_X1 U476 ( .A1(n413), .A2(n411), .ZN(n636) );
  NOR2_X1 U477 ( .A1(n625), .A2(n412), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n398), .B(n402), .ZN(n629) );
  XNOR2_X1 U479 ( .A(n400), .B(n724), .ZN(n398) );
  INV_X1 U480 ( .A(KEYINPUT114), .ZN(n436) );
  NAND2_X1 U481 ( .A1(n353), .A2(n383), .ZN(n563) );
  INV_X1 U482 ( .A(G472), .ZN(n374) );
  NOR2_X1 U483 ( .A1(n639), .A2(G902), .ZN(n554) );
  INV_X1 U484 ( .A(n493), .ZN(n725) );
  AND2_X1 U485 ( .A1(n444), .A2(G953), .ZN(n729) );
  INV_X1 U486 ( .A(G898), .ZN(n444) );
  XNOR2_X1 U487 ( .A(n443), .B(n441), .ZN(n712) );
  XNOR2_X1 U488 ( .A(n491), .B(n489), .ZN(n443) );
  NAND2_X1 U489 ( .A1(n385), .A2(G475), .ZN(n647) );
  XNOR2_X1 U490 ( .A(n645), .B(KEYINPUT59), .ZN(n646) );
  NAND2_X1 U491 ( .A1(n385), .A2(G210), .ZN(n631) );
  XNOR2_X1 U492 ( .A(KEYINPUT91), .B(n632), .ZN(n704) );
  AND2_X1 U493 ( .A1(n445), .A2(G953), .ZN(n632) );
  INV_X1 U494 ( .A(G952), .ZN(n445) );
  NAND2_X1 U495 ( .A1(n413), .A2(n410), .ZN(n414) );
  INV_X1 U496 ( .A(n625), .ZN(n410) );
  XNOR2_X1 U497 ( .A(n607), .B(KEYINPUT113), .ZN(n463) );
  INV_X1 U498 ( .A(KEYINPUT32), .ZN(n393) );
  XNOR2_X1 U499 ( .A(n569), .B(n415), .ZN(n653) );
  INV_X1 U500 ( .A(KEYINPUT27), .ZN(n415) );
  INV_X1 U501 ( .A(n570), .ZN(n651) );
  AND2_X1 U502 ( .A1(n532), .A2(n449), .ZN(n351) );
  AND2_X1 U503 ( .A1(n369), .A2(n362), .ZN(n352) );
  AND2_X1 U504 ( .A1(n418), .A2(n419), .ZN(n353) );
  XNOR2_X1 U505 ( .A(n503), .B(KEYINPUT81), .ZN(n354) );
  XOR2_X1 U506 ( .A(n348), .B(n391), .Z(n355) );
  AND2_X1 U507 ( .A1(n620), .A2(KEYINPUT77), .ZN(n356) );
  AND2_X1 U508 ( .A1(n352), .A2(n365), .ZN(n357) );
  INV_X1 U509 ( .A(n578), .ZN(n373) );
  AND2_X1 U510 ( .A1(n582), .A2(n581), .ZN(n358) );
  AND2_X1 U511 ( .A1(n465), .A2(n373), .ZN(n359) );
  NOR2_X1 U512 ( .A1(n386), .A2(n697), .ZN(n360) );
  NOR2_X1 U513 ( .A1(n680), .A2(n386), .ZN(n361) );
  AND2_X1 U514 ( .A1(n368), .A2(n429), .ZN(n362) );
  AND2_X1 U515 ( .A1(n585), .A2(n373), .ZN(n363) );
  INV_X1 U516 ( .A(n656), .ZN(n416) );
  INV_X1 U517 ( .A(n659), .ZN(n409) );
  XNOR2_X1 U518 ( .A(n610), .B(KEYINPUT86), .ZN(n364) );
  INV_X1 U519 ( .A(KEYINPUT2), .ZN(n412) );
  NAND2_X1 U520 ( .A1(n370), .A2(n620), .ZN(n625) );
  INV_X1 U521 ( .A(n370), .ZN(n367) );
  NOR2_X1 U522 ( .A1(n681), .A2(n358), .ZN(n372) );
  XNOR2_X1 U523 ( .A(n377), .B(n502), .ZN(n402) );
  NAND2_X1 U524 ( .A1(n689), .A2(n422), .ZN(n379) );
  XNOR2_X1 U525 ( .A(n568), .B(KEYINPUT101), .ZN(n380) );
  AND2_X1 U526 ( .A1(n381), .A2(n591), .ZN(n689) );
  XNOR2_X2 U527 ( .A(n468), .B(n382), .ZN(n381) );
  OR2_X1 U528 ( .A1(n386), .A2(n421), .ZN(n383) );
  XNOR2_X2 U529 ( .A(n390), .B(n560), .ZN(n386) );
  NAND2_X1 U530 ( .A1(n385), .A2(G469), .ZN(n708) );
  NAND2_X1 U531 ( .A1(n385), .A2(G478), .ZN(n711) );
  NAND2_X1 U532 ( .A1(n385), .A2(G217), .ZN(n715) );
  NAND2_X1 U533 ( .A1(n386), .A2(n561), .ZN(n418) );
  NAND2_X1 U534 ( .A1(n588), .A2(n684), .ZN(n388) );
  AND2_X1 U535 ( .A1(n426), .A2(n392), .ZN(n655) );
  AND2_X1 U536 ( .A1(n363), .A2(n348), .ZN(n392) );
  XNOR2_X2 U537 ( .A(n396), .B(n395), .ZN(n426) );
  XNOR2_X1 U538 ( .A(n433), .B(KEYINPUT36), .ZN(n584) );
  XNOR2_X1 U539 ( .A(n611), .B(n436), .ZN(n435) );
  NAND2_X1 U540 ( .A1(n516), .A2(n517), .ZN(n396) );
  NAND2_X1 U541 ( .A1(n574), .A2(n397), .ZN(n405) );
  NAND2_X1 U542 ( .A1(n435), .A2(n434), .ZN(n433) );
  NOR2_X1 U543 ( .A1(n747), .A2(KEYINPUT44), .ZN(n565) );
  INV_X2 U544 ( .A(n557), .ZN(n422) );
  NAND2_X1 U545 ( .A1(n430), .A2(n357), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n403), .B(n577), .ZN(n624) );
  NOR2_X2 U547 ( .A1(n406), .A2(n404), .ZN(n403) );
  NAND2_X1 U548 ( .A1(n408), .A2(n407), .ZN(n406) );
  XNOR2_X1 U549 ( .A(n556), .B(KEYINPUT67), .ZN(n407) );
  NAND2_X1 U550 ( .A1(n565), .A2(n564), .ZN(n408) );
  XNOR2_X1 U551 ( .A(n414), .B(n412), .ZN(n701) );
  NAND2_X1 U552 ( .A1(n422), .A2(n423), .ZN(n421) );
  INV_X1 U553 ( .A(n561), .ZN(n423) );
  NAND2_X1 U554 ( .A1(n637), .A2(n424), .ZN(n641) );
  NAND2_X1 U555 ( .A1(n427), .A2(n623), .ZN(n424) );
  INV_X1 U556 ( .A(n425), .ZN(n615) );
  XNOR2_X2 U557 ( .A(n504), .B(n354), .ZN(n425) );
  AND2_X1 U558 ( .A1(n425), .A2(n596), .ZN(n597) );
  NAND2_X1 U559 ( .A1(n426), .A2(n457), .ZN(n570) );
  XNOR2_X1 U560 ( .A(n428), .B(KEYINPUT84), .ZN(n427) );
  INV_X1 U561 ( .A(n621), .ZN(n429) );
  INV_X1 U562 ( .A(n624), .ZN(n430) );
  NAND2_X1 U563 ( .A1(n586), .A2(n512), .ZN(n513) );
  INV_X1 U564 ( .A(n456), .ZN(n434) );
  NAND2_X1 U565 ( .A1(n583), .A2(n355), .ZN(n611) );
  NAND2_X1 U566 ( .A1(n438), .A2(n609), .ZN(n437) );
  NOR2_X1 U567 ( .A1(n667), .A2(n439), .ZN(n438) );
  XNOR2_X1 U568 ( .A(n534), .B(n442), .ZN(n441) );
  NAND2_X1 U569 ( .A1(n446), .A2(G227), .ZN(n536) );
  AND2_X1 U570 ( .A1(n446), .A2(G224), .ZN(n497) );
  NAND2_X1 U571 ( .A1(n737), .A2(n446), .ZN(n743) );
  INV_X1 U572 ( .A(n714), .ZN(n450) );
  NAND2_X1 U573 ( .A1(n453), .A2(G902), .ZN(n451) );
  NAND2_X1 U574 ( .A1(n714), .A2(n453), .ZN(n452) );
  XNOR2_X2 U575 ( .A(KEYINPUT4), .B(G146), .ZN(n735) );
  XNOR2_X2 U576 ( .A(G125), .B(KEYINPUT18), .ZN(n499) );
  NOR2_X1 U577 ( .A1(n459), .A2(n670), .ZN(n671) );
  NAND2_X1 U578 ( .A1(n600), .A2(n459), .ZN(n602) );
  NAND2_X1 U579 ( .A1(n559), .A2(n684), .ZN(n468) );
  XNOR2_X2 U580 ( .A(n534), .B(n469), .ZN(n553) );
  BUF_X1 U581 ( .A(n624), .Z(n718) );
  NOR2_X1 U582 ( .A1(n557), .A2(n558), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n553), .B(n552), .ZN(n639) );
  XNOR2_X1 U584 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n470) );
  INV_X1 U585 ( .A(n745), .ZN(n599) );
  INV_X1 U586 ( .A(G110), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U589 ( .A(KEYINPUT39), .ZN(n601) );
  XNOR2_X1 U590 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U591 ( .A(n602), .B(n601), .ZN(n617) );
  XNOR2_X1 U592 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U593 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n643) );
  INV_X1 U594 ( .A(KEYINPUT56), .ZN(n634) );
  XNOR2_X1 U595 ( .A(n644), .B(n643), .ZN(G57) );
  XNOR2_X1 U596 ( .A(KEYINPUT13), .B(G475), .ZN(n484) );
  XOR2_X2 U597 ( .A(G113), .B(G104), .Z(n495) );
  XOR2_X1 U598 ( .A(n495), .B(n533), .Z(n472) );
  NOR2_X1 U599 ( .A1(G953), .A2(G237), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G214), .A2(n548), .ZN(n471) );
  XNOR2_X1 U601 ( .A(n472), .B(n471), .ZN(n476) );
  XOR2_X1 U602 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n474) );
  XNOR2_X1 U603 ( .A(KEYINPUT104), .B(KEYINPUT12), .ZN(n473) );
  XNOR2_X1 U604 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U605 ( .A(n476), .B(n475), .Z(n482) );
  XOR2_X1 U606 ( .A(G125), .B(KEYINPUT10), .Z(n477) );
  XNOR2_X1 U607 ( .A(G140), .B(n477), .ZN(n734) );
  XNOR2_X1 U608 ( .A(G146), .B(n734), .ZN(n527) );
  XOR2_X1 U609 ( .A(KEYINPUT105), .B(KEYINPUT102), .Z(n479) );
  XNOR2_X1 U610 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U611 ( .A(n527), .B(n480), .ZN(n481) );
  XNOR2_X1 U612 ( .A(n482), .B(n481), .ZN(n645) );
  NOR2_X1 U613 ( .A1(G902), .A2(n645), .ZN(n483) );
  XNOR2_X1 U614 ( .A(n484), .B(n483), .ZN(n572) );
  INV_X1 U615 ( .A(n572), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n518), .A2(G217), .ZN(n491) );
  XOR2_X2 U617 ( .A(G122), .B(G107), .Z(n494) );
  XOR2_X1 U618 ( .A(KEYINPUT7), .B(n494), .Z(n489) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(KEYINPUT106), .Z(n490) );
  NOR2_X1 U620 ( .A1(G902), .A2(n712), .ZN(n492) );
  XNOR2_X1 U621 ( .A(G478), .B(n492), .ZN(n571) );
  INV_X1 U622 ( .A(n672), .ZN(n517) );
  XOR2_X1 U623 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n496) );
  INV_X1 U624 ( .A(n540), .ZN(n498) );
  XOR2_X1 U625 ( .A(KEYINPUT17), .B(KEYINPUT79), .Z(n500) );
  XNOR2_X1 U626 ( .A(n501), .B(KEYINPUT90), .ZN(n502) );
  NAND2_X1 U627 ( .A1(n629), .A2(n621), .ZN(n504) );
  OR2_X1 U628 ( .A1(G237), .A2(G902), .ZN(n505) );
  NAND2_X1 U629 ( .A1(n505), .A2(G210), .ZN(n503) );
  NAND2_X1 U630 ( .A1(G214), .A2(n505), .ZN(n670) );
  NAND2_X1 U631 ( .A1(G234), .A2(G237), .ZN(n506) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n506), .ZN(n509) );
  NAND2_X1 U633 ( .A1(G902), .A2(n509), .ZN(n579) );
  INV_X1 U634 ( .A(n579), .ZN(n507) );
  NAND2_X1 U635 ( .A1(n729), .A2(n507), .ZN(n508) );
  XNOR2_X1 U636 ( .A(n508), .B(KEYINPUT94), .ZN(n511) );
  NAND2_X1 U637 ( .A1(G952), .A2(n509), .ZN(n696) );
  NOR2_X1 U638 ( .A1(n696), .A2(G953), .ZN(n510) );
  XNOR2_X1 U639 ( .A(n510), .B(KEYINPUT93), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n511), .A2(n582), .ZN(n512) );
  XNOR2_X2 U641 ( .A(n513), .B(KEYINPUT0), .ZN(n557) );
  NAND2_X1 U642 ( .A1(G234), .A2(n621), .ZN(n514) );
  XNOR2_X1 U643 ( .A(KEYINPUT20), .B(n514), .ZN(n529) );
  NAND2_X1 U644 ( .A1(G221), .A2(n529), .ZN(n515) );
  XNOR2_X1 U645 ( .A(KEYINPUT21), .B(n515), .ZN(n681) );
  XOR2_X1 U646 ( .A(KEYINPUT99), .B(n681), .Z(n558) );
  NAND2_X1 U647 ( .A1(n518), .A2(G221), .ZN(n526) );
  XOR2_X1 U648 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n520) );
  XNOR2_X1 U649 ( .A(G128), .B(KEYINPUT24), .ZN(n519) );
  XNOR2_X1 U650 ( .A(n520), .B(n519), .ZN(n524) );
  XNOR2_X1 U651 ( .A(n526), .B(n525), .ZN(n528) );
  XNOR2_X1 U652 ( .A(n528), .B(n527), .ZN(n714) );
  NAND2_X1 U653 ( .A1(n529), .A2(G217), .ZN(n531) );
  XNOR2_X1 U654 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n530) );
  XNOR2_X1 U655 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U656 ( .A(G140), .B(n538), .ZN(n542) );
  XNOR2_X1 U657 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U658 ( .A(n542), .B(n541), .ZN(n544) );
  XNOR2_X2 U659 ( .A(n547), .B(n546), .ZN(n588) );
  INV_X1 U660 ( .A(n559), .ZN(n585) );
  XOR2_X1 U661 ( .A(G113), .B(KEYINPUT5), .Z(n550) );
  NAND2_X1 U662 ( .A1(n548), .A2(G210), .ZN(n549) );
  XNOR2_X1 U663 ( .A(n550), .B(n549), .ZN(n551) );
  INV_X1 U664 ( .A(KEYINPUT44), .ZN(n555) );
  XNOR2_X1 U665 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n560) );
  XNOR2_X1 U666 ( .A(KEYINPUT34), .B(KEYINPUT80), .ZN(n561) );
  NOR2_X1 U667 ( .A1(n562), .A2(n571), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n563), .B(KEYINPUT35), .ZN(n566) );
  NAND2_X1 U669 ( .A1(n566), .A2(KEYINPUT44), .ZN(n574) );
  NOR2_X1 U670 ( .A1(n571), .A2(n572), .ZN(n567) );
  XNOR2_X1 U671 ( .A(n567), .B(KEYINPUT107), .ZN(n656) );
  NAND2_X1 U672 ( .A1(n422), .A2(n595), .ZN(n568) );
  NAND2_X1 U673 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U674 ( .A1(n572), .A2(n571), .ZN(n659) );
  NAND2_X1 U675 ( .A1(n656), .A2(n659), .ZN(n674) );
  INV_X1 U676 ( .A(KEYINPUT87), .ZN(n575) );
  INV_X1 U677 ( .A(KEYINPUT65), .ZN(n576) );
  NOR2_X1 U678 ( .A1(G900), .A2(n579), .ZN(n580) );
  NAND2_X1 U679 ( .A1(G953), .A2(n580), .ZN(n581) );
  NOR2_X1 U680 ( .A1(n659), .A2(n587), .ZN(n583) );
  INV_X1 U681 ( .A(n586), .ZN(n590) );
  NAND2_X1 U682 ( .A1(n589), .A2(n588), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n591), .A2(n670), .ZN(n592) );
  XNOR2_X1 U684 ( .A(KEYINPUT30), .B(n592), .ZN(n593) );
  NOR2_X1 U685 ( .A1(n593), .A2(n358), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n600), .A2(n597), .ZN(n598) );
  XNOR2_X1 U687 ( .A(KEYINPUT109), .B(n598), .ZN(n745) );
  NOR2_X1 U688 ( .A1(n617), .A2(n659), .ZN(n604) );
  XNOR2_X1 U689 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n603) );
  XNOR2_X1 U690 ( .A(n604), .B(n603), .ZN(n746) );
  XOR2_X1 U691 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n605) );
  XNOR2_X1 U692 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n607) );
  XNOR2_X1 U693 ( .A(n608), .B(n470), .ZN(n609) );
  XNOR2_X1 U694 ( .A(KEYINPUT48), .B(KEYINPUT71), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n349), .A2(n611), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n670), .A2(n612), .ZN(n614) );
  XNOR2_X1 U697 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n614), .B(n613), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n669) );
  INV_X1 U700 ( .A(n669), .ZN(n619) );
  OR2_X1 U701 ( .A1(n617), .A2(n656), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n618), .B(KEYINPUT115), .ZN(n748) );
  NOR2_X1 U703 ( .A1(n619), .A2(n748), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT85), .B(n621), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n622), .A2(KEYINPUT2), .ZN(n623) );
  XOR2_X1 U706 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT89), .B(KEYINPUT82), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U709 ( .A(n629), .B(n628), .Z(n630) );
  XNOR2_X1 U710 ( .A(n631), .B(n630), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n633), .A2(n704), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n635), .B(n634), .ZN(G51) );
  AND2_X1 U713 ( .A1(n636), .A2(G472), .ZN(n637) );
  XOR2_X1 U714 ( .A(KEYINPUT116), .B(KEYINPUT62), .Z(n638) );
  NAND2_X1 U715 ( .A1(n642), .A2(n704), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n648), .A2(n704), .ZN(n650) );
  INV_X1 U718 ( .A(KEYINPUT60), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(G60) );
  XOR2_X1 U720 ( .A(G101), .B(n651), .Z(G3) );
  XOR2_X1 U721 ( .A(n652), .B(G104), .Z(G6) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT26), .ZN(n654) );
  XNOR2_X1 U723 ( .A(G107), .B(n654), .ZN(G9) );
  XOR2_X1 U724 ( .A(n655), .B(G110), .Z(G12) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .Z(n658) );
  NAND2_X1 U726 ( .A1(n660), .A2(n416), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(G30) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n662) );
  NAND2_X1 U729 ( .A1(n660), .A2(n409), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(G146), .B(n663), .ZN(G48) );
  NAND2_X1 U732 ( .A1(n409), .A2(n350), .ZN(n664) );
  XNOR2_X1 U733 ( .A(G113), .B(n664), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n350), .A2(n416), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(G116), .ZN(G18) );
  XNOR2_X1 U736 ( .A(G125), .B(n667), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n668), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U738 ( .A(G140), .B(n669), .ZN(G42) );
  NOR2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT121), .B(n673), .Z(n678) );
  INV_X1 U741 ( .A(n674), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U744 ( .A(n679), .B(KEYINPUT122), .ZN(n680) );
  AND2_X1 U745 ( .A1(n373), .A2(n681), .ZN(n682) );
  XNOR2_X1 U746 ( .A(n682), .B(KEYINPUT49), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n348), .A2(n683), .ZN(n687) );
  NOR2_X1 U748 ( .A1(n684), .A2(n349), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U752 ( .A(KEYINPUT51), .B(n690), .Z(n691) );
  NOR2_X1 U753 ( .A1(n697), .A2(n691), .ZN(n692) );
  XNOR2_X1 U754 ( .A(n692), .B(KEYINPUT120), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n361), .A2(n693), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n694), .B(KEYINPUT52), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n699) );
  XOR2_X1 U758 ( .A(KEYINPUT123), .B(n360), .Z(n698) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n702), .A2(G953), .ZN(n703) );
  XNOR2_X1 U762 ( .A(n703), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U763 ( .A(n704), .ZN(n717) );
  XNOR2_X1 U764 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n707) );
  XNOR2_X1 U765 ( .A(n705), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n707), .B(n706), .ZN(n709) );
  XOR2_X1 U767 ( .A(n709), .B(n708), .Z(n710) );
  NOR2_X1 U768 ( .A1(n717), .A2(n710), .ZN(G54) );
  XNOR2_X1 U769 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n717), .A2(n713), .ZN(G63) );
  XNOR2_X1 U771 ( .A(n714), .B(n715), .ZN(n716) );
  NOR2_X1 U772 ( .A1(n717), .A2(n716), .ZN(G66) );
  OR2_X1 U773 ( .A1(G953), .A2(n718), .ZN(n722) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U776 ( .A1(n720), .A2(G898), .ZN(n721) );
  NAND2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U778 ( .A(n723), .B(KEYINPUT125), .ZN(n731) );
  XOR2_X1 U779 ( .A(G110), .B(n724), .Z(n727) );
  XNOR2_X1 U780 ( .A(G101), .B(n725), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U783 ( .A(n731), .B(n730), .Z(G69) );
  XOR2_X1 U784 ( .A(n732), .B(KEYINPUT126), .Z(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(n738) );
  XOR2_X1 U787 ( .A(n738), .B(n625), .Z(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(G227), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n739), .B(KEYINPUT127), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n741), .A2(G953), .ZN(n742) );
  NAND2_X1 U792 ( .A1(n743), .A2(n742), .ZN(G72) );
  XOR2_X1 U793 ( .A(n744), .B(G137), .Z(G39) );
  XOR2_X1 U794 ( .A(G143), .B(n745), .Z(G45) );
  XOR2_X1 U795 ( .A(n746), .B(G131), .Z(G33) );
  XOR2_X1 U796 ( .A(G122), .B(n747), .Z(G24) );
  XNOR2_X1 U797 ( .A(G134), .B(n748), .ZN(n749) );
  XNOR2_X1 U798 ( .A(n749), .B(KEYINPUT119), .ZN(G36) );
  BUF_X1 U799 ( .A(n750), .Z(n751) );
  XOR2_X1 U800 ( .A(G119), .B(n751), .Z(G21) );
endmodule

