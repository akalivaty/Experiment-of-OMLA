//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n463), .B2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G137), .A3(new_n466), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n466), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND2_X1   g066(.A1(KEYINPUT69), .A2(G138), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n466), .B(new_n492), .C1(new_n481), .C2(new_n482), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n470), .A2(KEYINPUT4), .A3(new_n466), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n470), .A2(G126), .A3(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G50), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n505), .B2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n512), .B2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n512), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT71), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n516), .A2(new_n529), .A3(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n533), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n528), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n513), .A2(new_n514), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n537), .A2(G89), .A3(new_n524), .A4(new_n516), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT73), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n505), .A2(new_n529), .B1(new_n532), .B2(new_n534), .ZN(new_n540));
  AND4_X1   g115(.A1(KEYINPUT73), .A2(new_n540), .A3(new_n538), .A4(new_n528), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  OAI211_X1 g118(.A(G64), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n537), .A2(G90), .A3(new_n524), .A4(new_n516), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n505), .A2(G52), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AOI22_X1  g127(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n519), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n505), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n517), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(new_n504), .ZN(new_n564));
  NOR2_X1   g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  OAI211_X1 g140(.A(G53), .B(G543), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n537), .A2(G91), .A3(new_n524), .A4(new_n516), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n515), .A2(new_n574), .A3(G91), .A4(new_n516), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n570), .A2(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(G65), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n577), .A2(KEYINPUT76), .A3(new_n578), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(G651), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n583), .ZN(G299));
  NAND2_X1  g159(.A1(new_n520), .A2(new_n521), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(new_n517), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G88), .ZN(new_n588));
  INV_X1    g163(.A(new_n509), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(new_n507), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(G303));
  OAI21_X1  g166(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n515), .A2(G87), .A3(new_n516), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n505), .A2(G49), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(new_n515), .A2(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n519), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n515), .A2(G86), .A3(new_n516), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n505), .A2(G48), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n587), .A2(G85), .B1(G47), .B2(new_n505), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n519), .B2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n515), .A2(G66), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n516), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n505), .A2(KEYINPUT77), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n610), .A2(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n517), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .A4(new_n516), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n607), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n607), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(G286), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G299), .B(KEYINPUT78), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G297));
  AOI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n623), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(new_n558), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n622), .A2(G559), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n634), .B1(new_n636), .B2(G868), .ZN(G323));
  XOR2_X1   g212(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n638));
  XNOR2_X1  g213(.A(G323), .B(new_n638), .ZN(G282));
  NAND2_X1  g214(.A1(new_n468), .A2(new_n470), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n484), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n486), .A2(G123), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n466), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n644), .A2(new_n645), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  INV_X1    g233(.A(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g240(.A(KEYINPUT82), .B(KEYINPUT14), .C1(new_n660), .C2(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XOR2_X1   g244(.A(G2443), .B(G2446), .Z(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n667), .B2(new_n668), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n657), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n656), .A3(new_n673), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n655), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G14), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n676), .A2(new_n678), .A3(new_n655), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT83), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT83), .ZN(new_n685));
  NAND4_X1  g260(.A1(new_n676), .A2(new_n678), .A3(new_n685), .A4(new_n655), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n681), .A2(KEYINPUT85), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(KEYINPUT85), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G401));
  INV_X1    g265(.A(KEYINPUT18), .ZN(new_n691));
  XOR2_X1   g266(.A(G2084), .B(G2090), .Z(new_n692));
  XNOR2_X1  g267(.A(G2067), .B(G2678), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT17), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT86), .B(G2100), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G2072), .B(G2078), .Z(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n694), .B2(KEYINPUT18), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(new_n651), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(G227));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1956), .B(G2474), .Z(new_n706));
  XOR2_X1   g281(.A(G1961), .B(G1966), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT87), .ZN(new_n709));
  XOR2_X1   g284(.A(G1971), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT19), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(KEYINPUT87), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n706), .A2(new_n707), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(new_n708), .ZN(new_n718));
  MUX2_X1   g293(.A(new_n718), .B(new_n717), .S(new_n711), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT89), .Z(new_n721));
  AND3_X1   g296(.A1(new_n715), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n715), .B2(new_n719), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(G1991), .B(G1996), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n724), .A2(new_n726), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n705), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n729), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n731), .A2(new_n704), .A3(new_n727), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(G229));
  XOR2_X1   g308(.A(KEYINPUT93), .B(G16), .Z(new_n734));
  MUX2_X1   g309(.A(G303), .B(G22), .S(new_n734), .Z(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G6), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n602), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT32), .B(G1981), .ZN(new_n740));
  MUX2_X1   g315(.A(G23), .B(G288), .S(G16), .Z(new_n741));
  XOR2_X1   g316(.A(KEYINPUT33), .B(G1976), .Z(new_n742));
  AOI22_X1  g317(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n739), .A2(new_n740), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n737), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT34), .ZN(new_n747));
  OR2_X1    g322(.A1(G25), .A2(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n484), .A2(G131), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n486), .A2(G119), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n466), .A2(G107), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT90), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n748), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT35), .B(G1991), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT92), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n746), .A2(KEYINPUT34), .ZN(new_n762));
  MUX2_X1   g337(.A(G290), .B(G24), .S(new_n734), .Z(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1986), .Z(new_n764));
  NAND4_X1  g339(.A1(new_n747), .A2(new_n761), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT36), .ZN(new_n766));
  MUX2_X1   g341(.A(G5), .B(G301), .S(G16), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G1961), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT101), .Z(new_n769));
  MUX2_X1   g344(.A(G21), .B(G286), .S(G16), .Z(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(G1966), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n770), .A2(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT99), .B(KEYINPUT31), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G11), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT100), .ZN(new_n777));
  AOI21_X1  g352(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n650), .B2(new_n757), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(KEYINPUT102), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n757), .A2(G26), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT28), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n484), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n486), .A2(G128), .ZN(new_n786));
  INV_X1    g361(.A(G104), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n787), .A2(new_n466), .A3(KEYINPUT96), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT96), .B1(new_n787), .B2(new_n466), .ZN(new_n789));
  OAI221_X1 g364(.A(G2104), .B1(G116), .B2(new_n466), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n785), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT97), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(KEYINPUT97), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n784), .B1(new_n794), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n623), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G4), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT94), .B(G1348), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n797), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n633), .B(G19), .S(new_n734), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT95), .B(G1341), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G1961), .B2(new_n767), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G141), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n486), .A2(G129), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n468), .A2(G105), .ZN(new_n810));
  NAND3_X1  g385(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT26), .Z(new_n812));
  NAND4_X1  g387(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n757), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n757), .B2(G32), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT27), .B(G1996), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2084), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT24), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(G34), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(G34), .ZN(new_n822));
  AOI21_X1  g397(.A(G29), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n479), .B2(G29), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n757), .A2(G33), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT25), .Z(new_n828));
  AOI22_X1  g403(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n829));
  INV_X1    g404(.A(new_n484), .ZN(new_n830));
  INV_X1    g405(.A(G139), .ZN(new_n831));
  OAI221_X1 g406(.A(new_n828), .B1(new_n829), .B2(new_n466), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n826), .B1(new_n833), .B2(new_n757), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(G2072), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n824), .A2(new_n819), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n818), .A2(new_n825), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(G2072), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n757), .A2(G35), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G162), .B2(new_n757), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT29), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n839), .B1(G2090), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n807), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n757), .A2(G27), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G164), .B2(new_n757), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G2078), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n782), .A2(new_n803), .A3(new_n844), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(G2090), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT104), .B(G1956), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n734), .A2(G20), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT23), .Z(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G299), .B2(G16), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n850), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n851), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(KEYINPUT105), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(KEYINPUT105), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n781), .B2(KEYINPUT102), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n849), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n766), .A2(new_n860), .ZN(G150));
  INV_X1    g436(.A(G150), .ZN(G311));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n515), .B2(G67), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n866));
  OAI21_X1  g441(.A(G651), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g442(.A(KEYINPUT106), .B(new_n864), .C1(new_n515), .C2(G67), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n537), .A2(G93), .A3(new_n524), .A4(new_n516), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n505), .A2(G55), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n869), .A2(KEYINPUT107), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT107), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  OAI22_X1  g447(.A1(new_n867), .A2(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n537), .A2(G67), .A3(new_n524), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n863), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT106), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n865), .A2(new_n866), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(G651), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n869), .A2(new_n870), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n869), .A2(KEYINPUT107), .A3(new_n870), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n885), .A3(KEYINPUT108), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n875), .A2(new_n633), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n873), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(KEYINPUT108), .A3(new_n558), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n623), .A2(G559), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n894));
  AOI21_X1  g469(.A(G860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n873), .A2(G860), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT37), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G145));
  NAND3_X1  g474(.A1(new_n792), .A2(G164), .A3(new_n793), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G164), .B1(new_n792), .B2(new_n793), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n833), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n832), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n813), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n814), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n484), .A2(G142), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n486), .A2(G130), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n466), .A2(G118), .ZN(new_n912));
  OAI21_X1  g487(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n641), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n754), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n909), .B1(KEYINPUT109), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n479), .B(new_n650), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G162), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n907), .A2(new_n922), .A3(new_n908), .A4(new_n916), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n909), .A2(new_n916), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n907), .A2(new_n908), .A3(new_n917), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n920), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g505(.A(G290), .B(G166), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n602), .B(G288), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n636), .B(new_n890), .ZN(new_n941));
  NOR2_X1   g516(.A1(G299), .A2(new_n622), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n583), .A2(new_n576), .B1(new_n616), .B2(new_n621), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n942), .B2(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(G299), .A2(new_n622), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n576), .A2(new_n583), .A3(new_n616), .A4(new_n621), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(KEYINPUT41), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n940), .A2(new_n945), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n940), .B1(new_n945), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G868), .B2(new_n888), .ZN(G295));
  OAI21_X1  g531(.A(new_n955), .B1(G868), .B2(new_n888), .ZN(G331));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT41), .B1(new_n948), .B2(new_n949), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n547), .A2(new_n550), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n519), .B1(new_n544), .B2(new_n545), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n548), .A2(new_n549), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT112), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n963), .B(new_n966), .C1(new_n539), .C2(new_n541), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT73), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n540), .A2(new_n528), .ZN(new_n969));
  INV_X1    g544(.A(new_n538), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n536), .A2(KEYINPUT73), .A3(new_n538), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(G301), .A3(new_n972), .A4(KEYINPUT112), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n974), .A2(new_n889), .A3(new_n887), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n887), .A2(new_n889), .B1(new_n973), .B2(new_n967), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n961), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n977), .A2(KEYINPUT113), .B1(new_n978), .B2(new_n944), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(new_n973), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n890), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n974), .A2(new_n887), .A3(new_n889), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n951), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n933), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n944), .A3(new_n982), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n977), .A2(new_n933), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n928), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n958), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n987), .B1(new_n983), .B2(new_n984), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n977), .A2(KEYINPUT113), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n934), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n988), .A2(new_n928), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT115), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n990), .A2(KEYINPUT43), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(new_n944), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n975), .A2(new_n976), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n934), .B1(new_n1001), .B2(new_n983), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n994), .A2(new_n998), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(new_n999), .A3(new_n928), .A4(new_n988), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT114), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n997), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n996), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n993), .A2(new_n994), .A3(new_n999), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1002), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT43), .B1(new_n1009), .B2(new_n989), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(G397));
  NAND4_X1  g589(.A1(new_n478), .A2(G40), .A3(new_n469), .A4(new_n471), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n472), .A2(KEYINPUT116), .A3(G40), .A4(new_n478), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n500), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n794), .B(G2067), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n813), .B(G1996), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1023), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n754), .B(new_n760), .Z(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G290), .B(G1986), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n500), .A2(new_n1020), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n592), .A2(new_n593), .A3(G1976), .A4(new_n594), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1033), .B(G8), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT119), .ZN(new_n1040));
  INV_X1    g615(.A(new_n598), .ZN(new_n1041));
  INV_X1    g616(.A(new_n601), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G1981), .B1(new_n598), .B2(new_n601), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1033), .A2(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT120), .A4(KEYINPUT49), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1049), .B(new_n1056), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1038), .A2(new_n1058), .A3(KEYINPUT52), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1040), .A2(new_n1054), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1032), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n500), .A2(new_n1020), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT50), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n500), .A2(new_n1063), .A3(new_n1020), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1019), .A2(new_n1021), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n1069), .A2(G2090), .B1(new_n1071), .B2(G1971), .ZN(new_n1072));
  NAND3_X1  g647(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G288), .A2(G1976), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1054), .A2(new_n1078), .B1(new_n1043), .B2(new_n602), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1049), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1060), .A2(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1072), .A2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1038), .A2(new_n1058), .A3(KEYINPUT52), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1058), .B1(new_n1038), .B2(KEYINPUT52), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(KEYINPUT121), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1076), .B1(new_n1072), .B2(G8), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1060), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1022), .A2(new_n1017), .A3(new_n1018), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1966), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1069), .B2(G2084), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1082), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1076), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1089), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1066), .A2(new_n1017), .A3(new_n1018), .A4(new_n1067), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G2090), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1104), .A2(new_n1105), .B1(new_n1094), .B2(new_n736), .ZN(new_n1106));
  INV_X1    g681(.A(G8), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1083), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1085), .A2(new_n1088), .A3(new_n1077), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1097), .A2(G8), .A3(G168), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1102), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1081), .B1(new_n1101), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1071), .A2(new_n1113), .B1(new_n1114), .B2(new_n1103), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n576), .A2(new_n583), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1103), .A2(new_n1114), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1070), .A2(new_n1021), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(new_n1061), .A3(new_n1113), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1122), .A2(new_n1124), .B1(new_n1118), .B2(new_n1116), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1068), .A2(new_n1066), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1064), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1061), .A2(new_n796), .A3(new_n1032), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n622), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1128), .A2(new_n1134), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1121), .A2(new_n1138), .A3(new_n1127), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1132), .A2(new_n622), .A3(new_n1133), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1134), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1135), .A2(new_n1119), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1137), .B1(new_n1143), .B2(new_n1125), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT123), .B(G1996), .Z(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1123), .A2(new_n1061), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1033), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g725(.A(new_n1145), .B(new_n633), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1094), .B2(new_n1146), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT59), .B1(new_n1152), .B2(new_n558), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n622), .A2(KEYINPUT60), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1132), .A2(new_n1133), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1144), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1136), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1097), .A2(G8), .A3(G286), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT124), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1096), .B(G168), .C1(new_n1069), .C2(G2084), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G8), .ZN(new_n1162));
  NOR2_X1   g737(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1161), .B(G8), .C1(KEYINPUT125), .C2(KEYINPUT51), .ZN(new_n1165));
  NAND2_X1  g740(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1160), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1109), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1060), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1172), .A2(KEYINPUT126), .A3(new_n1077), .A4(new_n1108), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n1174));
  INV_X1    g749(.A(G2078), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1071), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT53), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G1961), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1069), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1015), .A2(new_n1177), .A3(G2078), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1123), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1178), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1174), .B1(new_n1183), .B2(G171), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1176), .A2(new_n1177), .B1(new_n1069), .B2(new_n1179), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n1175), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1185), .A2(new_n1186), .A3(G301), .A4(new_n1187), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1178), .A2(G301), .A3(new_n1180), .A4(new_n1187), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1184), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1183), .A2(G171), .ZN(new_n1192));
  AOI21_X1  g767(.A(G301), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1174), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1171), .A2(new_n1173), .A3(new_n1191), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1112), .B1(new_n1169), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1171), .A2(new_n1173), .A3(new_n1193), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1168), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1160), .A2(new_n1167), .A3(KEYINPUT62), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1031), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1023), .B1(new_n1024), .B2(new_n813), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1027), .A2(G1996), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1204), .A2(KEYINPUT46), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1204), .A2(KEYINPUT46), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1203), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g782(.A(new_n1207), .B(KEYINPUT47), .Z(new_n1208));
  NOR3_X1   g783(.A1(new_n1027), .A2(G1986), .A3(G290), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT48), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n794), .A2(G2067), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n756), .A2(new_n760), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1211), .B1(new_n1026), .B2(new_n1212), .ZN(new_n1213));
  OAI22_X1  g788(.A1(new_n1029), .A2(new_n1210), .B1(new_n1213), .B2(new_n1027), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1208), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1202), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g791(.A1(G227), .A2(new_n461), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G229), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g793(.A(new_n929), .B(new_n1219), .C1(new_n688), .C2(new_n689), .ZN(new_n1220));
  INV_X1    g794(.A(new_n1011), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1220), .A2(new_n1221), .ZN(G308));
  OR2_X1    g796(.A1(new_n1220), .A2(new_n1221), .ZN(G225));
endmodule


