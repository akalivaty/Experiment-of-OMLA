

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U548 ( .A1(n533), .A2(n532), .ZN(G160) );
  INV_X1 U549 ( .A(n751), .ZN(n730) );
  NAND2_X1 U550 ( .A1(n700), .A2(G8), .ZN(n701) );
  XOR2_X1 U551 ( .A(n736), .B(KEYINPUT28), .Z(n513) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(KEYINPUT30), .ZN(n514) );
  INV_X1 U553 ( .A(KEYINPUT99), .ZN(n727) );
  XNOR2_X1 U554 ( .A(n701), .B(n514), .ZN(n702) );
  XNOR2_X1 U555 ( .A(n758), .B(KEYINPUT32), .ZN(n759) );
  NAND2_X1 U556 ( .A1(n697), .A2(n696), .ZN(n751) );
  NOR2_X1 U557 ( .A1(n630), .A2(G651), .ZN(n648) );
  NOR2_X1 U558 ( .A1(n525), .A2(n524), .ZN(G164) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n515), .Z(n873) );
  NAND2_X1 U561 ( .A1(G138), .A2(n873), .ZN(n516) );
  XNOR2_X1 U562 ( .A(n516), .B(KEYINPUT92), .ZN(n519) );
  INV_X1 U563 ( .A(G2105), .ZN(n520) );
  XOR2_X1 U564 ( .A(KEYINPUT65), .B(G2104), .Z(n521) );
  AND2_X1 U565 ( .A1(n520), .A2(n521), .ZN(n871) );
  NAND2_X1 U566 ( .A1(G102), .A2(n871), .ZN(n517) );
  XOR2_X1 U567 ( .A(KEYINPUT91), .B(n517), .Z(n518) );
  NAND2_X1 U568 ( .A1(n519), .A2(n518), .ZN(n525) );
  AND2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n867) );
  NAND2_X1 U570 ( .A1(G114), .A2(n867), .ZN(n523) );
  NOR2_X2 U571 ( .A1(n521), .A2(n520), .ZN(n868) );
  NAND2_X1 U572 ( .A1(G126), .A2(n868), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G125), .A2(n868), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n526), .B(KEYINPUT66), .ZN(n529) );
  NAND2_X1 U576 ( .A1(G101), .A2(n871), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(n527), .Z(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U579 ( .A1(G113), .A2(n867), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G137), .A2(n873), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U582 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U583 ( .A1(G123), .A2(n868), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n534), .B(KEYINPUT18), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT80), .ZN(n537) );
  NAND2_X1 U586 ( .A1(G135), .A2(n873), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U588 ( .A(KEYINPUT81), .B(n538), .ZN(n543) );
  NAND2_X1 U589 ( .A1(G111), .A2(n867), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G99), .A2(n871), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U592 ( .A(KEYINPUT82), .B(n541), .Z(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n992) );
  XNOR2_X1 U594 ( .A(G2096), .B(n992), .ZN(n544) );
  OR2_X1 U595 ( .A1(G2100), .A2(n544), .ZN(G156) );
  INV_X1 U596 ( .A(G57), .ZN(G237) );
  INV_X1 U597 ( .A(G108), .ZN(G238) );
  INV_X1 U598 ( .A(G69), .ZN(G235) );
  NAND2_X1 U599 ( .A1(G7), .A2(G661), .ZN(n545) );
  XNOR2_X1 U600 ( .A(n545), .B(KEYINPUT72), .ZN(n546) );
  XNOR2_X1 U601 ( .A(KEYINPUT10), .B(n546), .ZN(G223) );
  INV_X1 U602 ( .A(G223), .ZN(n820) );
  NAND2_X1 U603 ( .A1(n820), .A2(G567), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT11), .B(n547), .Z(G234) );
  INV_X1 U605 ( .A(G651), .ZN(n552) );
  NOR2_X1 U606 ( .A1(G543), .A2(n552), .ZN(n549) );
  XNOR2_X1 U607 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n548) );
  XNOR2_X2 U608 ( .A(n549), .B(n548), .ZN(n641) );
  NAND2_X1 U609 ( .A1(n641), .A2(G56), .ZN(n550) );
  XNOR2_X1 U610 ( .A(KEYINPUT14), .B(n550), .ZN(n557) );
  NOR2_X1 U611 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U612 ( .A1(n642), .A2(G81), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n551), .B(KEYINPUT12), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT0), .B(G543), .Z(n630) );
  NOR2_X1 U615 ( .A1(n630), .A2(n552), .ZN(n643) );
  NAND2_X1 U616 ( .A1(G68), .A2(n643), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U618 ( .A(KEYINPUT13), .B(n555), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT73), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n648), .A2(G43), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n971) );
  INV_X1 U623 ( .A(G860), .ZN(n603) );
  OR2_X1 U624 ( .A1(n971), .A2(n603), .ZN(G153) );
  NAND2_X1 U625 ( .A1(n642), .A2(G90), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT70), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G77), .A2(n643), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT9), .B(n564), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n648), .A2(G52), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT68), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G64), .A2(n641), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT69), .B(n568), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G92), .A2(n642), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G79), .A2(n643), .ZN(n571) );
  AND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n641), .A2(G66), .ZN(n573) );
  XOR2_X1 U640 ( .A(n573), .B(KEYINPUT74), .Z(n575) );
  AND2_X1 U641 ( .A1(n648), .A2(G54), .ZN(n574) );
  NOR2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X2 U644 ( .A(n578), .B(KEYINPUT15), .Z(n955) );
  INV_X1 U645 ( .A(n955), .ZN(n611) );
  NOR2_X1 U646 ( .A1(n611), .A2(G868), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT75), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U650 ( .A1(n642), .A2(G89), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G76), .A2(n643), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n585) );
  XNOR2_X1 U655 ( .A(KEYINPUT5), .B(n585), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n587), .B(n586), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G63), .A2(n641), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G51), .A2(n648), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U660 ( .A(KEYINPUT6), .B(n590), .Z(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT7), .B(n593), .ZN(G168) );
  XOR2_X1 U663 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U664 ( .A1(G65), .A2(n641), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G91), .A2(n642), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G78), .A2(n643), .ZN(n596) );
  XNOR2_X1 U668 ( .A(KEYINPUT71), .B(n596), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n648), .A2(G53), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(G299) );
  INV_X1 U672 ( .A(G868), .ZN(n651) );
  NOR2_X1 U673 ( .A1(G286), .A2(n651), .ZN(n602) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n604), .A2(n611), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U679 ( .A1(n611), .A2(G868), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G559), .A2(n606), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT79), .B(n607), .Z(n610) );
  NOR2_X1 U682 ( .A1(G868), .A2(n971), .ZN(n608) );
  XNOR2_X1 U683 ( .A(KEYINPUT78), .B(n608), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U685 ( .A1(n611), .A2(G559), .ZN(n661) );
  XNOR2_X1 U686 ( .A(n971), .B(n661), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n612), .A2(G860), .ZN(n619) );
  NAND2_X1 U688 ( .A1(G67), .A2(n641), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G93), .A2(n642), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G80), .A2(n643), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G55), .A2(n648), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n658) );
  XOR2_X1 U695 ( .A(n619), .B(n658), .Z(G145) );
  NAND2_X1 U696 ( .A1(G61), .A2(n641), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G86), .A2(n642), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n643), .A2(G73), .ZN(n622) );
  XOR2_X1 U700 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n648), .A2(G48), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U704 ( .A1(G49), .A2(n648), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n641), .A2(n629), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G88), .A2(n642), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G75), .A2(n643), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U713 ( .A(KEYINPUT84), .B(n635), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G62), .A2(n641), .ZN(n636) );
  XNOR2_X1 U715 ( .A(KEYINPUT83), .B(n636), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n648), .A2(G50), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  AND2_X1 U720 ( .A1(n641), .A2(G60), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G85), .A2(n642), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G72), .A2(n643), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n648), .A2(G47), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U727 ( .A1(n651), .A2(n658), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(KEYINPUT86), .ZN(n664) );
  XOR2_X1 U729 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n653) );
  XNOR2_X1 U730 ( .A(G288), .B(n653), .ZN(n654) );
  XNOR2_X1 U731 ( .A(G305), .B(n654), .ZN(n656) );
  INV_X1 U732 ( .A(G299), .ZN(n961) );
  XNOR2_X1 U733 ( .A(n961), .B(G166), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U735 ( .A(n658), .B(n657), .Z(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(G290), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n971), .B(n660), .ZN(n885) );
  XNOR2_X1 U738 ( .A(n885), .B(n661), .ZN(n662) );
  NAND2_X1 U739 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n670) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U750 ( .A1(n671), .A2(G218), .ZN(n672) );
  NAND2_X1 U751 ( .A1(G96), .A2(n672), .ZN(n824) );
  NAND2_X1 U752 ( .A1(G2106), .A2(n824), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT88), .B(n673), .Z(n679) );
  NOR2_X1 U754 ( .A1(G235), .A2(G238), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G120), .A2(n674), .ZN(n675) );
  NOR2_X1 U756 ( .A1(n675), .A2(G237), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(KEYINPUT89), .ZN(n825) );
  NAND2_X1 U758 ( .A1(G567), .A2(n825), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT90), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(n679), .A2(n678), .ZN(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U763 ( .A1(n681), .A2(n680), .ZN(n823) );
  NAND2_X1 U764 ( .A1(n823), .A2(G36), .ZN(G176) );
  XNOR2_X1 U765 ( .A(G2067), .B(KEYINPUT37), .ZN(n813) );
  NAND2_X1 U766 ( .A1(n867), .A2(G116), .ZN(n682) );
  XNOR2_X1 U767 ( .A(n682), .B(KEYINPUT94), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G128), .A2(n868), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT35), .ZN(n690) );
  NAND2_X1 U771 ( .A1(n871), .A2(G104), .ZN(n687) );
  NAND2_X1 U772 ( .A1(n873), .A2(G140), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT34), .B(n688), .Z(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U776 ( .A(n691), .B(KEYINPUT36), .Z(n881) );
  OR2_X1 U777 ( .A1(n813), .A2(n881), .ZN(n692) );
  XNOR2_X1 U778 ( .A(n692), .B(KEYINPUT95), .ZN(n1006) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n697) );
  NAND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n695) );
  NOR2_X1 U781 ( .A1(n697), .A2(n695), .ZN(n816) );
  NAND2_X1 U782 ( .A1(n1006), .A2(n816), .ZN(n811) );
  XNOR2_X1 U783 ( .A(G1986), .B(G290), .ZN(n960) );
  NAND2_X1 U784 ( .A1(n960), .A2(n816), .ZN(n693) );
  XOR2_X1 U785 ( .A(KEYINPUT93), .B(n693), .Z(n694) );
  NAND2_X1 U786 ( .A1(n811), .A2(n694), .ZN(n788) );
  INV_X1 U787 ( .A(n695), .ZN(n696) );
  NOR2_X1 U788 ( .A1(G2084), .A2(n751), .ZN(n698) );
  NAND2_X1 U789 ( .A1(G8), .A2(n698), .ZN(n749) );
  NAND2_X1 U790 ( .A1(G8), .A2(n751), .ZN(n783) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n783), .ZN(n747) );
  NOR2_X1 U792 ( .A1(n747), .A2(n698), .ZN(n699) );
  XOR2_X1 U793 ( .A(KEYINPUT101), .B(n699), .Z(n700) );
  NOR2_X1 U794 ( .A1(G168), .A2(n702), .ZN(n707) );
  XOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .Z(n919) );
  NOR2_X1 U796 ( .A1(n919), .A2(n751), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n730), .A2(G1961), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U799 ( .A(KEYINPUT98), .B(n705), .ZN(n739) );
  AND2_X1 U800 ( .A1(G301), .A2(n739), .ZN(n706) );
  NOR2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U802 ( .A(n708), .B(KEYINPUT31), .ZN(n744) );
  AND2_X1 U803 ( .A1(G1348), .A2(n955), .ZN(n711) );
  XNOR2_X1 U804 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n719) );
  INV_X1 U805 ( .A(G1341), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n719), .A2(n709), .ZN(n710) );
  NOR2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U808 ( .A1(n712), .A2(n730), .ZN(n713) );
  NOR2_X1 U809 ( .A1(n971), .A2(n713), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n955), .A2(G2067), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n719), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n716), .A2(n730), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n719), .ZN(n720) );
  NOR2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n751), .ZN(n723) );
  NAND2_X1 U818 ( .A1(G2067), .A2(n730), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n724), .A2(n955), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U822 ( .A(n728), .B(n727), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n730), .A2(G2072), .ZN(n729) );
  XNOR2_X1 U824 ( .A(n729), .B(KEYINPUT27), .ZN(n732) );
  INV_X1 U825 ( .A(G1956), .ZN(n927) );
  NOR2_X1 U826 ( .A1(n927), .A2(n730), .ZN(n731) );
  NOR2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n735) );
  NAND2_X1 U828 ( .A1(n735), .A2(n961), .ZN(n733) );
  NAND2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n735), .A2(n961), .ZN(n736) );
  NAND2_X1 U831 ( .A1(n737), .A2(n513), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n738), .B(KEYINPUT29), .ZN(n741) );
  NOR2_X1 U833 ( .A1(G301), .A2(n739), .ZN(n740) );
  NOR2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U835 ( .A(n742), .B(KEYINPUT100), .ZN(n743) );
  NOR2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U837 ( .A(n745), .B(KEYINPUT103), .ZN(n750) );
  XOR2_X1 U838 ( .A(n750), .B(KEYINPUT104), .Z(n746) );
  NOR2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n750), .A2(G286), .ZN(n756) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n783), .ZN(n753) );
  NOR2_X1 U843 ( .A1(G2090), .A2(n751), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U845 ( .A1(n754), .A2(G303), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n757), .A2(G8), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n777) );
  NOR2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U851 ( .A1(n766), .A2(n761), .ZN(n965) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n765) );
  AND2_X1 U853 ( .A1(n965), .A2(n765), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n777), .A2(n762), .ZN(n774) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n964) );
  INV_X1 U856 ( .A(n783), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n964), .A2(n763), .ZN(n764) );
  AND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n767), .A2(n783), .ZN(n770) );
  XNOR2_X1 U861 ( .A(G1981), .B(KEYINPUT105), .ZN(n768) );
  XNOR2_X1 U862 ( .A(n768), .B(G305), .ZN(n952) );
  INV_X1 U863 ( .A(n952), .ZN(n769) );
  OR2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n780) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n775) );
  NAND2_X1 U868 ( .A1(G8), .A2(n775), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n778), .A2(n783), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n786) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XNOR2_X1 U873 ( .A(n781), .B(KEYINPUT97), .ZN(n782) );
  XNOR2_X1 U874 ( .A(n782), .B(KEYINPUT24), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n804) );
  NAND2_X1 U878 ( .A1(G117), .A2(n867), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G141), .A2(n873), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n871), .A2(G105), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n868), .A2(G129), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n866) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n866), .ZN(n991) );
  NAND2_X1 U887 ( .A1(G131), .A2(n873), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G95), .A2(n871), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n868), .A2(G119), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT96), .B(n798), .Z(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n867), .A2(G107), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n860) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n860), .ZN(n996) );
  NAND2_X1 U896 ( .A1(n991), .A2(n996), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n816), .A2(n803), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n804), .A2(n805), .ZN(n818) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n866), .ZN(n984) );
  INV_X1 U900 ( .A(n805), .ZN(n808) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n860), .ZN(n989) );
  NOR2_X1 U903 ( .A1(n806), .A2(n989), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n984), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n881), .A2(n813), .ZN(n987) );
  NAND2_X1 U909 ( .A1(n814), .A2(n987), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n819), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U915 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(G188) );
  XNOR2_X1 U918 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U920 ( .A(G132), .ZN(G219) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G82), .ZN(G220) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XOR2_X1 U925 ( .A(G2100), .B(G2096), .Z(n827) );
  XNOR2_X1 U926 ( .A(KEYINPUT42), .B(G2678), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(G2090), .Z(n829) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U931 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2078), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(G227) );
  XNOR2_X1 U934 ( .A(G1991), .B(KEYINPUT110), .ZN(n843) );
  XOR2_X1 U935 ( .A(G1981), .B(G1956), .Z(n835) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1986), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n837) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1961), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U941 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U942 ( .A(G2474), .B(KEYINPUT41), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(G229) );
  NAND2_X1 U945 ( .A1(G112), .A2(n867), .ZN(n845) );
  NAND2_X1 U946 ( .A1(G136), .A2(n873), .ZN(n844) );
  NAND2_X1 U947 ( .A1(n845), .A2(n844), .ZN(n850) );
  NAND2_X1 U948 ( .A1(n868), .A2(G124), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U950 ( .A1(G100), .A2(n871), .ZN(n847) );
  NAND2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U952 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U953 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n859) );
  NAND2_X1 U954 ( .A1(G139), .A2(n873), .ZN(n852) );
  NAND2_X1 U955 ( .A1(G103), .A2(n871), .ZN(n851) );
  NAND2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G115), .A2(n867), .ZN(n854) );
  NAND2_X1 U958 ( .A1(G127), .A2(n868), .ZN(n853) );
  NAND2_X1 U959 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n855), .Z(n856) );
  NOR2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n1000) );
  XNOR2_X1 U962 ( .A(n1000), .B(KEYINPUT112), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n860), .B(G162), .ZN(n862) );
  XNOR2_X1 U965 ( .A(G164), .B(G160), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U967 ( .A(n864), .B(n863), .Z(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G118), .A2(n867), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G130), .A2(n868), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n871), .A2(G106), .ZN(n872) );
  XOR2_X1 U973 ( .A(KEYINPUT111), .B(n872), .Z(n875) );
  NAND2_X1 U974 ( .A1(n873), .A2(G142), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U976 ( .A(n876), .B(KEYINPUT45), .Z(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(n880), .B(n879), .Z(n883) );
  XNOR2_X1 U979 ( .A(n992), .B(n881), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  NOR2_X1 U981 ( .A1(G37), .A2(n884), .ZN(G395) );
  INV_X1 U982 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U983 ( .A(G286), .B(n955), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(G171), .ZN(n888) );
  NOR2_X1 U986 ( .A1(G37), .A2(n888), .ZN(G397) );
  XOR2_X1 U987 ( .A(KEYINPUT108), .B(G2438), .Z(n890) );
  XNOR2_X1 U988 ( .A(G2443), .B(KEYINPUT107), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U990 ( .A(G2451), .B(KEYINPUT106), .Z(n892) );
  XNOR2_X1 U991 ( .A(G2430), .B(G2454), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U994 ( .A(G2435), .B(G2446), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n899) );
  XOR2_X1 U996 ( .A(G1348), .B(G1341), .Z(n897) );
  XNOR2_X1 U997 ( .A(G2427), .B(n897), .ZN(n898) );
  XOR2_X1 U998 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U999 ( .A1(G14), .A2(n900), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(n906), .ZN(G401) );
  XOR2_X1 U1008 ( .A(G2090), .B(G35), .Z(n910) );
  XOR2_X1 U1009 ( .A(G2084), .B(G34), .Z(n907) );
  XNOR2_X1 U1010 ( .A(KEYINPUT118), .B(n907), .ZN(n908) );
  XNOR2_X1 U1011 ( .A(n908), .B(KEYINPUT54), .ZN(n909) );
  NAND2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n924) );
  XNOR2_X1 U1013 ( .A(G1996), .B(G32), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(G1991), .B(G25), .ZN(n911) );
  NOR2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n918) );
  XOR2_X1 U1016 ( .A(G2072), .B(G33), .Z(n913) );
  NAND2_X1 U1017 ( .A1(n913), .A2(G28), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT117), .B(G2067), .Z(n914) );
  XNOR2_X1 U1019 ( .A(G26), .B(n914), .ZN(n915) );
  NOR2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1021 ( .A1(n918), .A2(n917), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G27), .B(n919), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(n922), .B(KEYINPUT53), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1026 ( .A(KEYINPUT55), .B(n925), .Z(n926) );
  NOR2_X1 U1027 ( .A1(G29), .A2(n926), .ZN(n1017) );
  XOR2_X1 U1028 ( .A(KEYINPUT123), .B(G16), .Z(n951) );
  XNOR2_X1 U1029 ( .A(n927), .B(G20), .ZN(n935) );
  XOR2_X1 U1030 ( .A(G1341), .B(G19), .Z(n930) );
  XOR2_X1 U1031 ( .A(G6), .B(KEYINPUT124), .Z(n928) );
  XNOR2_X1 U1032 ( .A(G1981), .B(n928), .ZN(n929) );
  NAND2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1034 ( .A(KEYINPUT59), .B(G1348), .Z(n931) );
  XNOR2_X1 U1035 ( .A(G4), .B(n931), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(n936), .B(KEYINPUT60), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(KEYINPUT125), .B(n937), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(G5), .B(G1961), .ZN(n938) );
  NOR2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G1986), .B(G24), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n942) );
  NOR2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n945) );
  XOR2_X1 U1047 ( .A(G1976), .B(G23), .Z(n944) );
  NAND2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(n946), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1051 ( .A(KEYINPUT61), .B(n949), .Z(n950) );
  NOR2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n981) );
  XNOR2_X1 U1053 ( .A(KEYINPUT56), .B(G16), .ZN(n978) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1056 ( .A(n954), .B(KEYINPUT57), .ZN(n976) );
  XOR2_X1 U1057 ( .A(n955), .B(G1348), .Z(n958) );
  XNOR2_X1 U1058 ( .A(G1961), .B(G301), .ZN(n956) );
  XNOR2_X1 U1059 ( .A(KEYINPUT119), .B(n956), .ZN(n957) );
  NAND2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n961), .B(G1956), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(n968), .B(KEYINPUT120), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n974) );
  XOR2_X1 U1069 ( .A(G1341), .B(n971), .Z(n972) );
  XNOR2_X1 U1070 ( .A(KEYINPUT121), .B(n972), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT122), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT126), .B(n982), .ZN(n1015) );
  XOR2_X1 U1077 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT51), .B(n985), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n986), .B(KEYINPUT113), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n999) );
  INV_X1 U1082 ( .A(n989), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G160), .B(G2084), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(G2072), .B(n1000), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G164), .B(G2078), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1001), .B(KEYINPUT114), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT50), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(KEYINPUT115), .B(n1009), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1010), .Z(n1011) );
  NOR2_X1 U1098 ( .A1(KEYINPUT55), .A2(n1011), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT116), .B(n1012), .Z(n1013) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(G29), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(G11), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(n1019), .B(KEYINPUT62), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1020), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

