//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(KEYINPUT88), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(KEYINPUT88), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n214), .A2(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n217), .A2(new_n218), .B1(new_n213), .B2(new_n208), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n219), .B(new_n221), .C1(new_n211), .C2(new_n212), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT96), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(G85gat), .A3(G92gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228));
  INV_X1    g027(.A(G85gat), .ZN(new_n229));
  INV_X1    g028(.A(G92gat), .ZN(new_n230));
  AOI22_X1  g029(.A1(KEYINPUT8), .A2(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n227), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G99gat), .B(G106gat), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT89), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n243), .A3(new_n240), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n236), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n223), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n223), .B2(new_n240), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n239), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G190gat), .B(G218gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT98), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n207), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT97), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n251), .B2(new_n253), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n253), .B2(new_n251), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n251), .A2(KEYINPUT97), .A3(new_n253), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n254), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n251), .A2(new_n253), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(KEYINPUT98), .ZN(new_n265));
  INV_X1    g064(.A(new_n260), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n207), .A4(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G57gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(G64gat), .ZN(new_n270));
  INV_X1    g069(.A(G64gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G57gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT9), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G71gat), .A2(G78gat), .ZN(new_n274));
  INV_X1    g073(.A(G71gat), .ZN(new_n275));
  INV_X1    g074(.A(G78gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT93), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT93), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G71gat), .B2(G78gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n273), .A2(new_n274), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT9), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n274), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT94), .B1(new_n269), .B2(G64gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G57gat), .B2(new_n271), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n269), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT21), .ZN(new_n288));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(G127gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT16), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(G1gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(G1gat), .B2(new_n292), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G8gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(KEYINPUT21), .B2(new_n287), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n291), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G183gat), .B(G211gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT95), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n300), .B(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n304), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n235), .B(new_n287), .Z(new_n308));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT99), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n287), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n310), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G120gat), .B(G148gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT100), .ZN(new_n318));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  OR3_X1    g119(.A1(new_n313), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n313), .B2(new_n316), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n268), .A2(new_n307), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT101), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT36), .ZN(new_n327));
  AND2_X1   g126(.A1(G113gat), .A2(G120gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G113gat), .A2(G120gat), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT1), .ZN(new_n330));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G113gat), .A2(G120gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G134gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G127gat), .ZN(new_n341));
  INV_X1    g140(.A(G127gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n334), .A3(new_n338), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT69), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT68), .B1(new_n328), .B2(new_n329), .ZN(new_n350));
  AND4_X1   g149(.A1(KEYINPUT69), .A2(new_n349), .A3(new_n347), .A4(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n333), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n355), .A2(new_n356), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n357), .A2(new_n359), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G183gat), .ZN(new_n365));
  INV_X1    g164(.A(G190gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT24), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n364), .A2(new_n370), .B1(new_n355), .B2(new_n356), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n359), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n356), .ZN(new_n373));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n361), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n355), .A2(new_n356), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n372), .A2(new_n375), .A3(new_n376), .A4(new_n369), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT66), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT26), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n358), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(KEYINPUT66), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n384));
  NAND2_X1  g183(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n358), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n386), .A3(new_n374), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n365), .A2(KEYINPUT27), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G183gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n390), .A3(new_n366), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT28), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT27), .B(G183gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT28), .A3(new_n366), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n396), .A3(new_n368), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n350), .A2(new_n347), .A3(new_n344), .A4(new_n331), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT69), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n349), .A2(KEYINPUT69), .A3(new_n347), .A4(new_n350), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n332), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT70), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n354), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n352), .A2(new_n353), .A3(new_n397), .A4(new_n378), .ZN(new_n406));
  INV_X1    g205(.A(G227gat), .ZN(new_n407));
  INV_X1    g206(.A(G233gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n409), .B(KEYINPUT64), .Z(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT32), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n410), .A2(KEYINPUT34), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n405), .B2(new_n406), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n422));
  INV_X1    g221(.A(new_n409), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(KEYINPUT34), .ZN(new_n425));
  INV_X1    g224(.A(new_n417), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n411), .B(KEYINPUT32), .C1(new_n413), .C2(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n418), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n418), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n327), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n427), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n425), .A3(new_n427), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(KEYINPUT36), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G78gat), .B(G106gat), .Z(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT3), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT29), .ZN(new_n442));
  AND2_X1   g241(.A1(G211gat), .A2(G218gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT22), .ZN(new_n444));
  OR2_X1    g243(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(G204gat), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G204gat), .ZN(new_n448));
  AND2_X1   g247(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT73), .ZN(new_n453));
  NOR2_X1   g252(.A1(G211gat), .A2(G218gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n443), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G211gat), .ZN(new_n456));
  INV_X1    g255(.A(G218gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G211gat), .A2(G218gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(KEYINPUT73), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n442), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n452), .A2(new_n461), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n441), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G141gat), .B(G148gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT2), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(G155gat), .B2(G162gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G141gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G148gat), .ZN(new_n473));
  INV_X1    g272(.A(G148gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G141gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G155gat), .B(G162gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT2), .B1(new_n302), .B2(new_n206), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n479), .A3(new_n441), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n442), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT72), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n455), .A2(new_n460), .A3(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n452), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n485), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT82), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n455), .A2(new_n460), .A3(new_n484), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(new_n452), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n483), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G228gat), .A2(G233gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(KEYINPUT81), .Z(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT29), .B1(new_n486), .B2(new_n487), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n480), .B1(new_n498), .B2(KEYINPUT3), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n491), .B2(new_n483), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n440), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n439), .B1(new_n502), .B2(KEYINPUT83), .ZN(new_n503));
  INV_X1    g302(.A(new_n496), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n492), .B1(new_n491), .B2(new_n483), .ZN(new_n505));
  AND4_X1   g304(.A1(new_n492), .A2(new_n483), .A3(new_n486), .A4(new_n487), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n507), .B2(new_n481), .ZN(new_n508));
  INV_X1    g307(.A(new_n501), .ZN(new_n509));
  OAI21_X1  g308(.A(G22gat), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n494), .A2(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n440), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n510), .A2(KEYINPUT83), .A3(new_n512), .A4(new_n439), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(KEYINPUT84), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT84), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G226gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n408), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n398), .B2(new_n442), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n519), .B(new_n408), .C1(new_n378), .C2(new_n397), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n491), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n398), .A2(new_n520), .ZN(new_n524));
  INV_X1    g323(.A(new_n491), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT29), .B1(new_n378), .B2(new_n397), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n524), .B(new_n525), .C1(new_n520), .C2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G8gat), .B(G36gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT74), .ZN(new_n529));
  XNOR2_X1  g328(.A(G64gat), .B(G92gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n523), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n523), .A2(new_n527), .A3(KEYINPUT30), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n523), .A2(new_n527), .ZN(new_n536));
  INV_X1    g335(.A(new_n531), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n540));
  INV_X1    g339(.A(new_n480), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n403), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n352), .A2(new_n480), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G225gat), .A2(G233gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n352), .A2(new_n540), .A3(new_n480), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT5), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT75), .B1(new_n480), .B2(KEYINPUT3), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n480), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n352), .B(new_n482), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n541), .B(new_n333), .C1(new_n348), .C2(new_n351), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT4), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n541), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n552), .A2(new_n545), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G85gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT78), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT79), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G1gat), .B(G29gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT5), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n558), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT6), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n558), .A2(new_n568), .A3(KEYINPUT80), .A4(new_n565), .ZN(new_n573));
  INV_X1    g372(.A(new_n565), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n576), .A2(new_n545), .B1(new_n548), .B2(KEYINPUT5), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n577), .B2(new_n567), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n567), .B1(new_n557), .B2(new_n549), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(KEYINPUT6), .A3(new_n565), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n539), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n436), .B1(new_n518), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n515), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT83), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n511), .B2(new_n440), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n586), .A2(new_n439), .B1(new_n510), .B2(new_n512), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n575), .A2(new_n546), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n546), .B1(new_n544), .B2(new_n547), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n546), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n574), .B1(new_n594), .B2(KEYINPUT39), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n589), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n565), .B1(new_n590), .B2(new_n591), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n544), .A2(new_n547), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n594), .B(KEYINPUT39), .C1(new_n598), .C2(new_n546), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n599), .A3(KEYINPUT40), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n596), .A2(new_n569), .A3(new_n539), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n531), .B1(new_n536), .B2(KEYINPUT37), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT86), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n523), .A2(new_n527), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n523), .A2(new_n605), .A3(new_n527), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT86), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n609), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n603), .A2(new_n608), .A3(new_n611), .A4(new_n606), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n581), .A2(new_n612), .A3(new_n532), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT87), .B1(new_n609), .B2(KEYINPUT38), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n572), .B1(new_n580), .B2(new_n565), .ZN(new_n616));
  INV_X1    g415(.A(new_n569), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT85), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT85), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n578), .A2(new_n569), .A3(new_n619), .A4(new_n572), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n602), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623));
  AND4_X1   g422(.A1(new_n515), .A2(new_n433), .A3(new_n514), .A4(new_n434), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n582), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n581), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n618), .B2(new_n620), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n428), .A2(new_n429), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n588), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n583), .A2(new_n622), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n296), .B1(new_n242), .B2(new_n244), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n250), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n223), .A2(new_n296), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT91), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n223), .A2(new_n296), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n642), .A2(new_n635), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n637), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n634), .A2(KEYINPUT18), .A3(new_n635), .A4(new_n638), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(KEYINPUT92), .A3(new_n646), .ZN(new_n649));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G197gat), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT11), .B(G169gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT12), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n647), .A2(new_n646), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n656), .B(new_n641), .C1(KEYINPUT92), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n268), .A2(new_n660), .A3(new_n307), .A4(new_n324), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n326), .A2(new_n632), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n579), .A2(new_n581), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(G1gat), .Z(G1324gat));
  INV_X1    g464(.A(new_n539), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G8gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n667), .ZN(new_n671));
  MUX2_X1   g470(.A(new_n669), .B(new_n671), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n662), .B2(new_n436), .ZN(new_n673));
  INV_X1    g472(.A(new_n628), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n662), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n662), .A2(new_n518), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n261), .A2(new_n267), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n632), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n659), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n682), .A2(new_n307), .A3(new_n323), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n663), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n211), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n632), .A2(new_n680), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n632), .A2(KEYINPUT44), .A3(new_n680), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n683), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n691), .A2(KEYINPUT103), .A3(new_n683), .A4(new_n692), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n695), .A2(new_n685), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n688), .B1(new_n211), .B2(new_n697), .ZN(G1328gat));
  NAND3_X1  g497(.A1(new_n684), .A2(new_n212), .A3(new_n539), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT46), .Z(new_n700));
  AND3_X1   g499(.A1(new_n695), .A2(new_n539), .A3(new_n696), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n212), .B2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n681), .A2(new_n703), .A3(new_n628), .A4(new_n683), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT105), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n693), .B2(new_n436), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n436), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n710), .A3(new_n696), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n711), .A2(KEYINPUT104), .A3(G43gat), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT104), .B1(new_n711), .B2(G43gat), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n713), .A3(new_n705), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n693), .B2(new_n588), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n518), .A2(G50gat), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT106), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n684), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n518), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n695), .A2(new_n721), .A3(new_n696), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n722), .A2(G50gat), .B1(new_n684), .B2(new_n718), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n723), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g523(.A1(new_n682), .A2(new_n323), .ZN(new_n725));
  INV_X1    g524(.A(new_n307), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n726), .A3(new_n680), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n632), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(KEYINPUT107), .A3(new_n632), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n663), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n269), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n666), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT108), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n732), .B2(new_n436), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n628), .A2(new_n275), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g543(.A1(new_n732), .A2(new_n518), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n276), .ZN(G1335gat));
  NOR3_X1   g545(.A1(new_n689), .A2(new_n659), .A3(new_n307), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT51), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(new_n229), .A3(new_n685), .A4(new_n323), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n691), .A2(new_n692), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n307), .A2(new_n659), .A3(new_n324), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n663), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n539), .A3(new_n751), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n230), .B1(new_n755), .B2(KEYINPUT110), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT110), .B2(new_n755), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n323), .A2(new_n230), .A3(new_n539), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT109), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(new_n748), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n748), .A2(new_n759), .B1(new_n755), .B2(G92gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(G1337gat));
  NOR3_X1   g563(.A1(new_n324), .A2(new_n674), .A3(G99gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G99gat), .B1(new_n752), .B2(new_n436), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(G1338gat));
  OAI21_X1  g567(.A(G106gat), .B1(new_n752), .B2(new_n588), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n324), .A2(G106gat), .A3(new_n588), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n748), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(KEYINPUT111), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT53), .B(G106gat), .C1(new_n752), .C2(new_n518), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT111), .A2(KEYINPUT53), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n748), .B2(new_n770), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n776), .ZN(G1339gat));
  INV_X1    g576(.A(new_n316), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n314), .A2(new_n310), .A3(new_n315), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT54), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n320), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n316), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n321), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n314), .A2(new_n310), .A3(new_n315), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n787), .A2(new_n316), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n314), .A2(new_n315), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n309), .A3(new_n782), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n320), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n786), .C1(new_n789), .C2(new_n792), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n785), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n643), .A2(new_n645), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT114), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n653), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n641), .A2(new_n646), .A3(new_n647), .A4(new_n657), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n323), .A3(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n797), .A2(new_n659), .B1(KEYINPUT115), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n680), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n801), .A2(new_n802), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n680), .A2(new_n797), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n726), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n325), .A2(new_n659), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n721), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n663), .A2(new_n539), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n674), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n682), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n663), .B1(new_n809), .B2(new_n811), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n624), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n666), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n659), .A2(new_n335), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT116), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n817), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1340gat));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n323), .A3(new_n815), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n826), .A2(new_n827), .A3(G120gat), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n826), .B2(G120gat), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n323), .A2(new_n336), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n828), .A2(new_n829), .B1(new_n820), .B2(new_n830), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n816), .B2(new_n726), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n307), .A2(new_n342), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n820), .B2(new_n833), .ZN(G1342gat));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n340), .A3(new_n666), .A4(new_n680), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n816), .B2(new_n268), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(KEYINPUT56), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n814), .A2(new_n710), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n518), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n793), .A2(new_n321), .A3(new_n784), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n658), .B2(new_n655), .ZN(new_n844));
  INV_X1    g643(.A(new_n803), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n268), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n680), .A2(new_n797), .A3(new_n807), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n307), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n842), .B1(new_n848), .B2(new_n810), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT119), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n851), .B(new_n842), .C1(new_n848), .C2(new_n810), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n797), .A2(new_n659), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n805), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n808), .B1(new_n856), .B2(new_n268), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n811), .B1(new_n857), .B2(new_n307), .ZN(new_n858));
  INV_X1    g657(.A(new_n588), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n659), .B(new_n840), .C1(new_n853), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G141gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n710), .A2(new_n588), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n818), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n539), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n472), .A3(new_n659), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n862), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1344gat));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n474), .A3(new_n323), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n588), .B1(new_n809), .B2(new_n811), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(new_n841), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n326), .A2(new_n682), .A3(new_n661), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n841), .B(new_n721), .C1(new_n876), .C2(new_n848), .ZN(new_n877));
  INV_X1    g676(.A(new_n840), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT120), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n324), .B1(new_n878), .B2(KEYINPUT120), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n875), .A2(new_n877), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n873), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n323), .B(new_n840), .C1(new_n853), .C2(new_n860), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(new_n873), .A3(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n872), .B1(new_n882), .B2(new_n884), .ZN(G1345gat));
  OAI21_X1  g684(.A(new_n840), .B1(new_n853), .B2(new_n860), .ZN(new_n886));
  OAI21_X1  g685(.A(G155gat), .B1(new_n886), .B2(new_n726), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n865), .A2(new_n302), .A3(new_n307), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1346gat));
  NOR4_X1   g688(.A1(new_n864), .A2(G162gat), .A3(new_n539), .A4(new_n268), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G162gat), .B1(new_n886), .B2(new_n268), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1347gat));
  NAND2_X1  g693(.A1(new_n663), .A2(new_n539), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n674), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n812), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(G169gat), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n898), .A3(new_n682), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n685), .B1(new_n809), .B2(new_n811), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n624), .A2(new_n539), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n659), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n899), .B1(new_n898), .B2(new_n904), .ZN(G1348gat));
  OAI21_X1  g704(.A(G176gat), .B1(new_n897), .B2(new_n324), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n324), .A2(G176gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n902), .B2(new_n907), .ZN(G1349gat));
  OAI21_X1  g707(.A(G183gat), .B1(new_n897), .B2(new_n726), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n307), .A2(new_n394), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(G1350gat));
  NOR3_X1   g712(.A1(new_n902), .A2(G190gat), .A3(new_n268), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n812), .A2(new_n680), .A3(new_n896), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G190gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n915), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n917), .A2(new_n916), .A3(G190gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n895), .A2(new_n710), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n877), .B(new_n923), .C1(new_n874), .C2(new_n841), .ZN(new_n924));
  INV_X1    g723(.A(G197gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(new_n682), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n863), .A2(new_n539), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  AND2_X1   g727(.A1(new_n900), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n659), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n926), .A2(new_n930), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n324), .A2(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n900), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT125), .Z(new_n935));
  NOR2_X1   g734(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT126), .ZN(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n924), .B2(new_n324), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n929), .A2(new_n456), .A3(new_n307), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n924), .A2(new_n726), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT63), .B(G211gat), .C1(new_n924), .C2(new_n726), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(G1354gat));
  OAI21_X1  g744(.A(G218gat), .B1(new_n924), .B2(new_n268), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n457), .A3(new_n680), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1355gat));
endmodule


