//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G137), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n462), .B(KEYINPUT66), .C1(new_n464), .C2(new_n463), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n460), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AOI211_X1 g050(.A(KEYINPUT67), .B(new_n473), .C1(new_n467), .C2(new_n468), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n463), .A2(new_n464), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n479), .B(KEYINPUT68), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n470), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(new_n489), .B2(G124), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OR2_X1    g069(.A1(new_n470), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n463), .B2(new_n464), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n463), .B2(new_n464), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n503), .B(new_n506), .C1(new_n464), .C2(new_n463), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT69), .A3(G651), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(new_n513), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G50), .A3(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT5), .B1(KEYINPUT70), .B2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT71), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(KEYINPUT5), .A4(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OAI221_X1 g098(.A(new_n515), .B1(new_n521), .B2(new_n522), .C1(new_n523), .C2(new_n510), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  INV_X1    g100(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n514), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n520), .A2(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n528), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n521), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n510), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n510), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n528), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n526), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n518), .A2(new_n519), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(G651), .A2(new_n557), .B1(new_n526), .B2(G91), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n514), .A2(KEYINPUT73), .A3(G53), .A4(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT72), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n514), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n559), .A2(KEYINPUT72), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n558), .B1(new_n567), .B2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  NAND3_X1  g145(.A1(new_n514), .A2(new_n520), .A3(G87), .ZN(new_n571));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n518), .A2(new_n572), .A3(new_n519), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n511), .A2(new_n513), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n575), .A2(G49), .A3(G543), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n574), .A3(new_n577), .ZN(G288));
  NAND3_X1  g153(.A1(new_n514), .A2(new_n520), .A3(G86), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n518), .B2(new_n519), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n510), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n528), .A2(G47), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n526), .A2(G85), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G290));
  XOR2_X1   g166(.A(KEYINPUT75), .B(G66), .Z(new_n592));
  NOR2_X1   g167(.A1(new_n555), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G79), .ZN(new_n594));
  INV_X1    g169(.A(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT76), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n598));
  OAI221_X1 g173(.A(new_n598), .B1(new_n594), .B2(new_n595), .C1(new_n555), .C2(new_n592), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n599), .A3(G651), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n521), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n514), .A2(new_n520), .A3(KEYINPUT10), .A4(G92), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n603), .A2(new_n604), .B1(G54), .B2(new_n528), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(new_n558), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n563), .A2(new_n566), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT74), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n611), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n611), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(new_n606), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g200(.A1(new_n479), .A2(new_n471), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OAI22_X1  g203(.A1(new_n628), .A2(KEYINPUT13), .B1(KEYINPUT78), .B2(G2100), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(KEYINPUT13), .B2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n491), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n489), .A2(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(KEYINPUT80), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n637));
  OR3_X1    g212(.A1(new_n637), .A2(new_n470), .A3(G111), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(KEYINPUT80), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n637), .B1(new_n470), .B2(G111), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n636), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n633), .A2(new_n634), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n632), .A2(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n650), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n678), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n685), .C1(new_n675), .C2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT32), .B(G1981), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(G288), .A2(KEYINPUT89), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n571), .A2(new_n574), .A3(new_n699), .A4(new_n577), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G23), .B(new_n701), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT86), .B(G16), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  NOR4_X1   g284(.A1(new_n696), .A2(new_n697), .A3(new_n704), .A4(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n491), .A2(G131), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G107), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n489), .B2(G119), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT85), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n706), .A2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G290), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n706), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n712), .A2(new_n713), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT36), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n705), .A2(G20), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT23), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n616), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G1956), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n714), .A2(G32), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n489), .A2(G129), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  INV_X1    g321(.A(new_n471), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n747), .A2(new_n748), .A3(G105), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n747), .B2(G105), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n491), .B2(G141), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n741), .B1(new_n754), .B2(new_n714), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n755), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n714), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT3), .B(G2104), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n762), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n763), .B2(new_n470), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n491), .B2(G139), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(new_n714), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2072), .ZN(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT30), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n768), .B2(KEYINPUT30), .ZN(new_n770));
  OR2_X1    g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n642), .B2(new_n714), .ZN(new_n774));
  NOR2_X1   g349(.A1(G27), .A2(G29), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G164), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n767), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n706), .A2(G19), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n548), .B2(new_n706), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1341), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n737), .A2(G21), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G168), .B2(new_n737), .ZN(new_n783));
  INV_X1    g358(.A(G1966), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(KEYINPUT24), .B2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n483), .B2(G29), .ZN(new_n788));
  INV_X1    g363(.A(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n778), .A2(new_n781), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n714), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n714), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT29), .B(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n737), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n737), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1961), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n758), .A2(new_n791), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n788), .A2(new_n789), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n714), .A2(G26), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n491), .A2(G140), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n489), .A2(G128), .ZN(new_n805));
  OR2_X1    g380(.A1(G104), .A2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n806), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n808), .A2(KEYINPUT91), .A3(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(KEYINPUT91), .B1(new_n808), .B2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2067), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n737), .A2(G4), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n619), .B2(new_n737), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1348), .ZN(new_n817));
  AND4_X1   g392(.A1(new_n740), .A2(new_n799), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n734), .A2(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NAND2_X1  g395(.A1(new_n619), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n510), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n514), .A2(G55), .A3(G543), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n521), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(KEYINPUT96), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(KEYINPUT96), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n548), .B(new_n824), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n547), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n822), .B(new_n833), .Z(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n835), .A2(new_n836), .A3(G860), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n831), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  NAND2_X1  g415(.A1(new_n491), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n489), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n470), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n723), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n628), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n628), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(KEYINPUT100), .A3(new_n848), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n765), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n753), .B(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(new_n808), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n762), .A2(new_n499), .B1(new_n495), .B2(new_n497), .ZN(new_n857));
  INV_X1    g432(.A(new_n507), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n506), .B1(new_n762), .B2(new_n503), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n808), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n860), .B1(new_n856), .B2(new_n861), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n851), .B(new_n852), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n493), .B(new_n642), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n483), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n867), .B(new_n868), .Z(new_n869));
  INV_X1    g444(.A(new_n864), .ZN(new_n870));
  INV_X1    g445(.A(new_n852), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n862), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n865), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n869), .B1(new_n865), .B2(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT40), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n874), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n879), .A2(new_n880), .A3(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(G395));
  XNOR2_X1  g457(.A(G290), .B(KEYINPUT104), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n701), .ZN(new_n884));
  XNOR2_X1  g459(.A(G305), .B(G303), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(KEYINPUT105), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n885), .B(KEYINPUT105), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n558), .B(new_n606), .C1(new_n567), .C2(new_n568), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT101), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n614), .A2(new_n615), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n558), .A4(new_n606), .ZN(new_n897));
  NAND2_X1  g472(.A1(G299), .A2(new_n619), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(KEYINPUT102), .A3(new_n900), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n905));
  XOR2_X1   g480(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n833), .B(new_n622), .Z(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n905), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n892), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g489(.A(KEYINPUT106), .B(new_n912), .C1(new_n909), .C2(new_n910), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n891), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n909), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n892), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n889), .B(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n607), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n831), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(G868), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT107), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  INV_X1    g500(.A(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(new_n910), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n901), .A2(new_n902), .B1(new_n905), .B2(new_n907), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n904), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT106), .B1(new_n929), .B2(new_n912), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n919), .B1(new_n918), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n915), .A2(new_n891), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n925), .B(new_n926), .C1(new_n933), .C2(new_n607), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n924), .A2(new_n934), .ZN(G295));
  OAI21_X1  g510(.A(new_n926), .B1(new_n933), .B2(new_n607), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  XOR2_X1   g512(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n938));
  NAND2_X1  g513(.A1(new_n833), .A2(G171), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n830), .A2(new_n832), .A3(G301), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(G168), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n830), .A2(new_n832), .A3(G301), .ZN(new_n942));
  AOI21_X1  g517(.A(G301), .B1(new_n830), .B2(new_n832), .ZN(new_n943));
  OAI21_X1  g518(.A(G286), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n905), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n949), .B2(new_n889), .ZN(new_n950));
  INV_X1    g525(.A(new_n889), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n951), .B(new_n946), .C1(new_n947), .C2(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n938), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n948), .B1(new_n928), .B2(new_n904), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n954), .A2(new_n889), .A3(new_n945), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n894), .A2(new_n897), .A3(new_n898), .A4(new_n900), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n944), .A2(new_n941), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n899), .A2(new_n907), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n945), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n874), .B1(new_n959), .B2(new_n951), .ZN(new_n960));
  INV_X1    g535(.A(new_n938), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n955), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n937), .B1(new_n953), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  INV_X1    g539(.A(new_n948), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n945), .B1(new_n909), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n961), .B1(new_n966), .B2(new_n951), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n937), .B1(new_n950), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n955), .B2(new_n960), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n889), .B1(new_n954), .B2(new_n945), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(new_n952), .A3(new_n874), .A4(new_n938), .ZN(new_n972));
  AND4_X1   g547(.A1(new_n964), .A2(new_n969), .A3(new_n972), .A4(KEYINPUT44), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n963), .B1(new_n970), .B2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n481), .B2(G2105), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n477), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(G164), .B2(G1384), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n753), .B(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n808), .B(G2067), .Z(new_n983));
  AND2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n723), .B(new_n725), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(G290), .B(G1986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT110), .ZN(new_n989));
  NAND3_X1  g564(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(G166), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n976), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n860), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n1000), .B2(new_n978), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n505), .A2(new_n507), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1002), .B2(new_n857), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n477), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT111), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n860), .A2(new_n1009), .A3(new_n999), .ZN(new_n1013));
  INV_X1    g588(.A(new_n468), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT66), .B1(new_n762), .B2(new_n462), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n474), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT67), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n469), .A2(new_n460), .A3(new_n474), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1013), .A2(new_n1017), .A3(new_n1018), .A4(new_n976), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1012), .A2(G2090), .A3(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n997), .B(G8), .C1(new_n1007), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n581), .B2(new_n585), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n585), .A2(new_n1023), .A3(new_n579), .A4(new_n580), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT113), .B(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1017), .A2(new_n1003), .A3(new_n1018), .A4(new_n976), .ZN(new_n1030));
  INV_X1    g605(.A(new_n585), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n579), .A2(new_n580), .ZN(new_n1032));
  OAI21_X1  g607(.A(G1981), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n698), .A2(G1976), .A3(new_n700), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(new_n1030), .A3(new_n1029), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1030), .A3(new_n1029), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1035), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1025), .B(KEYINPUT114), .Z(new_n1043));
  NOR2_X1   g618(.A1(G288), .A2(G1976), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1030), .A2(new_n1029), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n1021), .A2(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n1049));
  INV_X1    g624(.A(G2090), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1019), .A2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1050), .A2(new_n1052), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1035), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1021), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n976), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n477), .A2(new_n979), .A3(KEYINPUT115), .A4(new_n976), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1004), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n784), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n789), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(G168), .A3(new_n1029), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1048), .B1(new_n1056), .B2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1062), .A2(new_n784), .B1(new_n1064), .B2(new_n789), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1069), .A2(G286), .A3(new_n1028), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1019), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1071), .A2(new_n1050), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n994), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1042), .B1(new_n997), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1070), .A2(new_n1075), .A3(KEYINPUT116), .A4(new_n1054), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1068), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1074), .A2(new_n997), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1070), .A2(new_n1075), .A3(new_n1079), .A4(KEYINPUT63), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1047), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n1052), .B2(G1956), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(new_n739), .C1(new_n1019), .C2(new_n1051), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n558), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(new_n613), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT56), .B(G2072), .Z(new_n1090));
  OR2_X1    g665(.A1(new_n1005), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1348), .B1(new_n1094), .B2(new_n1071), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1030), .A2(G2067), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n619), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1084), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n477), .A2(new_n1099), .A3(new_n976), .A4(new_n1013), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1083), .B1(new_n1100), .B2(new_n739), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1091), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n616), .A2(new_n1086), .B1(new_n613), .B2(new_n1087), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1093), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1348), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1096), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n600), .B2(new_n605), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n600), .A2(new_n605), .A3(new_n1110), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1111), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1116), .A2(KEYINPUT60), .A3(new_n1108), .A4(new_n1107), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT121), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1112), .A2(new_n1114), .A3(new_n1117), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n547), .B1(new_n1122), .B2(KEYINPUT59), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND3_X1  g699(.A1(new_n1030), .A2(KEYINPUT118), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1005), .B2(G1996), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT118), .B1(new_n1030), .B2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1122), .B2(KEYINPUT59), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(new_n1123), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1119), .A2(new_n1121), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1104), .A2(new_n1092), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT61), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1104), .A2(new_n1092), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1105), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G286), .A2(new_n1029), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1069), .B2(new_n994), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT51), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1028), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1146), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT122), .B(new_n1148), .C1(new_n1069), .C2(new_n1028), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1142), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1140), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1066), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT124), .B1(new_n475), .B2(new_n476), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1017), .A2(new_n1018), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1001), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1001), .A2(new_n1154), .A3(new_n1156), .A4(KEYINPUT125), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT53), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(G2078), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1004), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G2078), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1001), .A2(new_n1166), .A3(new_n477), .A4(new_n1004), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1162), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT123), .B(G1961), .Z(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(G301), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1060), .A2(new_n1061), .A3(new_n1004), .A4(new_n1163), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT54), .B1(new_n1174), .B2(G171), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1054), .B(new_n1075), .C1(new_n1172), .C2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1165), .A2(new_n1171), .A3(G301), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1174), .A2(G171), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT54), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1153), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1081), .B1(new_n1139), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT126), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1150), .A2(new_n1186), .A3(new_n1152), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1056), .A2(new_n1178), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1153), .A2(new_n1190), .A3(KEYINPUT62), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1185), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n989), .B1(new_n1183), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n980), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n808), .A2(G2067), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n718), .A2(new_n725), .A3(new_n722), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1195), .B1(new_n984), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1194), .B1(new_n984), .B2(new_n985), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n980), .A2(new_n731), .A3(new_n729), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT48), .Z(new_n1201));
  OAI22_X1  g776(.A1(new_n1194), .A2(new_n1198), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1194), .B1(new_n983), .B2(new_n754), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT46), .B1(new_n1194), .B2(G1996), .ZN(new_n1204));
  OR3_X1    g779(.A1(new_n1194), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT47), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT127), .B1(new_n1193), .B2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n988), .B(KEYINPUT110), .Z(new_n1211));
  AOI21_X1  g786(.A(new_n1190), .B1(new_n1153), .B2(KEYINPUT62), .ZN(new_n1212));
  AOI211_X1 g787(.A(KEYINPUT126), .B(new_n1186), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1211), .B1(new_n1215), .B2(new_n1182), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1216), .A2(new_n1217), .A3(new_n1208), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1210), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g794(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1221), .B1(new_n879), .B2(new_n876), .ZN(new_n1222));
  NOR2_X1   g796(.A1(new_n953), .A2(new_n962), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n1222), .A2(new_n1223), .ZN(G308));
  OAI221_X1 g798(.A(new_n1221), .B1(new_n879), .B2(new_n876), .C1(new_n953), .C2(new_n962), .ZN(G225));
endmodule


