//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1' ..
//Module:
 module locked_c1908( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  , KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0);
input KEYINPUT0;
input KEYINPUT1;
input KEYINPUT2;
input KEYINPUT3;
input KEYINPUT4;
input KEYINPUT5;
input KEYINPUT6;
input KEYINPUT7;
input KEYINPUT8;
input KEYINPUT9;
input KEYINPUT10;
input KEYINPUT11;
input KEYINPUT12;
input KEYINPUT13;
input KEYINPUT14;
input KEYINPUT15;
input KEYINPUT16;
input KEYINPUT17;
input KEYINPUT18;
input KEYINPUT19;
input KEYINPUT20;
input KEYINPUT21;
input KEYINPUT22;
input KEYINPUT23;
input KEYINPUT24;
input KEYINPUT25;
input KEYINPUT26;
input KEYINPUT27;
input KEYINPUT28;
input KEYINPUT29;
input KEYINPUT30;
input KEYINPUT31;
input KEYINPUT32;
input KEYINPUT33;
input KEYINPUT34;
input KEYINPUT35;
input KEYINPUT36;
input KEYINPUT37;
input KEYINPUT38;
input KEYINPUT39;
input KEYINPUT40;
input KEYINPUT41;
input KEYINPUT42;
input KEYINPUT43;
input KEYINPUT44;
input KEYINPUT45;
input KEYINPUT46;
input KEYINPUT47;
input KEYINPUT48;
input KEYINPUT49;
input KEYINPUT50;
input KEYINPUT51;
input KEYINPUT52;
input KEYINPUT53;
input KEYINPUT54;
input KEYINPUT55;
input KEYINPUT56;
input KEYINPUT57;
input KEYINPUT58;
input KEYINPUT59;
input KEYINPUT60;
input KEYINPUT61;
input KEYINPUT62;
input KEYINPUT63;
//Header:
   input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n335_, new_n336_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n343_, new_n345_, new_n347_, new_n348_, new_n350_, new_n352_,
    new_n353_, new_n355_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n369_, new_n370_, new_n371_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n424_,
    new_n425_, new_n426_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_;
wire RLL_wire_A_0;
wire RLL_wire_A_1;
wire RLL_wire_A_2;
wire RLL_wire_A_3;
wire RLL_wire_A_4;
wire RLL_wire_A_5;
wire RLL_wire_A_6;
wire RLL_wire_A_7;
wire RLL_wire_A_8;
wire RLL_wire_A_9;
wire RLL_wire_A_10;
wire RLL_wire_A_11;
wire RLL_wire_A_12;
wire RLL_wire_A_13;
wire RLL_wire_A_14;
wire RLL_wire_A_15;
wire RLL_wire_A_16;
wire RLL_wire_A_17;
wire RLL_wire_A_18;
wire RLL_wire_A_19;
wire RLL_wire_A_20;
wire RLL_wire_A_21;
wire RLL_wire_A_22;
wire RLL_wire_A_23;
wire RLL_wire_A_24;
wire RLL_wire_A_25;
wire RLL_wire_A_26;
wire RLL_wire_A_27;
wire RLL_wire_A_28;
wire RLL_wire_A_29;
wire RLL_wire_A_30;
wire RLL_wire_A_31;
wire RLL_wire_A_32;
wire RLL_wire_A_33;
wire RLL_wire_A_34;
wire RLL_wire_A_35;
wire RLL_wire_A_36;
wire RLL_wire_A_37;
wire RLL_wire_A_38;
wire RLL_wire_A_39;
wire RLL_wire_A_40;
wire RLL_wire_A_41;
wire RLL_wire_A_42;
wire RLL_wire_A_43;
wire RLL_wire_A_44;
wire RLL_wire_A_45;
wire RLL_wire_A_46;
wire RLL_wire_A_47;
wire RLL_wire_A_48;
wire RLL_wire_A_49;
wire RLL_wire_A_50;
wire RLL_wire_A_51;
wire RLL_wire_A_52;
wire RLL_wire_A_53;
wire RLL_wire_A_54;
wire RLL_wire_A_55;
wire RLL_wire_A_56;
wire RLL_wire_A_57;
wire RLL_wire_A_58;
wire RLL_wire_A_59;
wire RLL_wire_A_60;
wire RLL_wire_A_61;
wire RLL_wire_A_62;
wire RLL_wire_A_63;

//Body:
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n59_));
  INV_X1    g001(.A(new_n59_), .ZN(new_n60_));
  INV_X1    g002(.A(G902), .ZN(new_n61_));
  INV_X1    g003(.A(G224), .ZN(new_n62_));
  NOR2_X1   g004(.A1(new_n62_), .A2(G953), .ZN(new_n63_));
  INV_X1    g005(.A(G128), .ZN(new_n64_));
  INV_X1    g006(.A(G146), .ZN(new_n65_));
  NAND2_X1  g007(.A1(new_n65_), .A2(G143), .ZN(new_n66_));
  INV_X1    g008(.A(G143), .ZN(new_n67_));
  NAND2_X1  g009(.A1(new_n67_), .A2(G146), .ZN(new_n68_));
  AND3_X1   g010(.A1(new_n66_), .A2(new_n68_), .A3(new_n64_), .ZN(new_n69_));
  AOI21_X1  g011(.A(new_n64_), .B1(new_n66_), .B2(new_n68_), .ZN(RLL_wire_A_0));
  XNOR2_X1 RLL_XNOR_0 (.A(RLL_wire_A_0), .B(KEYINPUT0), .ZN(new_n70_) );
  OAI21_X1  g012(.A(G125), .B1(new_n69_), .B2(new_n70_), .ZN(new_n71_));
  INV_X1    g013(.A(G125), .ZN(new_n72_));
  NAND3_X1  g014(.A1(new_n66_), .A2(new_n68_), .A3(new_n64_), .ZN(new_n73_));
  NOR2_X1   g015(.A1(new_n67_), .A2(G146), .ZN(new_n74_));
  NOR2_X1   g016(.A1(new_n65_), .A2(G143), .ZN(RLL_wire_A_1));
  XOR2_X1 RLL_XOR_1 (.A(RLL_wire_A_1), .B(KEYINPUT1), .Z(new_n75_) );
  OAI21_X1  g017(.A(G128), .B1(new_n74_), .B2(new_n75_), .ZN(new_n76_));
  NAND3_X1  g018(.A1(new_n76_), .A2(new_n72_), .A3(new_n73_), .ZN(new_n77_));
  NAND3_X1  g019(.A1(new_n71_), .A2(new_n77_), .A3(new_n63_), .ZN(new_n78_));
  INV_X1    g020(.A(new_n78_), .ZN(new_n79_));
  AOI21_X1  g021(.A(new_n63_), .B1(new_n71_), .B2(new_n77_), .ZN(new_n80_));
  XNOR2_X1  g022(.A(G110), .B(G122), .ZN(new_n81_));
  INV_X1    g023(.A(G113), .ZN(RLL_wire_A_2));
  XNOR2_X1 RLL_XNOR_2 (.A(RLL_wire_A_2), .B(KEYINPUT2), .ZN(new_n82_) );
  INV_X1    g024(.A(G119), .ZN(new_n83_));
  NAND2_X1  g025(.A1(new_n83_), .A2(G116), .ZN(new_n84_));
  INV_X1    g026(.A(G116), .ZN(new_n85_));
  NAND2_X1  g027(.A1(new_n85_), .A2(G119), .ZN(new_n86_));
  NAND3_X1  g028(.A1(new_n84_), .A2(new_n86_), .A3(new_n82_), .ZN(new_n87_));
  INV_X1    g029(.A(new_n87_), .ZN(new_n88_));
  AOI21_X1  g030(.A(new_n82_), .B1(new_n84_), .B2(new_n86_), .ZN(new_n89_));
  INV_X1    g031(.A(G101), .ZN(new_n90_));
  INV_X1    g032(.A(G107), .ZN(new_n91_));
  NAND2_X1  g033(.A1(new_n91_), .A2(G104), .ZN(RLL_wire_A_3));
  XOR2_X1 RLL_XOR_3 (.A(RLL_wire_A_3), .B(KEYINPUT3), .Z(new_n92_) );
  INV_X1    g034(.A(G104), .ZN(new_n93_));
  NAND2_X1  g035(.A1(new_n93_), .A2(G107), .ZN(new_n94_));
  AND3_X1   g036(.A1(new_n92_), .A2(new_n94_), .A3(new_n90_), .ZN(new_n95_));
  AOI21_X1  g037(.A(new_n90_), .B1(new_n92_), .B2(new_n94_), .ZN(RLL_wire_A_4));
  XNOR2_X1 RLL_XNOR_4 (.A(RLL_wire_A_4), .B(KEYINPUT4), .ZN(new_n96_) );
  OAI22_X1  g038(.A1(new_n88_), .A2(new_n89_), .B1(new_n95_), .B2(new_n96_), .ZN(new_n97_));
  NOR2_X1   g039(.A1(new_n85_), .A2(G119), .ZN(RLL_wire_A_5));
  XNOR2_X1 RLL_XNOR_5 (.A(RLL_wire_A_5), .B(KEYINPUT5), .ZN(new_n98_) );
  NOR2_X1   g040(.A1(new_n83_), .A2(G116), .ZN(new_n99_));
  OAI21_X1  g041(.A(G113), .B1(new_n98_), .B2(new_n99_), .ZN(new_n100_));
  NAND3_X1  g042(.A1(new_n92_), .A2(new_n94_), .A3(new_n90_), .ZN(new_n101_));
  NOR2_X1   g043(.A1(new_n93_), .A2(G107), .ZN(new_n102_));
  NOR2_X1   g044(.A1(new_n91_), .A2(G104), .ZN(new_n103_));
  OAI21_X1  g045(.A(G101), .B1(new_n102_), .B2(new_n103_), .ZN(new_n104_));
  NAND4_X1  g046(.A1(new_n100_), .A2(new_n104_), .A3(new_n87_), .A4(new_n101_), .ZN(new_n105_));
  AND3_X1   g047(.A1(new_n97_), .A2(new_n105_), .A3(new_n81_), .ZN(new_n106_));
  AOI21_X1  g048(.A(new_n81_), .B1(new_n97_), .B2(new_n105_), .ZN(RLL_wire_A_6));
  XNOR2_X1 RLL_XNOR_6 (.A(RLL_wire_A_6), .B(KEYINPUT6), .ZN(new_n107_) );
  OAI22_X1  g049(.A1(new_n106_), .A2(new_n107_), .B1(new_n79_), .B2(new_n80_), .ZN(new_n108_));
  INV_X1    g050(.A(new_n63_), .ZN(new_n109_));
  NAND2_X1  g051(.A1(new_n71_), .A2(new_n77_), .ZN(RLL_wire_A_7));
  XNOR2_X1 RLL_XNOR_7 (.A(RLL_wire_A_7), .B(KEYINPUT7), .ZN(new_n110_) );
  NAND2_X1  g052(.A1(new_n110_), .A2(new_n109_), .ZN(new_n111_));
  NAND3_X1  g053(.A1(new_n97_), .A2(new_n105_), .A3(new_n81_), .ZN(new_n112_));
  INV_X1    g054(.A(new_n81_), .ZN(RLL_wire_A_8));
  XOR2_X1 RLL_XOR_8 (.A(RLL_wire_A_8), .B(KEYINPUT8), .Z(new_n113_) );
  AOI22_X1  g055(.A1(new_n87_), .A2(new_n100_), .B1(new_n104_), .B2(new_n101_), .ZN(new_n114_));
  AND4_X1   g056(.A1(new_n87_), .A2(new_n100_), .A3(new_n104_), .A4(new_n101_), .ZN(new_n115_));
  OAI21_X1  g057(.A(new_n113_), .B1(new_n115_), .B2(new_n114_), .ZN(new_n116_));
  NAND4_X1  g058(.A1(new_n116_), .A2(new_n78_), .A3(new_n111_), .A4(new_n112_), .ZN(new_n117_));
  NAND3_X1  g059(.A1(new_n108_), .A2(new_n117_), .A3(new_n61_), .ZN(new_n118_));
  OAI21_X1  g060(.A(G210), .B1(G237), .B2(G902), .ZN(new_n119_));
  INV_X1    g061(.A(new_n119_), .ZN(new_n120_));
  NAND2_X1  g062(.A1(new_n118_), .A2(new_n120_), .ZN(new_n121_));
  NAND4_X1  g063(.A1(new_n108_), .A2(new_n117_), .A3(new_n61_), .A4(new_n119_), .ZN(new_n122_));
  AOI21_X1  g064(.A(new_n60_), .B1(new_n121_), .B2(new_n122_), .ZN(new_n123_));
  INV_X1    g065(.A(G234), .ZN(RLL_wire_A_9));
  XOR2_X1 RLL_XOR_9 (.A(RLL_wire_A_9), .B(KEYINPUT9), .Z(new_n124_) );
  OAI21_X1  g066(.A(G221), .B1(new_n124_), .B2(G902), .ZN(new_n125_));
  INV_X1    g067(.A(new_n125_), .ZN(new_n126_));
  XNOR2_X1  g068(.A(G110), .B(G140), .ZN(new_n127_));
  INV_X1    g069(.A(G953), .ZN(new_n128_));
  AND2_X1   g070(.A1(new_n128_), .A2(G227), .ZN(new_n129_));
  XNOR2_X1  g071(.A(new_n127_), .B(new_n129_), .ZN(new_n130_));
  NAND4_X1  g072(.A1(new_n76_), .A2(new_n104_), .A3(new_n73_), .A4(new_n101_), .ZN(RLL_wire_A_10));
  XNOR2_X1 RLL_XNOR_10 (.A(RLL_wire_A_10), .B(KEYINPUT10), .ZN(new_n131_) );
  INV_X1    g073(.A(G131), .ZN(new_n132_));
  INV_X1    g074(.A(G137), .ZN(new_n133_));
  NAND2_X1  g075(.A1(new_n133_), .A2(G134), .ZN(RLL_wire_A_11));
  XNOR2_X1 RLL_XNOR_11 (.A(RLL_wire_A_11), .B(KEYINPUT11), .ZN(new_n134_) );
  INV_X1    g076(.A(G134), .ZN(new_n135_));
  NAND2_X1  g077(.A1(new_n135_), .A2(G137), .ZN(new_n136_));
  AOI21_X1  g078(.A(new_n132_), .B1(new_n134_), .B2(new_n136_), .ZN(new_n137_));
  AND3_X1   g079(.A1(new_n134_), .A2(new_n136_), .A3(new_n132_), .ZN(new_n138_));
  NOR2_X1   g080(.A1(new_n138_), .A2(new_n137_), .ZN(new_n139_));
  OAI22_X1  g081(.A1(new_n69_), .A2(new_n70_), .B1(new_n95_), .B2(new_n96_), .ZN(new_n140_));
  AND3_X1   g082(.A1(new_n140_), .A2(new_n131_), .A3(new_n139_), .ZN(new_n141_));
  AOI21_X1  g083(.A(new_n139_), .B1(new_n140_), .B2(new_n131_), .ZN(new_n142_));
  NOR3_X1   g084(.A1(new_n141_), .A2(new_n142_), .A3(new_n130_), .ZN(new_n143_));
  INV_X1    g085(.A(new_n130_), .ZN(new_n144_));
  AND4_X1   g086(.A1(new_n73_), .A2(new_n76_), .A3(new_n104_), .A4(new_n101_), .ZN(new_n145_));
  INV_X1    g087(.A(new_n139_), .ZN(new_n146_));
  AOI22_X1  g088(.A1(new_n73_), .A2(new_n76_), .B1(new_n104_), .B2(new_n101_), .ZN(new_n147_));
  OAI21_X1  g089(.A(new_n146_), .B1(new_n145_), .B2(new_n147_), .ZN(RLL_wire_A_12));
  XOR2_X1 RLL_XOR_12 (.A(RLL_wire_A_12), .B(KEYINPUT12), .Z(new_n148_) );
  NAND3_X1  g090(.A1(new_n140_), .A2(new_n131_), .A3(new_n139_), .ZN(new_n149_));
  AOI21_X1  g091(.A(new_n144_), .B1(new_n148_), .B2(new_n149_), .ZN(new_n150_));
  OAI21_X1  g092(.A(new_n61_), .B1(new_n143_), .B2(new_n150_), .ZN(new_n151_));
  NAND2_X1  g093(.A1(new_n151_), .A2(G469), .ZN(new_n152_));
  INV_X1    g094(.A(G469), .ZN(new_n153_));
  OAI21_X1  g095(.A(new_n130_), .B1(new_n141_), .B2(new_n142_), .ZN(new_n154_));
  NAND3_X1  g096(.A1(new_n148_), .A2(new_n144_), .A3(new_n149_), .ZN(new_n155_));
  NAND2_X1  g097(.A1(new_n154_), .A2(new_n155_), .ZN(new_n156_));
  NAND3_X1  g098(.A1(new_n156_), .A2(new_n153_), .A3(new_n61_), .ZN(new_n157_));
  AOI21_X1  g099(.A(new_n126_), .B1(new_n152_), .B2(new_n157_), .ZN(new_n158_));
  INV_X1    g100(.A(G217), .ZN(new_n159_));
  NOR3_X1   g101(.A1(new_n159_), .A2(new_n124_), .A3(G953), .ZN(new_n160_));
  NOR2_X1   g102(.A1(new_n64_), .A2(G143), .ZN(RLL_wire_A_13));
  XNOR2_X1 RLL_XNOR_13 (.A(RLL_wire_A_13), .B(KEYINPUT13), .ZN(new_n161_) );
  NOR2_X1   g103(.A1(new_n67_), .A2(G128), .ZN(new_n162_));
  OAI21_X1  g104(.A(G134), .B1(new_n161_), .B2(new_n162_), .ZN(new_n163_));
  NAND2_X1  g105(.A1(new_n67_), .A2(G128), .ZN(new_n164_));
  NAND2_X1  g106(.A1(new_n64_), .A2(G143), .ZN(new_n165_));
  NAND3_X1  g107(.A1(new_n164_), .A2(new_n165_), .A3(new_n135_), .ZN(new_n166_));
  INV_X1    g108(.A(G122), .ZN(new_n167_));
  NAND2_X1  g109(.A1(new_n167_), .A2(G116), .ZN(new_n168_));
  NAND2_X1  g110(.A1(new_n85_), .A2(G122), .ZN(new_n169_));
  AND3_X1   g111(.A1(new_n168_), .A2(new_n169_), .A3(new_n91_), .ZN(new_n170_));
  AOI21_X1  g112(.A(new_n91_), .B1(new_n168_), .B2(new_n169_), .ZN(new_n171_));
  OAI211_X1 g113(.A(new_n166_), .B(new_n163_), .C1(new_n170_), .C2(new_n171_), .ZN(new_n172_));
  AOI21_X1  g114(.A(new_n135_), .B1(new_n164_), .B2(new_n165_), .ZN(new_n173_));
  AND3_X1   g115(.A1(new_n164_), .A2(new_n165_), .A3(new_n135_), .ZN(new_n174_));
  NAND3_X1  g116(.A1(new_n168_), .A2(new_n169_), .A3(new_n91_), .ZN(new_n175_));
  NOR2_X1   g117(.A1(new_n85_), .A2(G122), .ZN(new_n176_));
  NOR2_X1   g118(.A1(new_n167_), .A2(G116), .ZN(RLL_wire_A_14));
  XOR2_X1 RLL_XOR_14 (.A(RLL_wire_A_14), .B(KEYINPUT14), .Z(new_n177_) );
  OAI21_X1  g119(.A(G107), .B1(new_n176_), .B2(new_n177_), .ZN(new_n178_));
  OAI211_X1 g120(.A(new_n175_), .B(new_n178_), .C1(new_n174_), .C2(new_n173_), .ZN(new_n179_));
  AND3_X1   g121(.A1(new_n172_), .A2(new_n179_), .A3(new_n160_), .ZN(new_n180_));
  AOI21_X1  g122(.A(new_n160_), .B1(new_n172_), .B2(new_n179_), .ZN(new_n181_));
  OAI21_X1  g123(.A(new_n61_), .B1(new_n180_), .B2(new_n181_), .ZN(RLL_wire_A_15));
  XOR2_X1 RLL_XOR_15 (.A(RLL_wire_A_15), .B(KEYINPUT15), .Z(new_n182_) );
  NAND2_X1  g124(.A1(new_n182_), .A2(G478), .ZN(new_n183_));
  INV_X1    g125(.A(G478), .ZN(new_n184_));
  OAI211_X1 g126(.A(new_n184_), .B(new_n61_), .C1(new_n180_), .C2(new_n181_), .ZN(new_n185_));
  NAND2_X1  g127(.A1(new_n183_), .A2(new_n185_), .ZN(new_n186_));
  INV_X1    g128(.A(G475), .ZN(new_n187_));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n188_));
  XNOR2_X1  g130(.A(new_n188_), .B(new_n93_), .ZN(new_n189_));
  NAND2_X1  g131(.A1(new_n72_), .A2(G140), .ZN(new_n190_));
  INV_X1    g132(.A(G140), .ZN(new_n191_));
  NAND2_X1  g133(.A1(new_n191_), .A2(G125), .ZN(RLL_wire_A_16));
  XNOR2_X1 RLL_XNOR_16 (.A(RLL_wire_A_16), .B(KEYINPUT16), .ZN(new_n192_) );
  AND3_X1   g134(.A1(new_n190_), .A2(new_n192_), .A3(new_n65_), .ZN(new_n193_));
  AOI21_X1  g135(.A(new_n65_), .B1(new_n190_), .B2(new_n192_), .ZN(new_n194_));
  NOR2_X1   g136(.A1(new_n193_), .A2(new_n194_), .ZN(new_n195_));
  INV_X1    g137(.A(G237), .ZN(new_n196_));
  NAND4_X1  g138(.A1(new_n196_), .A2(new_n128_), .A3(G143), .A4(G214), .ZN(new_n197_));
  INV_X1    g139(.A(G214), .ZN(new_n198_));
  NOR3_X1   g140(.A1(new_n198_), .A2(G237), .A3(G953), .ZN(new_n199_));
  OAI211_X1 g141(.A(new_n132_), .B(new_n197_), .C1(new_n199_), .C2(G143), .ZN(new_n200_));
  INV_X1    g142(.A(new_n200_), .ZN(new_n201_));
  NAND3_X1  g143(.A1(new_n196_), .A2(new_n128_), .A3(G214), .ZN(new_n202_));
  NAND2_X1  g144(.A1(new_n202_), .A2(new_n67_), .ZN(new_n203_));
  AOI21_X1  g145(.A(new_n132_), .B1(new_n203_), .B2(new_n197_), .ZN(RLL_wire_A_17));
  XOR2_X1 RLL_XOR_17 (.A(RLL_wire_A_17), .B(KEYINPUT17), .Z(new_n204_) );
  OAI21_X1  g146(.A(new_n195_), .B1(new_n201_), .B2(new_n204_), .ZN(new_n205_));
  NOR3_X1   g147(.A1(new_n198_), .A2(G237), .A3(G953), .ZN(new_n206_));
  OAI21_X1  g148(.A(new_n197_), .B1(new_n206_), .B2(G143), .ZN(RLL_wire_A_18));
  XNOR2_X1 RLL_XNOR_18 (.A(RLL_wire_A_18), .B(KEYINPUT18), .ZN(new_n207_) );
  NAND2_X1  g149(.A1(new_n207_), .A2(G131), .ZN(new_n208_));
  XNOR2_X1  g150(.A(G125), .B(G140), .ZN(new_n209_));
  AND2_X1   g151(.A1(G125), .A2(G140), .ZN(new_n210_));
  NOR2_X1   g152(.A1(G125), .A2(G140), .ZN(new_n211_));
  OAI21_X1  g153(.A(new_n65_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g154(.A(new_n212_), .B1(new_n209_), .B2(new_n65_), .ZN(new_n213_));
  NAND3_X1  g155(.A1(new_n208_), .A2(new_n200_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g156(.A1(new_n205_), .A2(new_n189_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g157(.A(new_n189_), .ZN(new_n216_));
  NAND2_X1  g158(.A1(new_n205_), .A2(new_n214_), .ZN(new_n217_));
  NAND2_X1  g159(.A1(new_n217_), .A2(new_n216_), .ZN(new_n218_));
  AOI21_X1  g160(.A(G902), .B1(new_n218_), .B2(new_n215_), .ZN(new_n219_));
  AND3_X1   g161(.A1(new_n205_), .A2(new_n189_), .A3(new_n214_), .ZN(new_n220_));
  NAND3_X1  g162(.A1(new_n196_), .A2(new_n128_), .A3(G214), .ZN(new_n221_));
  NAND2_X1  g163(.A1(new_n221_), .A2(new_n67_), .ZN(new_n222_));
  AOI21_X1  g164(.A(new_n132_), .B1(new_n222_), .B2(new_n197_), .ZN(new_n223_));
  OR2_X1    g165(.A1(new_n210_), .A2(new_n211_), .ZN(RLL_wire_A_19));
  XNOR2_X1 RLL_XNOR_19 (.A(RLL_wire_A_19), .B(KEYINPUT19), .ZN(new_n224_) );
  AOI21_X1  g166(.A(new_n194_), .B1(new_n65_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g167(.A(new_n225_), .B1(new_n201_), .B2(new_n223_), .ZN(new_n226_));
  AOI21_X1  g168(.A(new_n189_), .B1(new_n226_), .B2(new_n214_), .ZN(new_n227_));
  OAI211_X1 g169(.A(new_n187_), .B(new_n61_), .C1(new_n220_), .C2(new_n227_), .ZN(RLL_wire_A_20));
  XNOR2_X1 RLL_XNOR_20 (.A(RLL_wire_A_20), .B(KEYINPUT20), .ZN(new_n228_) );
  OAI21_X1  g170(.A(new_n228_), .B1(new_n219_), .B2(new_n187_), .ZN(new_n229_));
  INV_X1    g171(.A(G898), .ZN(RLL_wire_A_21));
  XOR2_X1 RLL_XOR_21 (.A(RLL_wire_A_21), .B(KEYINPUT21), .Z(new_n230_) );
  NAND2_X1  g172(.A1(G234), .A2(G237), .ZN(new_n231_));
  NAND4_X1  g173(.A1(new_n231_), .A2(new_n230_), .A3(G902), .A4(G953), .ZN(new_n232_));
  NAND3_X1  g174(.A1(new_n231_), .A2(G952), .A3(new_n128_), .ZN(new_n233_));
  NAND2_X1  g175(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g176(.A(new_n234_), .ZN(new_n235_));
  NOR3_X1   g177(.A1(new_n229_), .A2(new_n186_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g178(.A1(new_n128_), .A2(G221), .A3(G234), .ZN(new_n237_));
  XNOR2_X1  g179(.A(new_n237_), .B(new_n133_), .ZN(RLL_wire_A_22));
  XOR2_X1 RLL_XOR_22 (.A(RLL_wire_A_22), .B(KEYINPUT22), .Z(new_n238_) );
  INV_X1    g180(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g181(.A(new_n194_), .ZN(new_n240_));
  NOR2_X1   g182(.A1(new_n83_), .A2(G128), .ZN(RLL_wire_A_23));
  XNOR2_X1 RLL_XNOR_23 (.A(RLL_wire_A_23), .B(KEYINPUT23), .ZN(new_n241_) );
  NOR2_X1   g183(.A1(new_n64_), .A2(G119), .ZN(new_n242_));
  NOR3_X1   g184(.A1(new_n241_), .A2(new_n242_), .A3(G110), .ZN(new_n243_));
  INV_X1    g185(.A(G110), .ZN(RLL_wire_A_24));
  XNOR2_X1 RLL_XNOR_24 (.A(RLL_wire_A_24), .B(KEYINPUT24), .ZN(new_n244_) );
  XNOR2_X1  g186(.A(G119), .B(G128), .ZN(new_n245_));
  NOR2_X1   g187(.A1(new_n245_), .A2(new_n244_), .ZN(new_n246_));
  OAI211_X1 g188(.A(new_n240_), .B(new_n212_), .C1(new_n246_), .C2(new_n243_), .ZN(new_n247_));
  NAND2_X1  g189(.A1(new_n245_), .A2(new_n244_), .ZN(new_n248_));
  OAI21_X1  g190(.A(G110), .B1(new_n241_), .B2(new_n242_), .ZN(new_n249_));
  OAI211_X1 g191(.A(new_n248_), .B(new_n249_), .C1(new_n193_), .C2(new_n194_), .ZN(new_n250_));
  AND3_X1   g192(.A1(new_n247_), .A2(new_n239_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g193(.A(new_n239_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n252_));
  OAI21_X1  g194(.A(new_n61_), .B1(new_n251_), .B2(new_n252_), .ZN(RLL_wire_A_25));
  XOR2_X1 RLL_XOR_25 (.A(RLL_wire_A_25), .B(KEYINPUT25), .Z(new_n253_) );
  AOI21_X1  g195(.A(new_n159_), .B1(G234), .B2(new_n61_), .ZN(new_n254_));
  NAND2_X1  g196(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g197(.A(new_n254_), .ZN(new_n256_));
  OAI211_X1 g198(.A(new_n61_), .B(new_n256_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g199(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g200(.A1(new_n196_), .A2(new_n128_), .A3(G210), .ZN(RLL_wire_A_26));
  XOR2_X1 RLL_XOR_26 (.A(RLL_wire_A_26), .B(KEYINPUT26), .Z(new_n259_) );
  XNOR2_X1  g201(.A(new_n259_), .B(new_n90_), .ZN(RLL_wire_A_27));
  XNOR2_X1 RLL_XNOR_27 (.A(RLL_wire_A_27), .B(KEYINPUT27), .ZN(new_n260_) );
  INV_X1    g202(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g203(.A1(new_n88_), .A2(new_n89_), .ZN(new_n262_));
  NOR2_X1   g204(.A1(new_n135_), .A2(G137), .ZN(new_n263_));
  NOR2_X1   g205(.A1(new_n133_), .A2(G134), .ZN(new_n264_));
  OAI21_X1  g206(.A(G131), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g207(.A1(new_n134_), .A2(new_n136_), .A3(new_n132_), .ZN(new_n266_));
  NAND4_X1  g208(.A1(new_n76_), .A2(new_n265_), .A3(new_n73_), .A4(new_n266_), .ZN(new_n267_));
  OAI22_X1  g209(.A1(new_n69_), .A2(new_n70_), .B1(new_n138_), .B2(new_n137_), .ZN(new_n268_));
  AND3_X1   g210(.A1(new_n268_), .A2(new_n267_), .A3(new_n262_), .ZN(RLL_wire_A_28));
  XNOR2_X1 RLL_XNOR_28 (.A(RLL_wire_A_28), .B(KEYINPUT28), .ZN(new_n269_) );
  AOI21_X1  g211(.A(new_n262_), .B1(new_n268_), .B2(new_n267_), .ZN(new_n270_));
  NOR3_X1   g212(.A1(new_n269_), .A2(new_n270_), .A3(new_n261_), .ZN(RLL_wire_A_29));
  XOR2_X1 RLL_XOR_29 (.A(RLL_wire_A_29), .B(KEYINPUT29), .Z(new_n271_) );
  INV_X1    g213(.A(new_n262_), .ZN(new_n272_));
  NAND2_X1  g214(.A1(new_n268_), .A2(new_n267_), .ZN(RLL_wire_A_30));
  XNOR2_X1 RLL_XNOR_30 (.A(RLL_wire_A_30), .B(KEYINPUT30), .ZN(new_n273_) );
  NAND2_X1  g215(.A1(new_n273_), .A2(new_n272_), .ZN(new_n274_));
  NAND3_X1  g216(.A1(new_n268_), .A2(new_n267_), .A3(new_n262_), .ZN(new_n275_));
  AOI21_X1  g217(.A(new_n260_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g218(.A(new_n61_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g219(.A1(new_n277_), .A2(G472), .ZN(new_n278_));
  INV_X1    g220(.A(G472), .ZN(new_n279_));
  OAI21_X1  g221(.A(new_n261_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n280_));
  NAND3_X1  g222(.A1(new_n274_), .A2(new_n260_), .A3(new_n275_), .ZN(RLL_wire_A_31));
  XOR2_X1 RLL_XOR_31 (.A(RLL_wire_A_31), .B(KEYINPUT31), .Z(new_n281_) );
  NAND2_X1  g223(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g224(.A1(new_n282_), .A2(new_n279_), .A3(new_n61_), .ZN(RLL_wire_A_32));
  XNOR2_X1 RLL_XNOR_32 (.A(RLL_wire_A_32), .B(KEYINPUT32), .ZN(new_n283_) );
  AOI21_X1  g225(.A(new_n258_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g226(.A1(new_n284_), .A2(new_n158_), .A3(new_n236_), .A4(new_n123_), .ZN(new_n285_));
  XNOR2_X1  g227(.A(new_n285_), .B(G101), .ZN(G3));
  NAND3_X1  g228(.A1(new_n172_), .A2(new_n179_), .A3(new_n160_), .ZN(new_n287_));
  INV_X1    g229(.A(new_n160_), .ZN(new_n288_));
  NAND2_X1  g230(.A1(new_n172_), .A2(new_n179_), .ZN(new_n289_));
  NAND2_X1  g231(.A1(new_n289_), .A2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g232(.A1(new_n290_), .A2(new_n287_), .ZN(RLL_wire_A_33));
  XNOR2_X1 RLL_XNOR_33 (.A(RLL_wire_A_33), .B(KEYINPUT33), .ZN(new_n291_) );
  AOI21_X1  g233(.A(new_n184_), .B1(new_n291_), .B2(new_n61_), .ZN(new_n292_));
  INV_X1    g234(.A(new_n185_), .ZN(new_n293_));
  NOR2_X1   g235(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND3_X1   g236(.A1(new_n229_), .A2(new_n294_), .A3(new_n234_), .ZN(new_n295_));
  AOI21_X1  g237(.A(new_n279_), .B1(new_n282_), .B2(new_n61_), .ZN(new_n296_));
  AOI211_X1 g238(.A(G472), .B(G902), .C1(new_n280_), .C2(new_n281_), .ZN(new_n297_));
  NOR3_X1   g239(.A1(new_n296_), .A2(new_n297_), .A3(new_n258_), .ZN(new_n298_));
  NAND4_X1  g240(.A1(new_n298_), .A2(new_n158_), .A3(new_n295_), .A4(new_n123_), .ZN(new_n299_));
  XNOR2_X1  g241(.A(new_n299_), .B(G104), .ZN(RLL_wire_A_34));
  XOR2_X1 RLL_XOR_34 (.A(RLL_wire_A_34), .B(KEYINPUT34), .Z(G6) );
  AOI21_X1  g242(.A(new_n189_), .B1(new_n205_), .B2(new_n214_), .ZN(new_n301_));
  OAI21_X1  g243(.A(new_n61_), .B1(new_n220_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g244(.A1(new_n302_), .A2(G475), .ZN(new_n303_));
  AND4_X1   g245(.A1(new_n186_), .A2(new_n303_), .A3(new_n228_), .A4(new_n234_), .ZN(new_n304_));
  NAND4_X1  g246(.A1(new_n298_), .A2(new_n158_), .A3(new_n123_), .A4(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g247(.A(new_n305_), .B(G107), .ZN(RLL_wire_A_35));
  XOR2_X1 RLL_XOR_35 (.A(RLL_wire_A_35), .B(KEYINPUT35), .Z(G9) );
  NAND3_X1  g248(.A1(new_n247_), .A2(new_n239_), .A3(new_n250_), .ZN(new_n307_));
  NAND2_X1  g249(.A1(new_n247_), .A2(new_n250_), .ZN(RLL_wire_A_36));
  XOR2_X1 RLL_XOR_36 (.A(RLL_wire_A_36), .B(KEYINPUT36), .Z(new_n308_) );
  NAND2_X1  g250(.A1(new_n308_), .A2(new_n238_), .ZN(new_n309_));
  AOI21_X1  g251(.A(new_n254_), .B1(new_n309_), .B2(new_n307_), .ZN(new_n310_));
  AOI22_X1  g252(.A1(new_n61_), .A2(new_n310_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n311_));
  NOR3_X1   g253(.A1(new_n296_), .A2(new_n297_), .A3(new_n311_), .ZN(new_n312_));
  NAND4_X1  g254(.A1(new_n312_), .A2(new_n158_), .A3(new_n123_), .A4(new_n236_), .ZN(new_n313_));
  XNOR2_X1  g255(.A(new_n313_), .B(G110), .ZN(RLL_wire_A_37));
  XOR2_X1 RLL_XOR_37 (.A(RLL_wire_A_37), .B(KEYINPUT37), .Z(G12) );
  INV_X1    g256(.A(G900), .ZN(new_n315_));
  NAND4_X1  g257(.A1(new_n231_), .A2(new_n315_), .A3(G902), .A4(G953), .ZN(new_n316_));
  NAND2_X1  g258(.A1(new_n316_), .A2(new_n233_), .ZN(new_n317_));
  AND4_X1   g259(.A1(new_n186_), .A2(new_n303_), .A3(new_n228_), .A4(new_n317_), .ZN(new_n318_));
  AOI21_X1  g260(.A(new_n311_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n319_));
  NAND4_X1  g261(.A1(new_n319_), .A2(new_n158_), .A3(new_n123_), .A4(new_n318_), .ZN(new_n320_));
  XNOR2_X1  g262(.A(new_n320_), .B(G128), .ZN(G30));
  AND2_X1   g263(.A1(new_n229_), .A2(new_n186_), .ZN(new_n322_));
  NAND2_X1  g264(.A1(new_n121_), .A2(new_n122_), .ZN(RLL_wire_A_38));
  XNOR2_X1 RLL_XNOR_38 (.A(RLL_wire_A_38), .B(KEYINPUT38), .ZN(new_n323_) );
  NAND3_X1  g265(.A1(new_n268_), .A2(new_n267_), .A3(new_n262_), .ZN(new_n324_));
  NAND3_X1  g266(.A1(new_n274_), .A2(new_n260_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g267(.A(new_n275_), .ZN(new_n326_));
  OAI21_X1  g268(.A(new_n261_), .B1(new_n326_), .B2(new_n270_), .ZN(new_n327_));
  AOI21_X1  g269(.A(G902), .B1(new_n327_), .B2(new_n325_), .ZN(new_n328_));
  OAI21_X1  g270(.A(new_n283_), .B1(new_n279_), .B2(new_n328_), .ZN(new_n329_));
  AND3_X1   g271(.A1(new_n329_), .A2(new_n323_), .A3(new_n59_), .ZN(new_n330_));
  INV_X1    g272(.A(new_n317_), .ZN(RLL_wire_A_39));
  XNOR2_X1 RLL_XNOR_39 (.A(RLL_wire_A_39), .B(KEYINPUT39), .ZN(new_n331_) );
  AOI211_X1 g273(.A(new_n126_), .B(new_n331_), .C1(new_n152_), .C2(new_n157_), .ZN(RLL_wire_A_40));
  XNOR2_X1 RLL_XNOR_40 (.A(RLL_wire_A_40), .B(KEYINPUT40), .ZN(new_n332_) );
  NAND4_X1  g274(.A1(new_n330_), .A2(new_n332_), .A3(new_n311_), .A4(new_n322_), .ZN(new_n333_));
  XNOR2_X1  g275(.A(new_n333_), .B(G143), .ZN(G45));
  AND3_X1   g276(.A1(new_n229_), .A2(new_n294_), .A3(new_n317_), .ZN(new_n335_));
  NAND4_X1  g277(.A1(new_n158_), .A2(new_n319_), .A3(new_n335_), .A4(new_n123_), .ZN(new_n336_));
  XNOR2_X1  g278(.A(new_n336_), .B(G146), .ZN(G48));
  AOI21_X1  g279(.A(new_n153_), .B1(new_n156_), .B2(new_n61_), .ZN(new_n338_));
  AOI211_X1 g280(.A(G469), .B(G902), .C1(new_n154_), .C2(new_n155_), .ZN(new_n339_));
  NOR3_X1   g281(.A1(new_n338_), .A2(new_n339_), .A3(new_n126_), .ZN(new_n340_));
  NAND4_X1  g282(.A1(new_n340_), .A2(new_n284_), .A3(new_n295_), .A4(new_n123_), .ZN(new_n341_));
  XNOR2_X1  g283(.A(new_n341_), .B(G113), .ZN(RLL_wire_A_41));
  XNOR2_X1 RLL_XNOR_41 (.A(RLL_wire_A_41), .B(KEYINPUT41), .ZN(G15) );
  NAND4_X1  g284(.A1(new_n340_), .A2(new_n284_), .A3(new_n123_), .A4(new_n304_), .ZN(new_n343_));
  XNOR2_X1  g285(.A(new_n343_), .B(G116), .ZN(G18));
  NAND4_X1  g286(.A1(new_n340_), .A2(new_n319_), .A3(new_n123_), .A4(new_n236_), .ZN(new_n345_));
  XNOR2_X1  g287(.A(new_n345_), .B(G119), .ZN(G21));
  AOI211_X1 g288(.A(new_n60_), .B(new_n235_), .C1(new_n121_), .C2(new_n122_), .ZN(new_n347_));
  NAND4_X1  g289(.A1(new_n347_), .A2(new_n298_), .A3(new_n322_), .A4(new_n340_), .ZN(new_n348_));
  XNOR2_X1  g290(.A(new_n348_), .B(G122), .ZN(G24));
  NAND4_X1  g291(.A1(new_n312_), .A2(new_n340_), .A3(new_n335_), .A4(new_n123_), .ZN(new_n350_));
  XNOR2_X1  g292(.A(new_n350_), .B(G125), .ZN(G27));
  AND3_X1   g293(.A1(new_n121_), .A2(new_n59_), .A3(new_n122_), .ZN(new_n352_));
  NAND4_X1  g294(.A1(new_n158_), .A2(new_n284_), .A3(new_n352_), .A4(new_n335_), .ZN(RLL_wire_A_42));
  XOR2_X1 RLL_XOR_42 (.A(RLL_wire_A_42), .B(KEYINPUT42), .Z(new_n353_) );
  XNOR2_X1  g295(.A(new_n353_), .B(G131), .ZN(G33));
  NAND4_X1  g296(.A1(new_n158_), .A2(new_n284_), .A3(new_n352_), .A4(new_n318_), .ZN(new_n355_));
  XNOR2_X1  g297(.A(new_n355_), .B(G134), .ZN(G36));
  NOR2_X1   g298(.A1(new_n296_), .A2(new_n297_), .ZN(new_n357_));
  NAND3_X1  g299(.A1(new_n294_), .A2(new_n303_), .A3(new_n228_), .ZN(RLL_wire_A_43));
  XNOR2_X1 RLL_XNOR_43 (.A(RLL_wire_A_43), .B(KEYINPUT43), .ZN(new_n358_) );
  NOR3_X1   g300(.A1(new_n357_), .A2(new_n358_), .A3(new_n311_), .ZN(RLL_wire_A_44));
  XOR2_X1 RLL_XOR_44 (.A(RLL_wire_A_44), .B(KEYINPUT44), .Z(new_n359_) );
  NAND3_X1  g301(.A1(new_n140_), .A2(new_n131_), .A3(new_n139_), .ZN(new_n360_));
  NAND2_X1  g302(.A1(new_n148_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g303(.A1(new_n142_), .A2(new_n130_), .ZN(new_n362_));
  AOI22_X1  g304(.A1(new_n361_), .A2(new_n130_), .B1(new_n362_), .B2(new_n149_), .ZN(RLL_wire_A_45));
  XOR2_X1 RLL_XOR_45 (.A(RLL_wire_A_45), .B(KEYINPUT45), .Z(new_n363_) );
  OAI21_X1  g305(.A(G469), .B1(new_n363_), .B2(G902), .ZN(RLL_wire_A_46));
  XOR2_X1 RLL_XOR_46 (.A(RLL_wire_A_46), .B(KEYINPUT46), .Z(new_n364_) );
  NAND3_X1  g306(.A1(new_n156_), .A2(new_n153_), .A3(new_n61_), .ZN(new_n365_));
  AOI211_X1 g307(.A(new_n126_), .B(new_n331_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g308(.A1(new_n359_), .A2(new_n352_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g309(.A(new_n367_), .B(G137), .ZN(G39));
  AOI21_X1  g310(.A(new_n126_), .B1(new_n364_), .B2(new_n365_), .ZN(RLL_wire_A_47));
  XNOR2_X1 RLL_XNOR_47 (.A(RLL_wire_A_47), .B(KEYINPUT47), .ZN(new_n369_) );
  AND3_X1   g311(.A1(new_n278_), .A2(new_n258_), .A3(new_n283_), .ZN(new_n370_));
  NAND4_X1  g312(.A1(new_n370_), .A2(new_n369_), .A3(new_n335_), .A4(new_n352_), .ZN(new_n371_));
  XNOR2_X1  g313(.A(new_n371_), .B(G140), .ZN(G42));
  NAND2_X1  g314(.A1(new_n229_), .A2(new_n294_), .ZN(new_n373_));
  INV_X1    g315(.A(new_n373_), .ZN(new_n374_));
  NOR3_X1   g316(.A1(new_n329_), .A2(new_n233_), .A3(new_n258_), .ZN(new_n375_));
  NAND4_X1  g317(.A1(new_n375_), .A2(new_n374_), .A3(new_n340_), .A4(new_n352_), .ZN(new_n376_));
  NOR2_X1   g318(.A1(new_n358_), .A2(new_n233_), .ZN(new_n377_));
  NAND4_X1  g319(.A1(new_n377_), .A2(new_n284_), .A3(new_n340_), .A4(new_n352_), .ZN(RLL_wire_A_48));
  XNOR2_X1 RLL_XNOR_48 (.A(RLL_wire_A_48), .B(KEYINPUT48), .ZN(new_n378_) );
  NAND2_X1  g320(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g321(.A1(new_n338_), .A2(new_n339_), .ZN(RLL_wire_A_49));
  XNOR2_X1 RLL_XNOR_49 (.A(RLL_wire_A_49), .B(KEYINPUT49), .ZN(new_n380_) );
  NOR3_X1   g322(.A1(new_n329_), .A2(new_n323_), .A3(new_n229_), .ZN(new_n381_));
  NAND3_X1  g323(.A1(new_n381_), .A2(new_n294_), .A3(new_n380_), .ZN(new_n382_));
  NOR4_X1   g324(.A1(new_n382_), .A2(new_n60_), .A3(new_n126_), .A4(new_n258_), .ZN(new_n383_));
  AND2_X1   g325(.A1(new_n377_), .A2(new_n298_), .ZN(new_n384_));
  NAND3_X1  g326(.A1(new_n384_), .A2(new_n123_), .A3(new_n340_), .ZN(new_n385_));
  NAND3_X1  g327(.A1(new_n385_), .A2(G952), .A3(new_n128_), .ZN(new_n386_));
  NAND4_X1  g328(.A1(new_n377_), .A2(new_n312_), .A3(new_n340_), .A4(new_n352_), .ZN(new_n387_));
  NOR2_X1   g329(.A1(new_n323_), .A2(new_n59_), .ZN(new_n388_));
  NAND3_X1  g330(.A1(new_n384_), .A2(new_n340_), .A3(new_n388_), .ZN(RLL_wire_A_50));
  XOR2_X1 RLL_XOR_50 (.A(RLL_wire_A_50), .B(KEYINPUT50), .Z(new_n389_) );
  NOR2_X1   g331(.A1(new_n229_), .A2(new_n294_), .ZN(new_n390_));
  NAND4_X1  g332(.A1(new_n375_), .A2(new_n340_), .A3(new_n352_), .A4(new_n390_), .ZN(new_n391_));
  NOR3_X1   g333(.A1(new_n338_), .A2(new_n339_), .A3(new_n125_), .ZN(new_n392_));
  OAI211_X1 g334(.A(new_n384_), .B(new_n352_), .C1(new_n369_), .C2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g335(.A1(new_n393_), .A2(new_n389_), .A3(new_n387_), .A4(new_n391_), .ZN(RLL_wire_A_51));
  XOR2_X1 RLL_XOR_51 (.A(RLL_wire_A_51), .B(KEYINPUT51), .Z(new_n394_) );
  NOR4_X1   g336(.A1(new_n394_), .A2(new_n386_), .A3(new_n383_), .A4(new_n379_), .ZN(new_n395_));
  AND4_X1   g337(.A1(new_n285_), .A2(new_n299_), .A3(new_n313_), .A4(new_n305_), .ZN(new_n396_));
  AND4_X1   g338(.A1(new_n341_), .A2(new_n348_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n397_));
  NAND2_X1  g339(.A1(new_n158_), .A2(new_n317_), .ZN(new_n398_));
  NAND2_X1  g340(.A1(new_n312_), .A2(new_n335_), .ZN(new_n399_));
  NAND2_X1  g341(.A1(new_n158_), .A2(new_n352_), .ZN(new_n400_));
  NOR2_X1   g342(.A1(new_n229_), .A2(new_n186_), .ZN(new_n401_));
  NAND3_X1  g343(.A1(new_n319_), .A2(new_n352_), .A3(new_n401_), .ZN(new_n402_));
  OAI22_X1  g344(.A1(new_n402_), .A2(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n403_));
  NAND2_X1  g345(.A1(new_n353_), .A2(new_n355_), .ZN(new_n404_));
  NOR2_X1   g346(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g347(.A1(new_n322_), .A2(new_n123_), .A3(new_n311_), .A4(new_n329_), .ZN(new_n406_));
  OAI21_X1  g348(.A(new_n320_), .B1(new_n406_), .B2(new_n398_), .ZN(new_n407_));
  NAND2_X1  g349(.A1(new_n350_), .A2(new_n336_), .ZN(new_n408_));
  NOR2_X1   g350(.A1(new_n407_), .A2(new_n408_), .ZN(RLL_wire_A_52));
  XNOR2_X1 RLL_XNOR_52 (.A(RLL_wire_A_52), .B(KEYINPUT52), .ZN(new_n409_) );
  NAND4_X1  g351(.A1(new_n405_), .A2(new_n409_), .A3(new_n397_), .A4(new_n396_), .ZN(RLL_wire_A_53));
  XOR2_X1 RLL_XOR_53 (.A(RLL_wire_A_53), .B(KEYINPUT53), .Z(new_n410_) );
  INV_X1    g352(.A(new_n410_), .ZN(RLL_wire_A_54));
  XNOR2_X1 RLL_XNOR_54 (.A(RLL_wire_A_54), .B(KEYINPUT54), .ZN(new_n411_) );
  NOR3_X1   g353(.A1(new_n383_), .A2(G952), .A3(G953), .ZN(new_n412_));
  AOI21_X1  g354(.A(new_n412_), .B1(new_n395_), .B2(new_n411_), .ZN(G75));
  NOR2_X1   g355(.A1(new_n128_), .A2(G952), .ZN(new_n414_));
  NOR2_X1   g356(.A1(new_n119_), .A2(new_n61_), .ZN(new_n415_));
  NOR2_X1   g357(.A1(new_n79_), .A2(new_n80_), .ZN(new_n416_));
  NOR2_X1   g358(.A1(new_n106_), .A2(new_n107_), .ZN(new_n417_));
  XNOR2_X1  g359(.A(new_n417_), .B(new_n416_), .ZN(RLL_wire_A_55));
  XOR2_X1 RLL_XOR_55 (.A(RLL_wire_A_55), .B(KEYINPUT55), .Z(new_n418_) );
  NAND3_X1  g360(.A1(new_n410_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g361(.A(new_n418_), .ZN(RLL_wire_A_56));
  XOR2_X1 RLL_XOR_56 (.A(RLL_wire_A_56), .B(KEYINPUT56), .Z(new_n420_) );
  NAND2_X1  g362(.A1(new_n410_), .A2(new_n415_), .ZN(new_n421_));
  NAND2_X1  g363(.A1(new_n421_), .A2(new_n420_), .ZN(new_n422_));
  AOI21_X1  g364(.A(new_n414_), .B1(new_n422_), .B2(new_n419_), .ZN(G51));
  NAND4_X1  g365(.A1(new_n410_), .A2(G469), .A3(G902), .A4(new_n363_), .ZN(new_n424_));
  NAND2_X1  g366(.A1(G469), .A2(G902), .ZN(RLL_wire_A_57));
  XNOR2_X1 RLL_XNOR_57 (.A(RLL_wire_A_57), .B(KEYINPUT57), .ZN(new_n425_) );
  OAI21_X1  g367(.A(new_n156_), .B1(new_n411_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g368(.A(new_n414_), .B1(new_n426_), .B2(new_n424_), .ZN(G54));
  NOR2_X1   g369(.A1(new_n220_), .A2(new_n227_), .ZN(RLL_wire_A_58));
  XNOR2_X1 RLL_XNOR_58 (.A(RLL_wire_A_58), .B(KEYINPUT58), .ZN(new_n428_) );
  NAND4_X1  g370(.A1(new_n410_), .A2(G475), .A3(G902), .A4(new_n428_), .ZN(new_n429_));
  NAND3_X1  g371(.A1(new_n410_), .A2(G475), .A3(G902), .ZN(new_n430_));
  OAI21_X1  g372(.A(new_n430_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n431_));
  AOI21_X1  g373(.A(new_n414_), .B1(new_n431_), .B2(new_n429_), .ZN(G60));
  NAND2_X1  g374(.A1(G478), .A2(G902), .ZN(RLL_wire_A_59));
  XOR2_X1 RLL_XOR_59 (.A(RLL_wire_A_59), .B(KEYINPUT59), .Z(new_n433_) );
  OR3_X1    g375(.A1(new_n411_), .A2(new_n291_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g376(.A(new_n291_), .B1(new_n411_), .B2(new_n433_), .ZN(new_n435_));
  AOI21_X1  g377(.A(new_n414_), .B1(new_n434_), .B2(new_n435_), .ZN(G63));
  NOR2_X1   g378(.A1(new_n256_), .A2(new_n61_), .ZN(RLL_wire_A_60));
  XNOR2_X1 RLL_XNOR_60 (.A(RLL_wire_A_60), .B(KEYINPUT60), .ZN(new_n437_) );
  NAND4_X1  g379(.A1(new_n410_), .A2(new_n307_), .A3(new_n309_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g380(.A1(new_n410_), .A2(new_n437_), .ZN(new_n439_));
  OAI21_X1  g381(.A(new_n439_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n440_));
  AOI21_X1  g382(.A(new_n414_), .B1(new_n440_), .B2(new_n438_), .ZN(RLL_wire_A_61));
  XNOR2_X1 RLL_XNOR_61 (.A(RLL_wire_A_61), .B(KEYINPUT61), .ZN(G66) );
  OAI21_X1  g383(.A(new_n417_), .B1(G898), .B2(new_n128_), .ZN(new_n442_));
  NAND4_X1  g384(.A1(new_n348_), .A2(new_n341_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n443_));
  NAND4_X1  g385(.A1(new_n299_), .A2(new_n313_), .A3(new_n305_), .A4(new_n285_), .ZN(new_n444_));
  NOR2_X1   g386(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g387(.A1(new_n445_), .A2(G953), .ZN(new_n446_));
  NAND2_X1  g388(.A1(new_n446_), .A2(new_n442_), .ZN(new_n447_));
  INV_X1    g389(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g390(.A1(new_n446_), .A2(new_n442_), .ZN(new_n449_));
  OAI21_X1  g391(.A(G953), .B1(new_n62_), .B2(new_n230_), .ZN(new_n450_));
  OAI21_X1  g392(.A(new_n450_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n451_));
  OAI211_X1 g393(.A(new_n442_), .B(G953), .C1(new_n62_), .C2(new_n230_), .ZN(new_n452_));
  NAND2_X1  g394(.A1(new_n451_), .A2(new_n452_), .ZN(G69));
  INV_X1    g395(.A(new_n273_), .ZN(new_n454_));
  NOR2_X1   g396(.A1(new_n454_), .A2(new_n224_), .ZN(new_n455_));
  NAND2_X1  g397(.A1(new_n454_), .A2(new_n224_), .ZN(new_n456_));
  INV_X1    g398(.A(new_n456_), .ZN(new_n457_));
  AOI211_X1 g399(.A(new_n455_), .B(new_n457_), .C1(new_n315_), .C2(G953), .ZN(new_n458_));
  NAND4_X1  g400(.A1(new_n367_), .A2(new_n353_), .A3(new_n355_), .A4(new_n371_), .ZN(new_n459_));
  NAND4_X1  g401(.A1(new_n366_), .A2(new_n123_), .A3(new_n284_), .A4(new_n322_), .ZN(new_n460_));
  NAND4_X1  g402(.A1(new_n460_), .A2(new_n320_), .A3(new_n336_), .A4(new_n350_), .ZN(new_n461_));
  NOR2_X1   g403(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g404(.A(new_n458_), .B1(new_n462_), .B2(G953), .ZN(new_n463_));
  INV_X1    g405(.A(new_n458_), .ZN(new_n464_));
  NAND4_X1  g406(.A1(new_n333_), .A2(new_n320_), .A3(new_n336_), .A4(new_n350_), .ZN(RLL_wire_A_62));
  XNOR2_X1 RLL_XNOR_62 (.A(RLL_wire_A_62), .B(KEYINPUT62), .ZN(new_n465_) );
  NAND2_X1  g407(.A1(new_n367_), .A2(new_n371_), .ZN(new_n466_));
  NAND3_X1  g408(.A1(new_n186_), .A2(new_n303_), .A3(new_n228_), .ZN(new_n467_));
  AOI21_X1  g409(.A(new_n331_), .B1(new_n373_), .B2(new_n467_), .ZN(new_n468_));
  AND4_X1   g410(.A1(new_n158_), .A2(new_n468_), .A3(new_n284_), .A4(new_n352_), .ZN(new_n469_));
  OR3_X1    g411(.A1(new_n465_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g412(.A1(new_n470_), .A2(new_n128_), .A3(new_n464_), .ZN(new_n471_));
  NAND2_X1  g413(.A1(new_n471_), .A2(new_n463_), .ZN(new_n472_));
  AOI21_X1  g414(.A(new_n128_), .B1(G227), .B2(G900), .ZN(new_n473_));
  INV_X1    g415(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g416(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g417(.A1(new_n471_), .A2(new_n463_), .A3(new_n473_), .ZN(new_n476_));
  NAND2_X1  g418(.A1(new_n475_), .A2(new_n476_), .ZN(G72));
  NAND2_X1  g419(.A1(new_n274_), .A2(new_n324_), .ZN(new_n478_));
  NOR2_X1   g420(.A1(new_n279_), .A2(new_n61_), .ZN(RLL_wire_A_63));
  XNOR2_X1 RLL_XNOR_63 (.A(RLL_wire_A_63), .B(KEYINPUT63), .ZN(new_n479_) );
  INV_X1    g421(.A(new_n479_), .ZN(new_n480_));
  AOI211_X1 g422(.A(new_n478_), .B(new_n480_), .C1(new_n462_), .C2(new_n445_), .ZN(new_n481_));
  INV_X1    g423(.A(new_n478_), .ZN(new_n482_));
  AOI21_X1  g424(.A(new_n482_), .B1(new_n410_), .B2(new_n479_), .ZN(new_n483_));
  OAI21_X1  g425(.A(new_n261_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g426(.A1(new_n410_), .A2(new_n482_), .A3(new_n479_), .ZN(new_n485_));
  NOR3_X1   g427(.A1(new_n465_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n486_));
  NAND4_X1  g428(.A1(new_n299_), .A2(new_n313_), .A3(new_n305_), .A4(new_n285_), .ZN(new_n487_));
  NAND4_X1  g429(.A1(new_n348_), .A2(new_n341_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n488_));
  NOR2_X1   g430(.A1(new_n488_), .A2(new_n487_), .ZN(new_n489_));
  AOI21_X1  g431(.A(new_n480_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g432(.A(new_n260_), .B(new_n485_), .C1(new_n490_), .C2(new_n482_), .ZN(new_n491_));
  AOI21_X1  g433(.A(new_n414_), .B1(new_n484_), .B2(new_n491_), .ZN(G57));

endmodule
