

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596;

  INV_X1 U325 ( .A(n498), .ZN(n539) );
  XOR2_X1 U326 ( .A(n404), .B(n403), .Z(n498) );
  NOR2_X1 U327 ( .A1(n539), .A2(n542), .ZN(n480) );
  NOR2_X2 U328 ( .A1(n589), .A2(n593), .ZN(n590) );
  OR2_X1 U329 ( .A1(n468), .A2(n566), .ZN(n462) );
  XNOR2_X1 U330 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n307) );
  XNOR2_X1 U331 ( .A(n368), .B(n332), .ZN(n333) );
  XOR2_X1 U332 ( .A(n355), .B(KEYINPUT67), .Z(n293) );
  XOR2_X1 U333 ( .A(G197GAT), .B(KEYINPUT123), .Z(n294) );
  XNOR2_X1 U334 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U335 ( .A(n319), .B(n318), .ZN(n325) );
  XNOR2_X1 U336 ( .A(n383), .B(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U337 ( .A(n469), .B(KEYINPUT118), .ZN(n470) );
  XNOR2_X1 U338 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U339 ( .A(n465), .B(n294), .ZN(n466) );
  XNOR2_X1 U340 ( .A(n467), .B(n466), .ZN(G1352GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n296) );
  NAND2_X1 U342 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U344 ( .A(n297), .B(KEYINPUT30), .Z(n305) );
  XOR2_X1 U345 ( .A(G113GAT), .B(G50GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(G36GAT), .B(G43GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U348 ( .A(KEYINPUT29), .B(G8GAT), .Z(n301) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(G197GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G1GAT), .Z(n344) );
  XOR2_X1 U354 ( .A(n306), .B(n344), .Z(n310) );
  XNOR2_X1 U355 ( .A(n307), .B(KEYINPUT8), .ZN(n313) );
  BUF_X1 U356 ( .A(n313), .Z(n308) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G22GAT), .Z(n454) );
  XNOR2_X1 U358 ( .A(n308), .B(n454), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n578) );
  XOR2_X1 U360 ( .A(G43GAT), .B(G134GAT), .Z(n436) );
  INV_X1 U361 ( .A(n313), .ZN(n311) );
  NAND2_X1 U362 ( .A1(n436), .A2(n311), .ZN(n315) );
  INV_X1 U363 ( .A(n436), .ZN(n312) );
  NAND2_X1 U364 ( .A1(n313), .A2(n312), .ZN(n314) );
  NAND2_X1 U365 ( .A1(n315), .A2(n314), .ZN(n319) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  INV_X1 U367 ( .A(KEYINPUT11), .ZN(n316) );
  INV_X1 U368 ( .A(n325), .ZN(n323) );
  XOR2_X1 U369 ( .A(G92GAT), .B(G218GAT), .Z(n321) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n392) );
  XNOR2_X1 U372 ( .A(n392), .B(KEYINPUT68), .ZN(n324) );
  INV_X1 U373 ( .A(n324), .ZN(n322) );
  NAND2_X1 U374 ( .A1(n323), .A2(n322), .ZN(n327) );
  NAND2_X1 U375 ( .A1(n325), .A2(n324), .ZN(n326) );
  NAND2_X1 U376 ( .A1(n327), .A2(n326), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n328), .B(KEYINPUT9), .ZN(n334) );
  XOR2_X1 U378 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n330) );
  XNOR2_X1 U379 ( .A(G106GAT), .B(G85GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U381 ( .A(G99GAT), .B(n331), .Z(n368) );
  XOR2_X1 U382 ( .A(G50GAT), .B(G162GAT), .Z(n448) );
  XOR2_X1 U383 ( .A(n448), .B(KEYINPUT10), .Z(n332) );
  XNOR2_X2 U384 ( .A(n334), .B(n333), .ZN(n576) );
  XNOR2_X2 U385 ( .A(KEYINPUT76), .B(n576), .ZN(n562) );
  XNOR2_X1 U386 ( .A(KEYINPUT36), .B(n562), .ZN(n592) );
  XOR2_X1 U387 ( .A(G127GAT), .B(G71GAT), .Z(n336) );
  XNOR2_X1 U388 ( .A(G22GAT), .B(G183GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U390 ( .A(G64GAT), .B(G78GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G211GAT), .B(G155GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U393 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U394 ( .A(G57GAT), .B(KEYINPUT13), .Z(n363) );
  XOR2_X1 U395 ( .A(G8GAT), .B(KEYINPUT77), .Z(n396) );
  XOR2_X1 U396 ( .A(n363), .B(n396), .Z(n342) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n354) );
  XOR2_X1 U401 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X1 U402 ( .A(KEYINPUT82), .B(KEYINPUT14), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n350) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n352), .B(n351), .Z(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n490) );
  INV_X1 U409 ( .A(n490), .ZN(n589) );
  NOR2_X1 U410 ( .A1(n592), .A2(n589), .ZN(n356) );
  XNOR2_X1 U411 ( .A(KEYINPUT45), .B(KEYINPUT108), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n293), .ZN(n371) );
  XOR2_X1 U413 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n362) );
  XNOR2_X1 U414 ( .A(G78GAT), .B(KEYINPUT71), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n357), .B(G148GAT), .ZN(n450) );
  XOR2_X1 U416 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n359) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(G92GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n450), .B(n360), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U421 ( .A(G204GAT), .B(G64GAT), .Z(n388) );
  XOR2_X1 U422 ( .A(n388), .B(n363), .Z(n365) );
  NAND2_X1 U423 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U425 ( .A(n367), .B(n366), .Z(n370) );
  XOR2_X1 U426 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U427 ( .A(n434), .B(n368), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n586) );
  NAND2_X1 U429 ( .A1(n371), .A2(n586), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n372), .B(KEYINPUT109), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n373), .A2(n578), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n374), .B(KEYINPUT110), .ZN(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT107), .B(KEYINPUT47), .Z(n380) );
  XNOR2_X1 U434 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n586), .B(n375), .ZN(n580) );
  NOR2_X1 U436 ( .A1(n578), .A2(n580), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n376), .B(KEYINPUT46), .ZN(n377) );
  NOR2_X1 U438 ( .A1(n490), .A2(n377), .ZN(n378) );
  NAND2_X1 U439 ( .A1(n378), .A2(n576), .ZN(n379) );
  XOR2_X1 U440 ( .A(n380), .B(n379), .Z(n381) );
  AND2_X1 U441 ( .A1(n382), .A2(n381), .ZN(n385) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT111), .Z(n383) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n548) );
  XOR2_X1 U444 ( .A(G211GAT), .B(KEYINPUT21), .Z(n387) );
  XNOR2_X1 U445 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n445) );
  XOR2_X1 U447 ( .A(n388), .B(n445), .Z(n390) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U450 ( .A(n391), .B(KEYINPUT92), .Z(n394) );
  XNOR2_X1 U451 ( .A(n392), .B(KEYINPUT93), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U453 ( .A(n395), .B(KEYINPUT91), .Z(n398) );
  XNOR2_X1 U454 ( .A(n396), .B(KEYINPUT94), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n404) );
  XNOR2_X1 U456 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n399), .B(KEYINPUT17), .ZN(n400) );
  XOR2_X1 U458 ( .A(n400), .B(KEYINPUT18), .Z(n402) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(G176GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n437) );
  INV_X1 U461 ( .A(n437), .ZN(n403) );
  XOR2_X1 U462 ( .A(KEYINPUT117), .B(n539), .Z(n405) );
  NOR2_X1 U463 ( .A1(n548), .A2(n405), .ZN(n406) );
  XNOR2_X1 U464 ( .A(KEYINPUT54), .B(n406), .ZN(n426) );
  XOR2_X1 U465 ( .A(KEYINPUT4), .B(G57GAT), .Z(n408) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G148GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n425) );
  XOR2_X1 U468 ( .A(G162GAT), .B(G120GAT), .Z(n410) );
  XNOR2_X1 U469 ( .A(G141GAT), .B(G134GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U471 ( .A(G29GAT), .B(G85GAT), .Z(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n421) );
  XNOR2_X1 U473 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n413), .B(KEYINPUT1), .ZN(n414) );
  XOR2_X1 U475 ( .A(n414), .B(KEYINPUT5), .Z(n419) );
  XOR2_X1 U476 ( .A(G127GAT), .B(KEYINPUT83), .Z(n416) );
  XNOR2_X1 U477 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n431) );
  XNOR2_X1 U479 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n417), .B(KEYINPUT2), .ZN(n444) );
  XNOR2_X1 U481 ( .A(n431), .B(n444), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n423) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U486 ( .A(n425), .B(n424), .Z(n536) );
  AND2_X1 U487 ( .A1(n426), .A2(n536), .ZN(n428) );
  INV_X1 U488 ( .A(KEYINPUT66), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n468) );
  XOR2_X1 U490 ( .A(KEYINPUT84), .B(G99GAT), .Z(n430) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(G190GAT), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n441) );
  XOR2_X1 U493 ( .A(KEYINPUT20), .B(n431), .Z(n433) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n550) );
  INV_X1 U500 ( .A(n550), .ZN(n542) );
  XOR2_X1 U501 ( .A(KEYINPUT86), .B(KEYINPUT89), .Z(n443) );
  XNOR2_X1 U502 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n460) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n458) );
  XOR2_X1 U505 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n447) );
  XNOR2_X1 U506 ( .A(G218GAT), .B(G106GAT), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT23), .B(n450), .Z(n452) );
  NAND2_X1 U510 ( .A1(G228GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n460), .B(n459), .ZN(n481) );
  NAND2_X1 U516 ( .A1(n542), .A2(n481), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(n461), .ZN(n566) );
  XNOR2_X2 U518 ( .A(n462), .B(KEYINPUT122), .ZN(n593) );
  NOR2_X1 U519 ( .A1(n578), .A2(n593), .ZN(n467) );
  XOR2_X1 U520 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n464) );
  XNOR2_X1 U521 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n468), .A2(n481), .ZN(n471) );
  INV_X1 U524 ( .A(KEYINPUT55), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n472), .A2(n550), .ZN(n581) );
  NOR2_X1 U526 ( .A1(n581), .A2(n562), .ZN(n475) );
  XNOR2_X1 U527 ( .A(KEYINPUT121), .B(KEYINPUT58), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n473), .B(G190GAT), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  NOR2_X1 U530 ( .A1(n589), .A2(n581), .ZN(n478) );
  INV_X1 U531 ( .A(G183GAT), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT120), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n478), .B(n477), .ZN(G1350GAT) );
  XNOR2_X1 U534 ( .A(n539), .B(KEYINPUT27), .ZN(n484) );
  NOR2_X1 U535 ( .A1(n536), .A2(n484), .ZN(n569) );
  XOR2_X1 U536 ( .A(KEYINPUT28), .B(n481), .Z(n545) );
  NAND2_X1 U537 ( .A1(n569), .A2(n545), .ZN(n549) );
  XNOR2_X1 U538 ( .A(KEYINPUT85), .B(n542), .ZN(n479) );
  NOR2_X1 U539 ( .A1(n549), .A2(n479), .ZN(n489) );
  NOR2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT25), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(KEYINPUT95), .ZN(n486) );
  NOR2_X1 U543 ( .A1(n566), .A2(n484), .ZN(n485) );
  NOR2_X1 U544 ( .A1(n486), .A2(n485), .ZN(n487) );
  INV_X1 U545 ( .A(n536), .ZN(n495) );
  NOR2_X1 U546 ( .A1(n487), .A2(n495), .ZN(n488) );
  NOR2_X1 U547 ( .A1(n489), .A2(n488), .ZN(n509) );
  NAND2_X1 U548 ( .A1(n562), .A2(n490), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT16), .B(n491), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n509), .A2(n492), .ZN(n525) );
  INV_X1 U551 ( .A(n578), .ZN(n524) );
  NAND2_X1 U552 ( .A1(n524), .A2(n586), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT75), .ZN(n512) );
  NAND2_X1 U554 ( .A1(n525), .A2(n512), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT96), .B(n494), .Z(n504) );
  NAND2_X1 U556 ( .A1(n504), .A2(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(KEYINPUT34), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  XOR2_X1 U559 ( .A(G8GAT), .B(KEYINPUT97), .Z(n500) );
  NAND2_X1 U560 ( .A1(n504), .A2(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U563 ( .A1(n550), .A2(n504), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  INV_X1 U565 ( .A(n545), .ZN(n503) );
  NAND2_X1 U566 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(KEYINPUT98), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G22GAT), .B(n506), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n508) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n509), .A2(n592), .ZN(n510) );
  NAND2_X1 U573 ( .A1(n510), .A2(n589), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT37), .ZN(n535) );
  NAND2_X1 U575 ( .A1(n535), .A2(n512), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT38), .B(n513), .ZN(n522) );
  NOR2_X1 U577 ( .A1(n536), .A2(n522), .ZN(n514) );
  XOR2_X1 U578 ( .A(n515), .B(n514), .Z(n516) );
  XNOR2_X1 U579 ( .A(KEYINPUT99), .B(n516), .ZN(G1328GAT) );
  NOR2_X1 U580 ( .A1(n539), .A2(n522), .ZN(n517) );
  XOR2_X1 U581 ( .A(KEYINPUT102), .B(n517), .Z(n518) );
  XNOR2_X1 U582 ( .A(G36GAT), .B(n518), .ZN(G1329GAT) );
  NOR2_X1 U583 ( .A1(n522), .A2(n542), .ZN(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G43GAT), .B(n521), .ZN(G1330GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n545), .ZN(n523) );
  XOR2_X1 U588 ( .A(G50GAT), .B(n523), .Z(G1331GAT) );
  NOR2_X1 U589 ( .A1(n580), .A2(n524), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n525), .A2(n534), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n536), .A2(n531), .ZN(n527) );
  XNOR2_X1 U592 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(G57GAT), .B(n528), .Z(G1332GAT) );
  NOR2_X1 U595 ( .A1(n539), .A2(n531), .ZN(n529) );
  XOR2_X1 U596 ( .A(G64GAT), .B(n529), .Z(G1333GAT) );
  NOR2_X1 U597 ( .A1(n542), .A2(n531), .ZN(n530) );
  XOR2_X1 U598 ( .A(G71GAT), .B(n530), .Z(G1334GAT) );
  NOR2_X1 U599 ( .A1(n545), .A2(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1335GAT) );
  NAND2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n544) );
  NOR2_X1 U603 ( .A1(n536), .A2(n544), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G85GAT), .B(KEYINPUT105), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1336GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n544), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT106), .B(n540), .Z(n541) );
  XNOR2_X1 U608 ( .A(G92GAT), .B(n541), .ZN(G1337GAT) );
  NOR2_X1 U609 ( .A1(n542), .A2(n544), .ZN(n543) );
  XOR2_X1 U610 ( .A(G99GAT), .B(n543), .Z(G1338GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT44), .B(n546), .Z(n547) );
  XNOR2_X1 U613 ( .A(G106GAT), .B(n547), .ZN(G1339GAT) );
  XNOR2_X1 U614 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n554) );
  BUF_X1 U615 ( .A(n548), .Z(n567) );
  NOR2_X1 U616 ( .A1(n567), .A2(n549), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(KEYINPUT112), .ZN(n561) );
  NOR2_X1 U619 ( .A1(n578), .A2(n561), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G113GAT), .B(n555), .ZN(G1340GAT) );
  XNOR2_X1 U622 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n580), .A2(n561), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G120GAT), .B(n558), .Z(G1341GAT) );
  NOR2_X1 U626 ( .A1(n589), .A2(n561), .ZN(n559) );
  XOR2_X1 U627 ( .A(KEYINPUT50), .B(n559), .Z(n560) );
  XNOR2_X1 U628 ( .A(G127GAT), .B(n560), .ZN(G1342GAT) );
  XNOR2_X1 U629 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G134GAT), .B(n565), .ZN(G1343GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n575) );
  NOR2_X1 U635 ( .A1(n578), .A2(n575), .ZN(n570) );
  XOR2_X1 U636 ( .A(G141GAT), .B(n570), .Z(G1344GAT) );
  NOR2_X1 U637 ( .A1(n580), .A2(n575), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G148GAT), .B(n573), .ZN(G1345GAT) );
  NOR2_X1 U641 ( .A1(n589), .A2(n575), .ZN(n574) );
  XOR2_X1 U642 ( .A(G155GAT), .B(n574), .Z(G1346GAT) );
  NOR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(G162GAT), .B(n577), .Z(G1347GAT) );
  NOR2_X1 U645 ( .A1(n578), .A2(n581), .ZN(n579) );
  XOR2_X1 U646 ( .A(G169GAT), .B(n579), .Z(G1348GAT) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n583) );
  XNOR2_X1 U649 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1349GAT) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n586), .A2(n593), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT126), .B(n590), .Z(n591) );
  XNOR2_X1 U656 ( .A(G211GAT), .B(n591), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

