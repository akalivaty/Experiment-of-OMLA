//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n629, new_n631, new_n632, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g033(.A(G113), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n465), .B2(G125), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(G2105), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT68), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI22_X1  g046(.A1(new_n470), .A2(new_n471), .B1(new_n459), .B2(new_n460), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n462), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(new_n464), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n460), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G137), .B1(G101), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n468), .A2(new_n479), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n479), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(G136), .B2(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(G114), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G102), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n495), .B(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n477), .A2(new_n478), .A3(new_n464), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(G126), .A3(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(G138), .A3(new_n468), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n480), .A2(KEYINPUT71), .A3(G138), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n468), .A2(new_n465), .A3(G138), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G62), .ZN(new_n515));
  INV_X1    g090(.A(G75), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n513), .B2(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n511), .A2(new_n512), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT73), .B(G88), .Z(new_n525));
  AOI21_X1  g100(.A(new_n510), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(G51), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n511), .B2(new_n512), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT76), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n544));
  AND2_X1   g119(.A1(KEYINPUT5), .A2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(KEYINPUT5), .A2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n544), .B(new_n541), .C1(new_n547), .C2(new_n539), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n543), .A2(G651), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT77), .B(G90), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n524), .A2(new_n550), .B1(new_n526), .B2(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n521), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n526), .A2(G43), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  INV_X1    g132(.A(new_n523), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n513), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n547), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n526), .A2(G53), .ZN(new_n573));
  XOR2_X1   g148(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n524), .A2(G91), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n526), .A2(KEYINPUT78), .A3(KEYINPUT9), .A4(G53), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n572), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n524), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n526), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n584), .A2(KEYINPUT79), .A3(new_n521), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n584), .B2(new_n521), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n524), .A2(G86), .B1(new_n526), .B2(G48), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  INV_X1    g164(.A(G72), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n547), .A2(new_n589), .B1(new_n590), .B2(new_n510), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI221_X1 g168(.A(KEYINPUT80), .B1(new_n590), .B2(new_n510), .C1(new_n547), .C2(new_n589), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(G651), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n524), .A2(G85), .B1(new_n526), .B2(G47), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n595), .A2(KEYINPUT81), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT81), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT82), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n607), .A2(G79), .A3(G543), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(G66), .B1(new_n545), .B2(new_n546), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n521), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g186(.A(G54), .B(G543), .C1(new_n558), .C2(new_n557), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n511), .B2(new_n512), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n606), .A2(new_n608), .ZN(new_n617));
  OAI21_X1  g192(.A(G651), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n612), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n559), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n614), .A2(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n603), .B1(new_n602), .B2(new_n624), .ZN(G284));
  AOI21_X1  g200(.A(new_n603), .B1(new_n602), .B2(new_n624), .ZN(G321));
  MUX2_X1   g201(.A(G286), .B(G299), .S(new_n602), .Z(G297));
  MUX2_X1   g202(.A(G286), .B(G299), .S(new_n602), .Z(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n624), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n629), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(new_n602), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n602), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g208(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n634));
  XNOR2_X1  g209(.A(G323), .B(new_n634), .ZN(G282));
  NAND2_X1  g210(.A1(new_n465), .A2(new_n481), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  OAI221_X1 g214(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n488), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G135), .B2(new_n490), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT85), .B(G2096), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  INV_X1    g224(.A(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2427), .ZN(new_n652));
  INV_X1    g227(.A(G2430), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(KEYINPUT87), .ZN(new_n661));
  INV_X1    g236(.A(new_n659), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2451), .B(G2454), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n668));
  XOR2_X1   g243(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n660), .A2(new_n663), .A3(new_n669), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  INV_X1    g254(.A(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n680), .B2(new_n681), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n675), .A2(new_n677), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n676), .B1(new_n685), .B2(KEYINPUT17), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n679), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(KEYINPUT89), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G2096), .ZN(new_n691));
  INV_X1    g266(.A(G2096), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT90), .B(G2100), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(G1971), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1956), .B(G2474), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1961), .B(G1966), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT20), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(KEYINPUT92), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n700), .B2(new_n704), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n714), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  MUX2_X1   g294(.A(G6), .B(G305), .S(G16), .Z(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G23), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n582), .B2(new_n723), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT33), .B(G1976), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G166), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G22), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n722), .B(new_n731), .C1(new_n730), .C2(new_n729), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT34), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(KEYINPUT34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n600), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G16), .B2(G24), .ZN(new_n737));
  INV_X1    g312(.A(G1986), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(G25), .A2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n490), .A2(G131), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT93), .Z(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n744));
  INV_X1    g319(.A(G107), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n467), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n487), .B2(G119), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n741), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n750), .B(new_n752), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n735), .A2(new_n739), .A3(new_n740), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n734), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT36), .Z(new_n756));
  NAND2_X1  g331(.A1(G162), .A2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G29), .B2(G35), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT29), .ZN(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n490), .A2(G139), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n764), .B(new_n765), .C1(new_n468), .C2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G33), .B(new_n767), .S(G29), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2072), .Z(new_n769));
  NOR2_X1   g344(.A1(G171), .A2(new_n723), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G5), .B2(new_n723), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT24), .B(G34), .ZN(new_n774));
  INV_X1    g349(.A(G29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT98), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n483), .B2(new_n775), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n761), .A2(new_n769), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n759), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(G2090), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n624), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1348), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G11), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT30), .B(G28), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n644), .B2(new_n775), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT100), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n775), .A2(G32), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n487), .A2(G129), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n481), .A2(G105), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT26), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n796), .B(new_n798), .C1(new_n490), .C2(G141), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(new_n775), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT27), .B(G1996), .Z(new_n803));
  AOI211_X1 g378(.A(new_n786), .B(new_n791), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G19), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n562), .B2(G16), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1341), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n723), .A2(G21), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G168), .B2(new_n723), .ZN(new_n809));
  INV_X1    g384(.A(G1966), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n807), .B(new_n811), .C1(new_n779), .C2(new_n778), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n775), .A2(G26), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT28), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n487), .A2(G128), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n490), .A2(G140), .ZN(new_n816));
  NOR2_X1   g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT95), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT96), .B(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n802), .B2(new_n803), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n723), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT23), .ZN(new_n826));
  INV_X1    g401(.A(G299), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n723), .ZN(new_n828));
  INV_X1    g403(.A(G1956), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n772), .B2(new_n771), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n812), .A2(new_n824), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G27), .A2(G29), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G164), .B2(G29), .ZN(new_n834));
  INV_X1    g409(.A(G2078), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n783), .A2(new_n804), .A3(new_n832), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n756), .A2(new_n837), .ZN(G311));
  INV_X1    g413(.A(G311), .ZN(G150));
  AOI22_X1  g414(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n521), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n526), .A2(G55), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT101), .B(G93), .Z(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n559), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n562), .A2(new_n845), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n555), .A2(new_n561), .B1(new_n841), .B2(new_n844), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT38), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n624), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT102), .Z(new_n856));
  OAI21_X1  g431(.A(new_n846), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n848), .B1(new_n856), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(KEYINPUT105), .B(G37), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n487), .A2(G130), .ZN(new_n861));
  OAI221_X1 g436(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n490), .A2(G142), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n637), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n748), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n505), .A2(new_n507), .ZN(new_n867));
  INV_X1    g442(.A(new_n500), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n820), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n820), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n800), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n767), .A2(KEYINPUT104), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n800), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(new_n866), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n872), .A4(new_n873), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n767), .A2(KEYINPUT104), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n876), .B2(new_n879), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G162), .B(new_n483), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n643), .B(KEYINPUT103), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n860), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n881), .B2(new_n882), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NOR3_X1   g466(.A1(new_n841), .A2(new_n844), .A3(G868), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n624), .B2(G299), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n622), .A2(new_n623), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n612), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT83), .B1(new_n618), .B2(new_n612), .ZN(new_n898));
  OAI211_X1 g473(.A(G299), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(KEYINPUT106), .A3(new_n827), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n894), .A2(new_n895), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n827), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT41), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n631), .B(new_n851), .ZN(new_n907));
  MUX2_X1   g482(.A(new_n906), .B(new_n904), .S(new_n907), .Z(new_n908));
  XOR2_X1   g483(.A(G303), .B(G305), .Z(new_n909));
  INV_X1    g484(.A(new_n599), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n582), .B1(new_n910), .B2(new_n597), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n598), .A2(G288), .A3(new_n599), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G305), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n911), .B2(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT42), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n908), .B(new_n920), .Z(new_n921));
  INV_X1    g496(.A(new_n918), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n922), .B2(KEYINPUT108), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n921), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n892), .B1(new_n924), .B2(G868), .ZN(G295));
  AOI21_X1  g500(.A(new_n892), .B1(new_n924), .B2(G868), .ZN(G331));
  AND3_X1   g501(.A1(new_n549), .A2(KEYINPUT109), .A3(new_n551), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT109), .B1(new_n549), .B2(new_n551), .ZN(new_n928));
  OAI21_X1  g503(.A(G168), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(G301), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n549), .A2(KEYINPUT109), .A3(new_n551), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G286), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n933), .A3(new_n851), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n929), .A2(new_n933), .A3(new_n851), .A4(KEYINPUT110), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n933), .ZN(new_n938));
  INV_X1    g513(.A(new_n851), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n929), .A2(new_n933), .A3(new_n851), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n851), .B1(new_n929), .B2(new_n933), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n941), .A2(new_n906), .B1(new_n944), .B2(new_n904), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n918), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n902), .A2(new_n905), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n935), .B2(new_n934), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n937), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n944), .A2(new_n904), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n922), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT111), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT111), .B(new_n952), .C1(new_n945), .C2(new_n918), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n946), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  INV_X1    g533(.A(new_n946), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n941), .A2(new_n906), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n944), .A2(new_n904), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n918), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n963), .B2(G37), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n959), .B1(new_n964), .B2(new_n954), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n959), .A2(new_n860), .ZN(new_n968));
  AND4_X1   g543(.A1(KEYINPUT41), .A2(new_n894), .A3(new_n899), .A4(new_n901), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n944), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n895), .B1(new_n942), .B2(new_n943), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n941), .A2(new_n974), .B1(new_n903), .B2(new_n899), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n922), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n966), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n957), .A2(new_n967), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n968), .A2(new_n976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(KEYINPUT43), .B2(new_n956), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(KEYINPUT44), .B2(new_n982), .ZN(G397));
  NAND2_X1  g558(.A1(new_n572), .A2(new_n576), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT121), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n985), .A2(new_n577), .A3(new_n575), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(KEYINPUT121), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT57), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n827), .A2(KEYINPUT57), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT122), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G164), .B2(G1384), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  INV_X1    g569(.A(new_n507), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT4), .ZN(new_n996));
  INV_X1    g571(.A(G138), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n479), .A2(new_n997), .A3(new_n467), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(KEYINPUT71), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n999), .B2(new_n503), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT50), .B(new_n994), .C1(new_n1000), .C2(new_n500), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n475), .A2(G40), .A3(new_n482), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n829), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n867), .B2(new_n868), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(KEYINPUT115), .A3(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n475), .A2(G40), .A3(new_n482), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n994), .B1(new_n1000), .B2(new_n500), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n994), .C1(new_n1000), .C2(new_n500), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT56), .B(G2072), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1007), .A2(new_n1011), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n991), .B1(new_n1005), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2067), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n869), .A2(new_n994), .A3(new_n1019), .A4(new_n1003), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT123), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1006), .A2(KEYINPUT123), .A3(new_n1019), .A4(new_n1003), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1348), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1004), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n900), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1005), .A2(new_n991), .A3(new_n1017), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1018), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT61), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1005), .A2(new_n991), .A3(new_n1017), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(new_n1018), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1008), .B1(new_n993), .B2(new_n1001), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G1348), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(new_n1024), .A3(new_n624), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT60), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  OR4_X1    g612(.A1(KEYINPUT60), .A2(new_n1035), .A3(new_n1024), .A4(new_n900), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n991), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1017), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(G1956), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT61), .A3(new_n1029), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1007), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1009), .A2(new_n1008), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT58), .B(G1341), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1046), .A2(G1996), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1049), .B2(new_n562), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1049), .A2(new_n1045), .A3(new_n562), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1030), .B1(new_n1039), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1002), .A2(new_n1054), .A3(new_n779), .A4(new_n1003), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1003), .A3(new_n1012), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n810), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1034), .B2(new_n779), .ZN(new_n1060));
  OAI21_X1  g635(.A(G286), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT51), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1002), .A2(new_n779), .A3(new_n1003), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT120), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(G168), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(G8), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1065), .B2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1007), .A2(new_n1011), .A3(new_n835), .A4(new_n1014), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT124), .B(G1961), .Z(new_n1074));
  OR2_X1    g649(.A1(new_n1034), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n472), .A2(new_n467), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1072), .A2(G2078), .ZN(new_n1077));
  AND4_X1   g652(.A1(G40), .A2(new_n482), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1007), .A2(new_n1056), .A3(new_n1014), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1073), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1077), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1034), .A2(new_n1074), .B1(new_n1057), .B2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1081), .B(KEYINPUT54), .C1(new_n1085), .C2(G171), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n582), .A2(G1976), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT117), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  INV_X1    g664(.A(G8), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1047), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n869), .A2(new_n994), .A3(new_n1003), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n582), .B2(G1976), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1088), .B(new_n1097), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT118), .B(G1981), .Z(new_n1100));
  NAND4_X1  g675(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n587), .B1(new_n521), .B2(new_n584), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G1981), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1047), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT116), .B1(new_n1092), .B2(G8), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT119), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1107), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G166), .A2(new_n1090), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(KEYINPUT55), .Z(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1046), .A2(new_n730), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1004), .A2(G2090), .ZN(new_n1120));
  OAI211_X1 g695(.A(G8), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1046), .A2(new_n730), .B1(new_n1034), .B2(new_n760), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(new_n1090), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1099), .A2(new_n1115), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G171), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1073), .A2(new_n1075), .A3(G301), .A4(new_n1079), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT54), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1053), .A2(new_n1070), .A3(new_n1086), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1064), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1067), .B1(new_n1131), .B2(G286), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1065), .A2(G8), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1068), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1101), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G288), .A2(G1976), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1115), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1112), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1097), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1094), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1113), .B1(new_n1112), .B2(new_n1107), .ZN(new_n1145));
  AOI211_X1 g720(.A(KEYINPUT119), .B(new_n1106), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1146));
  OAI221_X1 g721(.A(new_n1144), .B1(new_n1095), .B2(new_n1094), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1141), .A2(new_n1142), .B1(new_n1147), .B2(new_n1121), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1149), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1131), .A2(G8), .A3(G168), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1150), .A2(new_n1151), .A3(KEYINPUT63), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1124), .B2(new_n1152), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1148), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1129), .A2(new_n1138), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1003), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n820), .B(new_n1019), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1160), .A2(KEYINPUT114), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT114), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1160), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1161), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n800), .B(G1996), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1162), .B(new_n1166), .C1(new_n1164), .C2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n748), .A2(new_n752), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n749), .A2(new_n751), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1164), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n600), .B(new_n738), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1158), .A2(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1160), .A2(G1996), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT46), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1164), .B1(new_n800), .B2(new_n1165), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1160), .A2(G1986), .A3(G290), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT48), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n820), .A2(G2067), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT125), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1160), .B1(new_n1185), .B2(KEYINPUT125), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1175), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1191));
  INV_X1    g765(.A(G319), .ZN(new_n1192));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(G227), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n1194), .B(G319), .C1(new_n695), .C2(new_n696), .ZN(new_n1195));
  NAND4_X1  g769(.A1(new_n673), .A2(new_n1193), .A3(new_n718), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n887), .B2(new_n889), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n978), .A2(new_n1191), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1191), .B1(new_n978), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  NAND2_X1  g774(.A1(new_n978), .A2(new_n1197), .ZN(G225));
endmodule


