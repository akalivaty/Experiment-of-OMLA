

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U324 ( .A(n406), .B(n405), .ZN(n439) );
  XNOR2_X1 U325 ( .A(n408), .B(n407), .ZN(n409) );
  NOR2_X1 U326 ( .A1(n395), .A2(n394), .ZN(n498) );
  XNOR2_X1 U327 ( .A(KEYINPUT28), .B(n480), .ZN(n548) );
  XOR2_X1 U328 ( .A(n445), .B(n444), .Z(n292) );
  XOR2_X1 U329 ( .A(n469), .B(n468), .Z(n293) );
  INV_X1 U330 ( .A(KEYINPUT54), .ZN(n475) );
  AND2_X1 U331 ( .A1(n388), .A2(n530), .ZN(n382) );
  INV_X1 U332 ( .A(KEYINPUT92), .ZN(n355) );
  XNOR2_X1 U333 ( .A(n382), .B(KEYINPUT95), .ZN(n543) );
  XNOR2_X1 U334 ( .A(n439), .B(n409), .ZN(n410) );
  XNOR2_X1 U335 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U336 ( .A(n358), .B(n357), .ZN(n359) );
  NOR2_X1 U337 ( .A1(n486), .A2(n559), .ZN(n583) );
  NAND2_X1 U338 ( .A1(n460), .A2(n459), .ZN(n563) );
  NOR2_X1 U339 ( .A1(n545), .A2(n482), .ZN(n577) );
  INV_X1 U340 ( .A(G43GAT), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n451), .B(KEYINPUT38), .ZN(n514) );
  XNOR2_X1 U342 ( .A(n483), .B(G176GAT), .ZN(n484) );
  XNOR2_X1 U343 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n485), .B(n484), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(G169GAT), .B(G113GAT), .Z(n424) );
  XNOR2_X1 U347 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n294), .B(KEYINPUT18), .ZN(n360) );
  XOR2_X1 U349 ( .A(n424), .B(n360), .Z(n296) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(n297), .B(G71GAT), .Z(n301) );
  XOR2_X1 U353 ( .A(G120GAT), .B(G127GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n371) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(n371), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n309) );
  XOR2_X1 U358 ( .A(G134GAT), .B(G190GAT), .Z(n303) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G99GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U361 ( .A(G176GAT), .B(G183GAT), .Z(n305) );
  XNOR2_X1 U362 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U364 ( .A(n307), .B(n306), .Z(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n545) );
  INV_X1 U366 ( .A(n545), .ZN(n534) );
  XOR2_X1 U367 ( .A(G64GAT), .B(G211GAT), .Z(n311) );
  XNOR2_X1 U368 ( .A(G127GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U370 ( .A(KEYINPUT14), .B(KEYINPUT84), .Z(n313) );
  XNOR2_X1 U371 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n325) );
  XOR2_X1 U374 ( .A(G8GAT), .B(G183GAT), .Z(n347) );
  XNOR2_X1 U375 ( .A(G15GAT), .B(G1GAT), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n316), .B(KEYINPUT69), .ZN(n425) );
  XOR2_X1 U377 ( .A(n425), .B(KEYINPUT83), .Z(n318) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U380 ( .A(n347), .B(n319), .Z(n323) );
  XOR2_X1 U381 ( .A(G22GAT), .B(G155GAT), .Z(n337) );
  XOR2_X1 U382 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n321) );
  XNOR2_X1 U383 ( .A(G71GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n447) );
  XNOR2_X1 U385 ( .A(n337), .B(n447), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n593) );
  INV_X1 U388 ( .A(n593), .ZN(n495) );
  XOR2_X1 U389 ( .A(KEYINPUT74), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U390 ( .A(G148GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U392 ( .A(KEYINPUT73), .B(n328), .Z(n450) );
  XOR2_X1 U393 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n330) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U396 ( .A(n331), .B(KEYINPUT24), .Z(n336) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n332), .B(KEYINPUT3), .ZN(n379) );
  XOR2_X1 U399 ( .A(G211GAT), .B(KEYINPUT21), .Z(n334) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n334), .B(n333), .ZN(n354) );
  XNOR2_X1 U402 ( .A(n379), .B(n354), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U404 ( .A(KEYINPUT87), .B(KEYINPUT89), .Z(n339) );
  XOR2_X1 U405 ( .A(G218GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U406 ( .A(n415), .B(n337), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U408 ( .A(n341), .B(n340), .Z(n343) );
  XNOR2_X1 U409 ( .A(G50GAT), .B(G106GAT), .ZN(n342) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n450), .B(n344), .ZN(n480) );
  XOR2_X1 U412 ( .A(KEYINPUT93), .B(G92GAT), .Z(n346) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U415 ( .A(G190GAT), .B(KEYINPUT81), .Z(n401) );
  XOR2_X1 U416 ( .A(n347), .B(n401), .Z(n349) );
  XNOR2_X1 U417 ( .A(G36GAT), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U419 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n353), .B(n352), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n354), .B(KEYINPUT94), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G64GAT), .ZN(n361) );
  XOR2_X1 U425 ( .A(n361), .B(KEYINPUT75), .Z(n446) );
  XNOR2_X1 U426 ( .A(n362), .B(n446), .ZN(n503) );
  XOR2_X1 U427 ( .A(KEYINPUT27), .B(n503), .Z(n388) );
  XOR2_X1 U428 ( .A(G85GAT), .B(G162GAT), .Z(n364) );
  XNOR2_X1 U429 ( .A(G29GAT), .B(G148GAT), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U431 ( .A(G57GAT), .B(G155GAT), .Z(n366) );
  XNOR2_X1 U432 ( .A(G113GAT), .B(G1GAT), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U434 ( .A(n368), .B(n367), .Z(n377) );
  XOR2_X1 U435 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n370) );
  XNOR2_X1 U436 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U438 ( .A(G134GAT), .B(KEYINPUT80), .Z(n402) );
  XOR2_X1 U439 ( .A(n402), .B(n371), .Z(n373) );
  NAND2_X1 U440 ( .A1(G225GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U444 ( .A(n378), .B(KEYINPUT4), .Z(n381) );
  XNOR2_X1 U445 ( .A(n379), .B(KEYINPUT5), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n530) );
  NOR2_X1 U447 ( .A1(n548), .A2(n543), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n383), .A2(n545), .ZN(n384) );
  XOR2_X1 U449 ( .A(KEYINPUT96), .B(n384), .Z(n395) );
  NOR2_X1 U450 ( .A1(n545), .A2(n503), .ZN(n385) );
  NOR2_X1 U451 ( .A1(n480), .A2(n385), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n386), .B(KEYINPUT25), .ZN(n391) );
  NAND2_X1 U453 ( .A1(n480), .A2(n545), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n387), .B(KEYINPUT26), .ZN(n559) );
  INV_X1 U455 ( .A(n559), .ZN(n389) );
  NAND2_X1 U456 ( .A1(n389), .A2(n388), .ZN(n390) );
  NAND2_X1 U457 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U458 ( .A(KEYINPUT97), .B(n392), .ZN(n393) );
  NOR2_X1 U459 ( .A1(n530), .A2(n393), .ZN(n394) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n419) );
  XOR2_X1 U461 ( .A(G43GAT), .B(G29GAT), .Z(n397) );
  XNOR2_X1 U462 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U464 ( .A(n398), .B(KEYINPUT68), .Z(n400) );
  XNOR2_X1 U465 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n400), .B(n399), .ZN(n438) );
  XOR2_X1 U467 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n404) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n411) );
  XOR2_X1 U470 ( .A(G92GAT), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U471 ( .A(G99GAT), .B(G106GAT), .ZN(n405) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n408) );
  INV_X1 U473 ( .A(KEYINPUT10), .ZN(n407) );
  XOR2_X1 U474 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U475 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n413) );
  XNOR2_X1 U476 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U480 ( .A(n438), .B(n418), .Z(n466) );
  XOR2_X1 U481 ( .A(KEYINPUT82), .B(n466), .Z(n578) );
  XOR2_X1 U482 ( .A(n419), .B(n578), .Z(n487) );
  NOR2_X1 U483 ( .A1(n498), .A2(n487), .ZN(n420) );
  NAND2_X1 U484 ( .A1(n495), .A2(n420), .ZN(n423) );
  XNOR2_X1 U485 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n421), .B(KEYINPUT37), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n529) );
  XOR2_X1 U488 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(G141GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U491 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n429) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n436) );
  XOR2_X1 U495 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n433) );
  XNOR2_X1 U496 ( .A(G197GAT), .B(G8GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n434), .B(KEYINPUT66), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n584) );
  INV_X1 U501 ( .A(n584), .ZN(n516) );
  XNOR2_X1 U502 ( .A(n516), .B(KEYINPUT71), .ZN(n573) );
  XOR2_X1 U503 ( .A(KEYINPUT76), .B(n439), .Z(n441) );
  NAND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U506 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n443) );
  XNOR2_X1 U507 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n442) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U509 ( .A(n447), .B(n446), .Z(n448) );
  XNOR2_X1 U510 ( .A(n292), .B(n448), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n456) );
  BUF_X1 U512 ( .A(n456), .Z(n588) );
  NAND2_X1 U513 ( .A1(n573), .A2(n588), .ZN(n500) );
  NOR2_X1 U514 ( .A1(n529), .A2(n500), .ZN(n451) );
  NAND2_X1 U515 ( .A1(n534), .A2(n514), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n453) );
  NAND2_X1 U517 ( .A1(KEYINPUT41), .A2(n456), .ZN(n460) );
  INV_X1 U518 ( .A(KEYINPUT41), .ZN(n458) );
  INV_X1 U519 ( .A(n456), .ZN(n457) );
  NAND2_X1 U520 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U521 ( .A(n563), .B(KEYINPUT107), .Z(n551) );
  INV_X1 U522 ( .A(KEYINPUT64), .ZN(n479) );
  NOR2_X1 U523 ( .A1(n487), .A2(n495), .ZN(n462) );
  INV_X1 U524 ( .A(KEYINPUT45), .ZN(n461) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(n465) );
  INV_X1 U526 ( .A(n573), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n588), .A2(n463), .ZN(n464) );
  NOR2_X1 U528 ( .A1(n465), .A2(n464), .ZN(n473) );
  BUF_X1 U529 ( .A(n466), .Z(n571) );
  XNOR2_X1 U530 ( .A(n593), .B(KEYINPUT114), .ZN(n575) );
  XOR2_X1 U531 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n467) );
  XNOR2_X1 U532 ( .A(KEYINPUT115), .B(n467), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n584), .A2(n563), .ZN(n468) );
  NOR2_X1 U534 ( .A1(n575), .A2(n293), .ZN(n470) );
  NAND2_X1 U535 ( .A1(n571), .A2(n470), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n471), .B(KEYINPUT47), .ZN(n472) );
  NOR2_X1 U537 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n474), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U539 ( .A1(n542), .A2(n503), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U541 ( .A1(n530), .A2(n477), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(n486) );
  NOR2_X1 U543 ( .A1(n486), .A2(n480), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NAND2_X1 U545 ( .A1(n551), .A2(n577), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n483) );
  INV_X1 U547 ( .A(n583), .ZN(n589) );
  NOR2_X1 U548 ( .A1(n487), .A2(n589), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT126), .B(n490), .ZN(n492) );
  XOR2_X1 U552 ( .A(G218GAT), .B(KEYINPUT125), .Z(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1355GAT) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT34), .ZN(n494) );
  XOR2_X1 U556 ( .A(KEYINPUT100), .B(n494), .Z(n502) );
  NOR2_X1 U557 ( .A1(n578), .A2(n495), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT16), .B(n496), .Z(n497) );
  NOR2_X1 U559 ( .A1(n498), .A2(n497), .ZN(n499) );
  XOR2_X1 U560 ( .A(KEYINPUT98), .B(n499), .Z(n518) );
  NOR2_X1 U561 ( .A1(n518), .A2(n500), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n530), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1324GAT) );
  XOR2_X1 U564 ( .A(G8GAT), .B(KEYINPUT101), .Z(n505) );
  INV_X1 U565 ( .A(n503), .ZN(n532) );
  NAND2_X1 U566 ( .A1(n508), .A2(n532), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1325GAT) );
  XOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U569 ( .A1(n508), .A2(n534), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n548), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U573 ( .A(G29GAT), .B(KEYINPUT39), .Z(n511) );
  NAND2_X1 U574 ( .A1(n530), .A2(n514), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  XOR2_X1 U576 ( .A(G36GAT), .B(KEYINPUT105), .Z(n513) );
  NAND2_X1 U577 ( .A1(n532), .A2(n514), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1329GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n548), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n520) );
  NAND2_X1 U582 ( .A1(n551), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT108), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n518), .A2(n528), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n525), .A2(n530), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n532), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U590 ( .A1(n525), .A2(n534), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT110), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G71GAT), .B(n524), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U594 ( .A1(n525), .A2(n548), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n530), .A2(n537), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G85GAT), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U601 ( .A(G99GAT), .B(KEYINPUT111), .Z(n536) );
  NAND2_X1 U602 ( .A1(n537), .A2(n534), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1338GAT) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n541) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U606 ( .A1(n537), .A2(n548), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(KEYINPUT117), .ZN(n560) );
  NOR2_X1 U611 ( .A1(n545), .A2(n560), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n546), .Z(n547) );
  NOR2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n573), .A2(n556), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT119), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G113GAT), .B(n550), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(G120GAT), .B(KEYINPUT49), .Z(n553) );
  NAND2_X1 U618 ( .A1(n556), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1341GAT) );
  NAND2_X1 U620 ( .A1(n575), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT50), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G127GAT), .B(n555), .ZN(G1342GAT) );
  XOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U624 ( .A1(n556), .A2(n578), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT120), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n584), .A2(n569), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G141GAT), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n569), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G148GAT), .B(n566), .ZN(G1345GAT) );
  XOR2_X1 U634 ( .A(G155GAT), .B(KEYINPUT121), .Z(n568) );
  NAND2_X1 U635 ( .A1(n593), .A2(n569), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(G1346GAT) );
  INV_X1 U637 ( .A(n569), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(G162GAT), .B(n572), .Z(G1347GAT) );
  NAND2_X1 U640 ( .A1(n577), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(G169GAT), .B(n574), .ZN(G1348GAT) );
  NAND2_X1 U642 ( .A1(n575), .A2(n577), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n582) );
  XNOR2_X1 U645 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT122), .ZN(n580) );
  XNOR2_X1 U647 ( .A(KEYINPUT58), .B(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1351GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n586) );
  NAND2_X1 U650 ( .A1(n583), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(n587), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n591) );
  OR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G204GAT), .B(n592), .ZN(G1353GAT) );
  NAND2_X1 U657 ( .A1(n583), .A2(n593), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
endmodule

