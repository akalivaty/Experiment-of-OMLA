//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1305, new_n1306, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n206), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n211), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT14), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G226), .A2(G1698), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(new_n232), .B2(G1698), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n225), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT13), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT65), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n258), .B2(new_n225), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n257), .A2(KEYINPUT65), .A3(G1), .A4(G13), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n263), .A2(G274), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n266), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n263), .A2(new_n269), .A3(G238), .A4(new_n267), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n260), .A2(new_n261), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n252), .A2(new_n253), .B1(G33), .B2(G97), .ZN(new_n272));
  INV_X1    g0072(.A(new_n259), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n268), .B(new_n270), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n250), .B1(new_n276), .B2(G169), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(new_n275), .A3(G179), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(G169), .A3(new_n250), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT71), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n225), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT66), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G68), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n286), .A2(G50), .B1(G20), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n206), .A2(G33), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n213), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT11), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(new_n225), .A3(new_n283), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n205), .A2(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G68), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT68), .B1(new_n296), .B2(new_n300), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT12), .B1(new_n295), .B2(G68), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n295), .A2(KEYINPUT12), .A3(G68), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT69), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n293), .B(new_n294), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n303), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n304), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n282), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n293), .A2(new_n294), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n306), .A2(new_n307), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n314), .A2(KEYINPUT71), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n281), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n276), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n314), .A2(new_n316), .A3(new_n315), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n271), .B2(new_n275), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n273), .B1(new_n213), .B2(new_n333), .ZN(new_n334));
  MUX2_X1   g0134(.A(G222), .B(G223), .S(G1698), .Z(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n263), .A2(new_n267), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n269), .ZN(new_n338));
  INV_X1    g0138(.A(G226), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n268), .B(new_n336), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n286), .A2(G150), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT8), .B(G58), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n289), .ZN(new_n345));
  INV_X1    g0145(.A(G50), .ZN(new_n346));
  INV_X1    g0146(.A(new_n295), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(new_n285), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT66), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n284), .B(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n350), .A2(G50), .A3(new_n295), .A4(new_n299), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n341), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(KEYINPUT9), .A3(new_n351), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n340), .A2(new_n322), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT10), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n355), .A2(new_n360), .A3(new_n356), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n340), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g0164(.A(KEYINPUT67), .B(G179), .Z(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(new_n352), .C1(new_n366), .C2(new_n340), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n299), .A2(G77), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n296), .A2(new_n368), .B1(G77), .B2(new_n295), .ZN(new_n369));
  INV_X1    g0169(.A(new_n344), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n289), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(new_n284), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G1698), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n253), .A2(G232), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n375), .B(new_n377), .C1(new_n215), .C2(new_n253), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n259), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n268), .C1(new_n214), .C2(new_n338), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n374), .B1(new_n380), .B2(new_n363), .ZN(new_n381));
  INV_X1    g0181(.A(new_n338), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G244), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n383), .A2(new_n268), .A3(new_n365), .A4(new_n379), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(G200), .ZN(new_n387));
  INV_X1    g0187(.A(new_n374), .ZN(new_n388));
  INV_X1    g0188(.A(new_n380), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(G190), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n328), .A2(new_n362), .A3(new_n367), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n350), .A2(new_n295), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n370), .A2(new_n299), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n295), .B2(new_n370), .ZN(new_n395));
  INV_X1    g0195(.A(new_n284), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n253), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n333), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G68), .ZN(new_n401));
  INV_X1    g0201(.A(G58), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n287), .ZN(new_n403));
  OAI21_X1  g0203(.A(G20), .B1(new_n403), .B2(new_n201), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n286), .A2(G159), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n396), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT72), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n329), .A3(KEYINPUT3), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT7), .A2(G20), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n411), .A2(new_n206), .A3(new_n413), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n287), .B1(new_n420), .B2(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n395), .B1(new_n410), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n376), .A2(G223), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT75), .B1(new_n414), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT75), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n429), .B(new_n426), .C1(new_n411), .C2(new_n413), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n376), .B1(new_n411), .B2(new_n413), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n273), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n263), .A2(new_n269), .A3(G232), .A4(new_n267), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n268), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n425), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n331), .A2(KEYINPUT72), .A3(G33), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n253), .B2(KEYINPUT72), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n429), .B1(new_n439), .B2(new_n426), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G87), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n414), .A2(G226), .A3(G1698), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n414), .A2(KEYINPUT75), .A3(new_n427), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n259), .ZN(new_n445));
  INV_X1    g0245(.A(new_n436), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(KEYINPUT76), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(G200), .B1(new_n437), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n434), .A2(G190), .A3(new_n436), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n424), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT76), .B1(new_n445), .B2(new_n446), .ZN(new_n453));
  AOI211_X1 g0253(.A(new_n425), .B(new_n436), .C1(new_n444), .C2(new_n259), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n363), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n395), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n409), .B(new_n406), .C1(new_n419), .C2(new_n421), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n406), .B1(new_n400), .B2(G68), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n284), .B1(new_n458), .B2(KEYINPUT16), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n456), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT74), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(KEYINPUT74), .B(new_n456), .C1(new_n457), .C2(new_n459), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n434), .A2(new_n436), .A3(new_n366), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n455), .A2(new_n462), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT18), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n437), .A2(new_n447), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n464), .B1(new_n468), .B2(new_n363), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n462), .A4(new_n463), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n325), .B1(new_n453), .B2(new_n454), .ZN(new_n472));
  INV_X1    g0272(.A(new_n449), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT17), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n452), .A2(new_n467), .A3(new_n471), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n205), .A2(G45), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(G257), .A3(new_n263), .A4(new_n267), .ZN(new_n483));
  INV_X1    g0283(.A(new_n481), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n477), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(G274), .A3(new_n263), .A4(new_n267), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n488));
  AND2_X1   g0288(.A1(KEYINPUT4), .A2(G244), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n330), .A2(new_n332), .A3(new_n489), .A4(new_n376), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n414), .A2(G244), .A3(new_n376), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n487), .B1(new_n495), .B2(new_n273), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT77), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT77), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n487), .C1(new_n495), .C2(new_n273), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n350), .B(new_n295), .C1(G1), .C2(new_n329), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  OR2_X1    g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  XOR2_X1   g0304(.A(G97), .B(G107), .Z(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n400), .A2(G107), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n284), .B1(new_n502), .B2(new_n347), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n500), .A2(new_n363), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n365), .B(new_n487), .C1(new_n495), .C2(new_n273), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT78), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n497), .A2(G190), .A3(new_n499), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n496), .A2(G200), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n503), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n511), .A2(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n216), .A2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G257), .B2(G1698), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n413), .B2(new_n411), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n253), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n259), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n482), .A2(G270), .A3(new_n263), .A4(new_n267), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(G190), .A3(new_n486), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n205), .B2(G33), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n297), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(KEYINPUT79), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT79), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n532), .A3(G20), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G13), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(G1), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n491), .B(new_n206), .C1(G33), .C2(new_n502), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n284), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n533), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n539), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n526), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n525), .A2(new_n486), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n325), .B1(new_n546), .B2(new_n524), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT82), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n524), .A2(new_n486), .A3(new_n525), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n544), .A4(new_n526), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n542), .A2(new_n543), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n297), .A2(new_n528), .B1(new_n534), .B2(new_n536), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n363), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(KEYINPUT21), .A3(new_n549), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n555), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(G179), .A3(new_n524), .A4(new_n546), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT21), .B1(new_n556), .B2(new_n549), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n214), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G238), .B2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n413), .B2(new_n411), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n329), .B1(new_n530), .B2(new_n532), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n259), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n478), .A2(G250), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n477), .A2(G274), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n263), .A3(new_n267), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(KEYINPUT80), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT80), .B1(new_n568), .B2(new_n571), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n372), .A2(new_n347), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n414), .A2(new_n206), .A3(G68), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  INV_X1    g0378(.A(G87), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n578), .A2(new_n579), .B1(new_n255), .B2(new_n206), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G97), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n580), .A2(new_n581), .B1(new_n289), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n576), .B1(new_n584), .B2(new_n396), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n501), .A2(new_n579), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n568), .A2(new_n571), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G190), .A3(new_n572), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n575), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n363), .B1(new_n573), .B2(new_n574), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n365), .A3(new_n572), .ZN(new_n594));
  XOR2_X1   g0394(.A(new_n372), .B(KEYINPUT81), .Z(new_n595));
  OAI221_X1 g0395(.A(new_n576), .B1(new_n501), .B2(new_n595), .C1(new_n584), .C2(new_n396), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n563), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(KEYINPUT22), .A2(G87), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n439), .A2(G20), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n567), .A2(new_n206), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n206), .A2(G87), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n333), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT23), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n206), .B2(G107), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n215), .A2(KEYINPUT23), .A3(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n602), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT24), .B1(new_n601), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n414), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n567), .A2(new_n206), .B1(new_n607), .B2(new_n608), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n605), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n284), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n347), .A2(new_n215), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT25), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n501), .B2(new_n215), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT83), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n396), .B1(new_n611), .B2(new_n615), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n624), .A2(new_n625), .A3(new_n621), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n486), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n414), .A2(G250), .A3(new_n376), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n414), .A2(G257), .A3(G1698), .ZN(new_n630));
  NAND2_X1  g0430(.A1(G33), .A2(G294), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n628), .B1(new_n632), .B2(new_n259), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n482), .A2(G264), .A3(new_n263), .A4(new_n267), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G169), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n259), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n337), .A2(new_n638), .A3(G264), .A4(new_n482), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(KEYINPUT84), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n637), .A2(new_n641), .A3(G179), .A4(new_n486), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT85), .B1(new_n636), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n634), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n644), .B(new_n628), .C1(new_n632), .C2(new_n259), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n642), .B(KEYINPUT85), .C1(new_n645), .C2(new_n363), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n627), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n635), .A2(G190), .ZN(new_n649));
  AOI21_X1  g0449(.A(G200), .B1(new_n633), .B2(new_n641), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n617), .B(new_n622), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n518), .A2(new_n599), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n392), .A2(new_n476), .A3(new_n652), .ZN(G372));
  XNOR2_X1  g0453(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n469), .A2(new_n460), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n455), .A2(new_n460), .A3(new_n465), .ZN(new_n656));
  INV_X1    g0456(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n474), .A2(KEYINPUT17), .ZN(new_n660));
  AOI211_X1 g0460(.A(new_n451), .B(new_n460), .C1(new_n472), .C2(new_n473), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n321), .B1(new_n664), .B2(new_n386), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n659), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n362), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n367), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n392), .A2(new_n476), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n511), .A2(new_n513), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n517), .A2(new_n514), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n562), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n636), .A2(new_n642), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n617), .A2(new_n622), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n588), .A2(G200), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n587), .A2(new_n591), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n588), .A2(new_n363), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n594), .A2(new_n596), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n651), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n672), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT26), .B1(new_n670), .B2(new_n598), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n500), .A2(new_n363), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n686), .A2(new_n513), .A3(new_n516), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n682), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n689), .A3(new_n680), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n669), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n668), .A2(new_n691), .ZN(G369));
  AND2_X1   g0492(.A1(new_n648), .A2(new_n651), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n536), .A2(new_n206), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n536), .A2(new_n696), .A3(new_n206), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(G213), .A3(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT87), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n627), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n693), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT88), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT88), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n693), .A2(new_n707), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n703), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n648), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n544), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n673), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n563), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n562), .A2(new_n703), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n706), .A2(new_n708), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n674), .A2(new_n675), .A3(new_n710), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT89), .Z(G399));
  INV_X1    g0524(.A(new_n209), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n578), .A2(new_n579), .A3(new_n527), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(G1), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT91), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(new_n223), .B2(new_n727), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n731), .B2(new_n730), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT28), .Z(new_n734));
  NAND4_X1  g0534(.A1(new_n693), .A2(new_n518), .A3(new_n599), .A4(new_n710), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n549), .A2(new_n365), .A3(new_n588), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n633), .A2(new_n641), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n736), .A2(new_n737), .A3(new_n496), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT92), .ZN(new_n739));
  AND4_X1   g0539(.A1(G179), .A2(new_n524), .A3(new_n486), .A4(new_n525), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n632), .A2(new_n259), .B1(new_n639), .B2(new_n640), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n590), .A4(new_n572), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n739), .B1(new_n500), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n739), .B(new_n745), .C1(new_n500), .C2(new_n742), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n703), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n710), .B1(new_n744), .B2(new_n746), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT31), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n735), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n672), .A2(new_n683), .ZN(new_n756));
  INV_X1    g0556(.A(new_n648), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(KEYINPUT94), .C1(new_n757), .C2(new_n673), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT94), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(new_n673), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n518), .A2(new_n651), .A3(new_n682), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n687), .A2(new_n688), .A3(new_n597), .A4(new_n592), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT26), .B1(new_n670), .B2(new_n681), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n763), .A2(new_n680), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n758), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n710), .B1(new_n690), .B2(new_n684), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n755), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n734), .B1(new_n771), .B2(G1), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT95), .ZN(G364));
  NOR2_X1   g0573(.A1(new_n535), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n205), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n726), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n716), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G330), .B2(new_n714), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n209), .A2(new_n253), .ZN(new_n780));
  INV_X1    g0580(.A(G355), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n209), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n224), .A2(G45), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G45), .B2(new_n246), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n415), .A2(new_n417), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n725), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n782), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n225), .B1(G20), .B2(new_n363), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n777), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n206), .A2(G190), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G179), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT32), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n365), .A2(new_n206), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(new_n322), .A3(G200), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n800), .A2(new_n801), .B1(new_n287), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n801), .B2(new_n800), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n365), .A2(new_n796), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G77), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n206), .A2(G179), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n322), .A3(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n215), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(G190), .A3(G200), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n253), .B1(new_n815), .B2(new_n579), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n206), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n814), .B(new_n816), .C1(G97), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n802), .A2(G190), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n325), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(G200), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G50), .A2(new_n822), .B1(new_n823), .B2(G58), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n805), .A2(new_n811), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n815), .A2(new_n522), .ZN(new_n826));
  INV_X1    g0626(.A(new_n806), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n827), .A2(new_n828), .B1(new_n818), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n826), .B(new_n830), .C1(G329), .C2(new_n797), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n333), .B1(new_n813), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n803), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT98), .B(KEYINPUT33), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(G317), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G322), .ZN(new_n839));
  INV_X1    g0639(.A(new_n823), .ZN(new_n840));
  INV_X1    g0640(.A(new_n822), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT97), .B(G326), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n839), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n825), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n794), .B1(new_n844), .B2(new_n791), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n714), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n779), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  INV_X1    g0649(.A(KEYINPUT103), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT101), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n385), .B(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n390), .A2(new_n387), .B1(new_n388), .B2(new_n703), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n381), .A2(new_n384), .A3(new_n703), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n768), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n857), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n710), .B(new_n859), .C1(new_n690), .C2(new_n684), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n850), .B1(new_n861), .B2(new_n754), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n755), .A2(KEYINPUT103), .A3(new_n858), .A4(new_n860), .ZN(new_n863));
  INV_X1    g0663(.A(new_n777), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n754), .B2(new_n861), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n791), .A2(new_n788), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n777), .B1(G77), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT99), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n822), .A2(G137), .B1(new_n834), .B2(G150), .ZN(new_n875));
  INV_X1    g0675(.A(G143), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n876), .B2(new_n840), .C1(new_n799), .C2(new_n809), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT34), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G132), .A2(new_n797), .B1(new_n819), .B2(G58), .ZN(new_n879));
  INV_X1    g0679(.A(new_n815), .ZN(new_n880));
  INV_X1    g0680(.A(new_n813), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n880), .A2(G50), .B1(new_n881), .B2(G68), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n878), .A2(new_n785), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n834), .A2(KEYINPUT100), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n834), .A2(KEYINPUT100), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(G283), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n530), .A2(new_n532), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n810), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(G294), .A2(new_n823), .B1(new_n822), .B2(G303), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n333), .B1(new_n818), .B2(new_n502), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n798), .A2(new_n828), .B1(new_n813), .B2(new_n579), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n892), .B(new_n893), .C1(G107), .C2(new_n880), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n888), .A2(new_n890), .A3(new_n891), .A4(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n883), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n791), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n874), .B1(new_n789), .B2(new_n859), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n870), .A2(new_n898), .ZN(G384));
  NOR2_X1   g0699(.A1(new_n774), .A2(new_n205), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n423), .A2(new_n285), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n422), .B2(new_n407), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n456), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n701), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n476), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n455), .A2(new_n903), .A3(new_n465), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n450), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n701), .B(KEYINPUT106), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n462), .A2(new_n463), .A3(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n466), .A2(new_n450), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n907), .B2(new_n915), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT108), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT107), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n656), .B(new_n913), .C1(new_n474), .C2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n450), .A2(KEYINPUT107), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n654), .B1(new_n469), .B2(new_n460), .ZN(new_n925));
  AND4_X1   g0725(.A1(new_n460), .A2(new_n455), .A3(new_n465), .A4(new_n654), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n452), .B(new_n475), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n913), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n924), .A2(new_n914), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n929), .B2(KEYINPUT38), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  AND4_X1   g0732(.A1(new_n911), .A2(new_n466), .A3(new_n450), .A4(new_n913), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n450), .A2(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n472), .A2(new_n473), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n921), .A3(new_n424), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n934), .A2(new_n656), .A3(new_n936), .A4(new_n913), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n933), .B1(new_n937), .B2(KEYINPUT37), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n913), .B1(new_n662), .B2(new_n659), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT108), .B(new_n932), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n930), .A2(new_n931), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n919), .B1(new_n941), .B2(new_n918), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n320), .A2(new_n703), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n852), .A2(new_n703), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n860), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n313), .A2(new_n317), .A3(new_n703), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n280), .A2(new_n279), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n277), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n664), .B(new_n948), .C1(new_n950), .C2(new_n318), .ZN(new_n951));
  INV_X1    g0751(.A(new_n948), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT105), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n281), .C2(new_n327), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n952), .B1(new_n281), .B2(new_n327), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n947), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n916), .A2(new_n917), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(new_n659), .B2(new_n912), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n944), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n767), .A2(new_n669), .A3(new_n770), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n668), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n963), .B(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(G330), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n907), .A2(new_n915), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n932), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n931), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n857), .B1(new_n955), .B2(new_n957), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n652), .A2(new_n703), .B1(new_n751), .B2(KEYINPUT31), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n748), .A2(new_n749), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT109), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n753), .A2(new_n976), .A3(new_n971), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n970), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT40), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n974), .A2(new_n979), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n940), .A2(new_n931), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n927), .A2(new_n928), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n921), .B1(new_n935), .B2(new_n424), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n656), .A2(new_n913), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n911), .B1(new_n986), .B2(new_n936), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n983), .B1(new_n987), .B2(new_n933), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT108), .B1(new_n988), .B2(new_n932), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n981), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n753), .A2(new_n669), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n967), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n900), .B1(new_n966), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n966), .B2(new_n994), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n527), .B(new_n227), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(KEYINPUT35), .B2(new_n506), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT36), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n223), .A2(new_n213), .A3(new_n403), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n287), .A2(G50), .ZN(new_n1001));
  OAI211_X1 g0801(.A(G1), .B(new_n535), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n999), .A3(new_n1002), .ZN(G367));
  NAND2_X1  g0803(.A1(new_n516), .A2(new_n703), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n518), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n687), .A2(new_n703), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n720), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT42), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n757), .A2(new_n671), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n703), .B1(new_n1011), .B2(new_n670), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1009), .B2(KEYINPUT42), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n710), .A2(new_n587), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n682), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n680), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT43), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1014), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1010), .A2(new_n1013), .A3(new_n1021), .A4(new_n1020), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n717), .A2(new_n1008), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n726), .B(KEYINPUT41), .Z(new_n1029));
  NAND3_X1  g0829(.A1(new_n720), .A2(new_n721), .A3(new_n1007), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT110), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT110), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n720), .A2(new_n1032), .A3(new_n721), .A4(new_n1007), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT45), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n722), .A2(KEYINPUT44), .A3(new_n1008), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT44), .B1(new_n722), .B2(new_n1008), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1031), .A2(KEYINPUT45), .A3(new_n1033), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1038), .A3(new_n717), .A4(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n720), .A2(KEYINPUT111), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n711), .A2(new_n719), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n720), .A2(KEYINPUT111), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n716), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n715), .B(new_n1041), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1045), .A2(new_n771), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1034), .A2(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1039), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n718), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1040), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1029), .B1(new_n1051), .B2(new_n771), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1028), .B1(new_n1052), .B2(new_n776), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n792), .B1(new_n209), .B2(new_n372), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n786), .B2(new_n238), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(new_n864), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n887), .A2(G159), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n810), .A2(G50), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G143), .A2(new_n822), .B1(new_n823), .B2(G150), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n253), .B1(new_n813), .B2(new_n213), .ZN(new_n1060));
  INV_X1    g0860(.A(G137), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n798), .A2(new_n1061), .B1(new_n815), .B2(new_n402), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(G68), .C2(new_n819), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n785), .B1(new_n822), .B2(G311), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n840), .B2(new_n522), .C1(new_n832), .C2(new_n809), .ZN(new_n1066));
  INV_X1    g0866(.A(G317), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n798), .A2(new_n1067), .B1(new_n813), .B2(new_n502), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n880), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n215), .B2(new_n818), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT46), .B1(new_n880), .B2(new_n889), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n886), .B2(new_n829), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1064), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT47), .Z(new_n1075));
  OAI221_X1 g0875(.A(new_n1056), .B1(new_n846), .B2(new_n1019), .C1(new_n1075), .C2(new_n897), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1053), .A2(new_n1076), .ZN(G387));
  OAI21_X1  g0877(.A(new_n786), .B1(new_n235), .B2(new_n265), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n729), .B2(new_n780), .ZN(new_n1079));
  OR3_X1    g0879(.A1(new_n344), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT50), .B1(new_n344), .B2(G50), .ZN(new_n1081));
  AOI21_X1  g0881(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n729), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1079), .A2(new_n1083), .B1(new_n215), .B2(new_n725), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n777), .B1(new_n1084), .B2(new_n793), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n711), .A2(new_n846), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n785), .B1(new_n841), .B2(new_n799), .C1(new_n346), .C2(new_n840), .ZN(new_n1087));
  INV_X1    g0887(.A(G150), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n798), .A2(new_n1088), .B1(new_n815), .B2(new_n213), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT112), .Z(new_n1090));
  AOI22_X1  g0890(.A1(new_n806), .A2(G68), .B1(G97), .B2(new_n881), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n803), .B2(new_n344), .C1(new_n595), .C2(new_n818), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1087), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT113), .Z(new_n1094));
  OAI22_X1  g0894(.A1(new_n818), .A2(new_n832), .B1(new_n815), .B2(new_n829), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n810), .A2(G303), .B1(G322), .B2(new_n822), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n1067), .B2(new_n840), .C1(new_n886), .C2(new_n828), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT48), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT49), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n889), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n798), .A2(new_n842), .B1(new_n1103), .B2(new_n813), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(new_n785), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1094), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1085), .B(new_n1086), .C1(new_n791), .C2(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n776), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1047), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n726), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1109), .A2(new_n771), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(G393));
  NAND3_X1  g0914(.A1(new_n1040), .A2(KEYINPUT114), .A3(new_n1050), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1116), .B(new_n718), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1007), .A2(new_n846), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT115), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G311), .A2(new_n823), .B1(new_n822), .B2(G317), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT52), .Z(new_n1122));
  OAI22_X1  g0922(.A1(new_n827), .A2(new_n829), .B1(new_n832), .B2(new_n815), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n798), .A2(new_n839), .B1(new_n1103), .B2(new_n818), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n253), .A4(new_n814), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1122), .B(new_n1125), .C1(new_n522), .C2(new_n886), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n818), .A2(new_n213), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n798), .A2(new_n876), .B1(new_n813), .B2(new_n579), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(G68), .C2(new_n880), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1129), .A2(new_n785), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n346), .B2(new_n886), .C1(new_n344), .C2(new_n809), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G150), .A2(new_n822), .B1(new_n823), .B2(G159), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT51), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1126), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT116), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n897), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n786), .A2(new_n243), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n793), .B1(G97), .B2(new_n725), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n864), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1118), .A2(new_n776), .B1(new_n1120), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1115), .A2(new_n1111), .A3(new_n1117), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n726), .A3(new_n1051), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(G390));
  NOR2_X1   g0943(.A1(new_n942), .A2(new_n789), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n886), .A2(new_n1061), .B1(new_n809), .B2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT120), .Z(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n798), .A2(new_n1148), .B1(new_n813), .B2(new_n346), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n333), .B(new_n1149), .C1(G159), .C2(new_n819), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n815), .A2(new_n1088), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G128), .A2(new_n822), .B1(new_n823), .B2(G132), .ZN(new_n1153));
  AND4_X1   g0953(.A1(new_n1147), .A2(new_n1150), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n841), .A2(new_n832), .B1(new_n809), .B2(new_n502), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1127), .B1(G68), .B2(new_n881), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n829), .B2(new_n798), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n253), .B(new_n1157), .C1(G87), .C2(new_n880), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n215), .B2(new_n886), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1155), .B(new_n1159), .C1(G116), .C2(new_n823), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n791), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n777), .C1(new_n370), .C2(new_n872), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1144), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n753), .A2(G330), .A3(new_n859), .A4(new_n958), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT117), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n943), .B1(new_n947), .B2(new_n958), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n918), .B1(new_n982), .B2(new_n989), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n919), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1164), .A2(KEYINPUT117), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n940), .A2(new_n931), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n943), .B1(new_n1172), .B2(new_n930), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n766), .A2(new_n710), .A3(new_n859), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n946), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n958), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1171), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1165), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n982), .A2(new_n989), .B1(new_n320), .B2(new_n703), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n958), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1174), .B2(new_n946), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1180), .A2(new_n1182), .B1(KEYINPUT117), .B2(new_n1164), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1165), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1183), .A2(new_n1169), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1163), .B1(new_n1187), .B2(new_n776), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n753), .A2(G330), .A3(new_n859), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1181), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1164), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n947), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT119), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n946), .A3(new_n1164), .A4(new_n1174), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n753), .A2(new_n669), .A3(G330), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT118), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n965), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1175), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1200), .A2(KEYINPUT119), .A3(new_n1164), .A4(new_n1190), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1195), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n726), .B1(new_n1187), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1178), .B2(new_n1185), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1188), .B1(new_n1203), .B2(new_n1205), .ZN(G378));
  INV_X1    g1006(.A(KEYINPUT123), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n362), .A2(new_n367), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n904), .A2(new_n352), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1210), .B(new_n1211), .Z(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n990), .A2(G330), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n931), .A2(new_n969), .B1(new_n974), .B2(KEYINPUT109), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT40), .B1(new_n1215), .B2(new_n977), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n967), .B1(new_n941), .B2(new_n981), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT122), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n980), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1213), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1218), .B2(new_n980), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(new_n1212), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1207), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(KEYINPUT124), .B(new_n961), .C1(new_n942), .C2(new_n943), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n944), .B2(new_n962), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1224), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1204), .A2(new_n1199), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1228), .B(new_n1207), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n963), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1218), .A2(new_n980), .A3(new_n1219), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1212), .B1(new_n1238), .B2(new_n1222), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1217), .A2(new_n1213), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n963), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1234), .B1(new_n1204), .B2(new_n1199), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n727), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1235), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1230), .A2(new_n776), .A3(new_n1232), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n864), .B1(new_n346), .B2(new_n871), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n806), .A2(G137), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n819), .A2(G150), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n815), .A2(new_n1145), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n823), .A2(G128), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n841), .B2(new_n1148), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1252), .B(new_n1254), .C1(G132), .C2(new_n834), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G33), .A2(G41), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT121), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n813), .A2(new_n799), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(G124), .C2(new_n797), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(new_n1258), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G41), .B1(new_n819), .B2(G68), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n595), .B2(new_n827), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n798), .A2(new_n832), .B1(new_n815), .B2(new_n213), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n813), .A2(new_n402), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1266), .A2(new_n785), .A3(new_n1267), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n215), .B2(new_n840), .C1(new_n527), .C2(new_n841), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1265), .B(new_n1269), .C1(G97), .C2(new_n834), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1270), .A2(KEYINPUT58), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(KEYINPUT58), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n346), .B(new_n1260), .C1(new_n785), .C2(G41), .ZN(new_n1273));
  AND4_X1   g1073(.A1(new_n1263), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n1248), .B1(new_n897), .B2(new_n1274), .C1(new_n1213), .C2(new_n789), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1247), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1246), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(G375));
  NAND2_X1  g1078(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n965), .B2(new_n1198), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1029), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1195), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1195), .A2(new_n776), .A3(new_n1201), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n777), .B1(G68), .B2(new_n872), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G150), .A2(new_n806), .B1(new_n797), .B2(G128), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n346), .B2(new_n818), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1267), .B(new_n1287), .C1(G159), .C2(new_n880), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n886), .B2(new_n1145), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n822), .A2(G132), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1290), .B(new_n785), .C1(new_n840), .C2(new_n1061), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n798), .A2(new_n522), .B1(new_n815), .B2(new_n502), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n595), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n819), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n1294), .B1(new_n215), .B2(new_n809), .C1(new_n886), .C2(new_n1103), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT125), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n333), .B1(new_n813), .B2(new_n213), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n822), .A2(G294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n1298), .B1(new_n1296), .B2(new_n1297), .C1(new_n832), .C2(new_n840), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1289), .A2(new_n1291), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1285), .B1(new_n1300), .B2(new_n791), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n958), .B2(new_n789), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1284), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1283), .A2(new_n1303), .ZN(G381));
  OR4_X1    g1104(.A1(G396), .A2(G384), .A3(G381), .A4(G393), .ZN(new_n1305));
  NOR4_X1   g1105(.A1(new_n1305), .A2(G387), .A3(G390), .A4(G378), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1277), .ZN(G407));
  INV_X1    g1107(.A(G378), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n702), .A2(G213), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(KEYINPUT126), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1277), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(G407), .A2(G213), .A3(new_n1311), .ZN(G409));
  INV_X1    g1112(.A(new_n1276), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1245), .A2(G378), .A3(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1281), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1237), .A2(new_n1241), .A3(new_n776), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1275), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1316), .B2(new_n1275), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1308), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1314), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1282), .A2(KEYINPUT60), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n726), .B1(new_n1280), .B2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1280), .A2(new_n1323), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1303), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(G384), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G384), .B(new_n1303), .C1(new_n1324), .C2(new_n1325), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1322), .A2(new_n1309), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(G387), .A2(new_n1142), .A3(new_n1140), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(G393), .B(new_n848), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(G390), .A2(new_n1053), .A3(new_n1076), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1335), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1336), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1338), .A2(new_n1339), .A3(KEYINPUT61), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1322), .A2(new_n1309), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n702), .A2(G213), .A3(G2897), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1328), .A2(new_n1329), .A3(new_n1342), .ZN(new_n1343));
  AOI22_X1  g1143(.A1(new_n1328), .A2(new_n1329), .B1(G2897), .B2(new_n1310), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1341), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1310), .B1(new_n1314), .B2(new_n1321), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1334), .A2(new_n1340), .A3(new_n1347), .A4(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT61), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1351), .B1(new_n1348), .B2(new_n1345), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1332), .A2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1348), .A2(KEYINPUT62), .A3(new_n1331), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1352), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1350), .B1(new_n1356), .B2(new_n1357), .ZN(G405));
  OAI21_X1  g1158(.A(new_n1308), .B1(new_n1246), .B2(new_n1276), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1314), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1331), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1359), .A2(new_n1330), .A3(new_n1314), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1357), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1361), .A2(new_n1357), .A3(new_n1362), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(G402));
endmodule


