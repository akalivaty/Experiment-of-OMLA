//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n463), .A2(new_n465), .A3(new_n469), .A4(G125), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n463), .A2(new_n465), .A3(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n463), .A2(new_n465), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n482), .A2(KEYINPUT69), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT69), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n479), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n480), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n484), .A2(new_n485), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n462), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(KEYINPUT70), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(new_n480), .B2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(new_n494), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT3), .B(G2104), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(G126), .A3(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n480), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n501), .A2(KEYINPUT4), .A3(G138), .A4(new_n480), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n500), .A2(new_n502), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(new_n510), .A3(new_n512), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  INV_X1    g098(.A(new_n518), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  INV_X1    g100(.A(new_n520), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n515), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n518), .A2(new_n535), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n510), .A2(new_n512), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT71), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n545), .A3(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT72), .B(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n526), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n524), .A2(G81), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT73), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n547), .A2(new_n553), .A3(new_n549), .A4(new_n550), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(KEYINPUT76), .B(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n540), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n524), .A2(G91), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n526), .A2(KEYINPUT9), .A3(G53), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n520), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT75), .B1(new_n567), .B2(new_n570), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n566), .B1(new_n573), .B2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  XNOR2_X1  g151(.A(new_n531), .B(KEYINPUT77), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n518), .A2(new_n579), .B1(new_n520), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT78), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(G651), .C1(new_n513), .C2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n540), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n590), .A2(KEYINPUT79), .A3(G651), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT79), .B1(new_n590), .B2(G651), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n513), .A2(G86), .A3(new_n517), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n518), .A2(new_n599), .B1(new_n520), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n540), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(KEYINPUT80), .A3(G651), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n602), .A2(new_n608), .A3(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n540), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(G54), .A2(new_n526), .B1(new_n613), .B2(G651), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n518), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT10), .B1(new_n518), .B2(new_n615), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G171), .ZN(G284));
  OAI21_X1  g196(.A(new_n620), .B1(new_n619), .B2(G171), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n619), .ZN(new_n623));
  INV_X1    g198(.A(G286), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n619), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n619), .ZN(G280));
  INV_X1    g201(.A(new_n618), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(G559), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(G860), .B2(new_n629), .ZN(G148));
  INV_X1    g205(.A(new_n555), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n619), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n618), .A2(new_n628), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n619), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n481), .A2(G123), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n486), .A2(G135), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n480), .B2(G111), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n664), .B2(new_n665), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n666), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n672), .B(new_n675), .Z(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AOI21_X1  g256(.A(KEYINPUT85), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT85), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n684), .A2(new_n685), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(new_n681), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n678), .A3(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n687), .B(new_n690), .C1(new_n685), .C2(new_n684), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT86), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1981), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n696), .B(new_n698), .Z(G229));
  MUX2_X1   g274(.A(G6), .B(G305), .S(G16), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(G1971), .Z(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n702), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT34), .Z(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1986), .Z(new_n715));
  AOI22_X1  g290(.A1(G119), .A2(new_n481), .B1(new_n486), .B2(G131), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(new_n480), .B2(G107), .ZN(new_n717));
  NOR2_X1   g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT89), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT88), .B(G29), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n720), .S(new_n721), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n713), .A2(new_n715), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT36), .ZN(new_n726));
  INV_X1    g301(.A(new_n721), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n727), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT29), .B(G2090), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n627), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G4), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT97), .B(G2078), .ZN(new_n736));
  NAND2_X1  g311(.A1(G164), .A2(new_n721), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G27), .B2(new_n721), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(G5), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G171), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n739), .B1(new_n740), .B2(new_n743), .C1(new_n736), .C2(new_n738), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G32), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n486), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n481), .A2(G129), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n480), .A2(G105), .A3(G2104), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND4_X1  g327(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n640), .A2(new_n727), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n703), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n703), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1966), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n743), .A2(new_n740), .B1(new_n755), .B2(new_n756), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(G28), .ZN(new_n766));
  INV_X1    g341(.A(G29), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n762), .B(new_n769), .C1(new_n734), .C2(new_n733), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n746), .A2(new_n757), .A3(new_n759), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  INV_X1    g347(.A(G127), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n479), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2105), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n486), .A2(G139), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  AND3_X1   g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G29), .B2(G33), .ZN(new_n783));
  INV_X1    g358(.A(G2072), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT95), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n727), .A2(KEYINPUT28), .A3(G26), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n481), .A2(G128), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n486), .A2(G140), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n767), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT28), .B1(new_n727), .B2(G26), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT24), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n727), .B1(new_n800), .B2(G34), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(G34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n477), .B2(new_n767), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  INV_X1    g383(.A(G2084), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n783), .A2(new_n784), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n786), .A2(new_n799), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n703), .A2(KEYINPUT23), .A3(G20), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT23), .ZN(new_n814));
  INV_X1    g389(.A(G20), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G299), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n813), .B(new_n816), .C1(new_n817), .C2(new_n703), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1956), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n771), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n726), .A2(new_n731), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n808), .A2(new_n809), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT96), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n703), .A2(G19), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n555), .B2(new_n703), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT90), .Z(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1341), .Z(new_n827));
  NOR3_X1   g402(.A1(new_n821), .A2(new_n823), .A3(new_n827), .ZN(G311));
  INV_X1    g403(.A(new_n820), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n823), .ZN(new_n833));
  INV_X1    g408(.A(new_n827), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n731), .ZN(G150));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n540), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G651), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  INV_X1    g417(.A(G55), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n518), .A2(new_n842), .B1(new_n520), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n627), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT39), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n845), .B1(new_n552), .B2(new_n554), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n845), .A2(new_n551), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n852), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n848), .B1(new_n856), .B2(G860), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT100), .ZN(G145));
  NAND2_X1  g433(.A1(new_n481), .A2(G130), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n486), .A2(G142), .ZN(new_n860));
  NOR2_X1   g435(.A1(G106), .A2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(new_n480), .B2(G118), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n720), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n781), .A2(new_n792), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n793), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n507), .B(new_n643), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n866), .B2(new_n868), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n871), .A2(new_n872), .A3(new_n754), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n868), .ZN(new_n874));
  INV_X1    g449(.A(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n753), .B1(new_n876), .B2(new_n870), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n865), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n754), .B1(new_n871), .B2(new_n872), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n753), .A3(new_n870), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n864), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n477), .B(new_n640), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n490), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT101), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n878), .A2(new_n884), .A3(new_n881), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n882), .A2(new_n891), .A3(new_n885), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT102), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n887), .A2(new_n890), .A3(new_n895), .A4(new_n892), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(KEYINPUT40), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT40), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(G395));
  NAND2_X1  g474(.A1(new_n846), .A2(new_n619), .ZN(new_n900));
  NAND2_X1  g475(.A1(G299), .A2(new_n618), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n627), .B(new_n566), .C1(new_n574), .C2(new_n573), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(KEYINPUT103), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n902), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT41), .B1(new_n901), .B2(new_n902), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n855), .B(new_n633), .ZN(new_n912));
  MUX2_X1   g487(.A(new_n907), .B(new_n911), .S(new_n912), .Z(new_n913));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(G305), .B(G303), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n708), .A2(G290), .ZN(new_n916));
  NAND4_X1  g491(.A1(G288), .A2(new_n602), .A3(new_n608), .A4(new_n609), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT104), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n915), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G305), .B(G166), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n914), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n925), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  INV_X1    g503(.A(new_n921), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n923), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n915), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n926), .B1(new_n933), .B2(new_n914), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n913), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n900), .B1(new_n935), .B2(new_n619), .ZN(G295));
  OAI21_X1  g511(.A(new_n900), .B1(new_n935), .B2(new_n619), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  INV_X1    g514(.A(new_n903), .ZN(new_n940));
  NOR2_X1   g515(.A1(G171), .A2(new_n531), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(G286), .B2(G171), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n853), .B2(new_n854), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n942), .A2(new_n853), .A3(new_n854), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n855), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n910), .A2(new_n948), .A3(new_n943), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT105), .B1(new_n922), .B2(new_n925), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n930), .A2(new_n928), .A3(new_n931), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n939), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n933), .A2(KEYINPUT106), .A3(new_n949), .A4(new_n946), .ZN(new_n955));
  INV_X1    g530(.A(new_n949), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n907), .B1(new_n948), .B2(new_n943), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n889), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n950), .A2(new_n953), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(new_n955), .A3(new_n962), .A4(new_n889), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n963), .B2(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n938), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n960), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT126), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT70), .B1(new_n493), .B2(new_n495), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n498), .A2(new_n497), .A3(new_n494), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n502), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n505), .A2(new_n506), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n983), .B(new_n475), .C1(new_n471), .C2(G2105), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n507), .A2(new_n985), .A3(new_n976), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n982), .A2(new_n809), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n985), .B1(new_n507), .B2(new_n976), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n472), .A2(G40), .A3(new_n476), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(KEYINPUT116), .A3(new_n809), .A4(new_n986), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT110), .B(G8), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n531), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n981), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n984), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1966), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1001), .A2(new_n997), .A3(new_n1002), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n994), .B(new_n996), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1001), .A2(new_n997), .A3(new_n1002), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(new_n989), .B2(new_n993), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n996), .A2(G8), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1005), .B(KEYINPUT51), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  INV_X1    g587(.A(new_n995), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1012), .B(new_n996), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1011), .A2(KEYINPUT122), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT122), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1015), .A2(new_n1016), .A3(KEYINPUT62), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT109), .B(G1971), .Z(new_n1018));
  NAND2_X1  g593(.A1(new_n1001), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2090), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT55), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n986), .A2(KEYINPUT113), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n507), .A2(new_n1030), .A3(new_n985), .A4(new_n976), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n992), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1032), .A2(new_n1019), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1027), .B(new_n1025), .C1(new_n1033), .C2(new_n1013), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1024), .B(KEYINPUT55), .Z(new_n1035));
  AOI21_X1  g610(.A(new_n1013), .B1(new_n1032), .B2(new_n1019), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1026), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G2078), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n999), .A2(new_n1039), .A3(new_n984), .A4(new_n1000), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1040), .A2(new_n1041), .B1(new_n1021), .B2(new_n740), .ZN(new_n1042));
  NOR2_X1   g617(.A1(KEYINPUT123), .A2(KEYINPUT53), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(G301), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g621(.A(new_n981), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1013), .B1(new_n1047), .B2(new_n984), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n708), .A2(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1048), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n596), .A2(KEYINPUT111), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n590), .A2(G651), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT79), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n590), .A2(KEYINPUT79), .A3(G651), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n594), .A2(new_n1061), .A3(new_n595), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(G1981), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1062), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n594), .B2(new_n595), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1069), .B2(new_n593), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n597), .A2(new_n1059), .A3(new_n1066), .A4(new_n1060), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT112), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1065), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1055), .B1(new_n1073), .B2(KEYINPUT49), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1065), .B(new_n1075), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1050), .B(new_n1054), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1038), .A2(new_n1045), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n975), .B1(new_n1017), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1078), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1011), .A2(KEYINPUT122), .A3(new_n1014), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT126), .B(new_n1080), .C1(new_n1085), .C2(KEYINPUT62), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1079), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT56), .B(G2072), .Z(new_n1090));
  OR3_X1    g665(.A1(new_n1001), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n992), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1092));
  INV_X1    g667(.A(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1089), .B1(new_n1001), .B2(new_n1090), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n817), .A2(new_n1097), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1097), .A2(new_n566), .A3(new_n570), .A4(new_n567), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1091), .A2(new_n1094), .A3(new_n1101), .A4(new_n1095), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1105), .A3(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1001), .A2(G1996), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n991), .B2(new_n981), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n631), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT59), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1021), .A2(new_n734), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n991), .A2(new_n981), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n798), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n627), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT120), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1021), .A2(new_n734), .B1(new_n1114), .B2(new_n798), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(KEYINPUT60), .A4(new_n618), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT119), .B1(new_n1116), .B2(new_n627), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1116), .A2(new_n1123), .A3(new_n627), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1125), .A2(KEYINPUT121), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT121), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1107), .B(new_n1112), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1100), .B1(new_n618), .B2(new_n1119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1102), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT124), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1042), .A2(new_n1044), .A3(G301), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1045), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1137), .A2(KEYINPUT54), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT54), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1141), .A2(new_n1143), .A3(new_n1038), .A4(new_n1077), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1133), .B1(new_n1134), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1143), .A2(new_n1038), .A3(new_n1077), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1085), .A2(KEYINPUT125), .A3(new_n1146), .A4(new_n1141), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1132), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1077), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n994), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(new_n624), .A3(new_n995), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(KEYINPUT63), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1026), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1050), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1048), .A3(new_n1076), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .A4(new_n1053), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT63), .B1(new_n1161), .B2(new_n1151), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1051), .A3(new_n708), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1071), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1048), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT117), .B1(new_n1156), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1009), .A2(G286), .A3(new_n1013), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1168), .A2(new_n1077), .A3(new_n1157), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1169), .A2(KEYINPUT63), .B1(new_n1048), .B2(new_n1164), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1026), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1170), .B(new_n1171), .C1(new_n1149), .C2(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1088), .A2(new_n1148), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n999), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n984), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT108), .Z(new_n1178));
  XNOR2_X1  g753(.A(new_n792), .B(new_n798), .ZN(new_n1179));
  INV_X1    g754(.A(G1996), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(new_n754), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1177), .A2(G1996), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n754), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n720), .B(new_n723), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1178), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1177), .ZN(new_n1189));
  XNOR2_X1  g764(.A(G290), .B(G1986), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1175), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1185), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1193), .A2(new_n723), .A3(new_n720), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n792), .A2(G2067), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1178), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1183), .B(KEYINPUT46), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1179), .A2(new_n754), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n1178), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT47), .Z(new_n1200));
  NAND2_X1  g775(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1177), .A2(G1986), .A3(G290), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  XOR2_X1   g778(.A(new_n1188), .B(KEYINPUT127), .Z(new_n1204));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1192), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g781(.A1(G401), .A2(G227), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n894), .B2(new_n896), .ZN(new_n1209));
  INV_X1    g783(.A(G229), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n460), .B1(new_n969), .B2(new_n970), .ZN(new_n1211));
  AND3_X1   g785(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(G308));
  NAND3_X1  g786(.A1(new_n1209), .A2(new_n1211), .A3(new_n1210), .ZN(G225));
endmodule


