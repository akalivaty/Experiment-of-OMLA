//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT69), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n461), .B2(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n467), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n468), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n471), .B2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n473), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n462), .C1(new_n472), .C2(new_n473), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n462), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT71), .B1(new_n478), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n489), .A2(new_n462), .A3(G138), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n461), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n481), .B2(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(new_n511), .A3(G62), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n502), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n508), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n513), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(KEYINPUT74), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(G543), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT75), .B(G51), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(new_n515), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n526), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  INV_X1    g109(.A(new_n530), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n536), .B1(new_n537), .B2(new_n524), .C1(new_n502), .C2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n505), .A2(new_n507), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n502), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n520), .A2(G543), .A3(new_n523), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G43), .B1(new_n535), .B2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n542), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n535), .B2(G91), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n520), .A2(G53), .A3(G543), .A4(new_n523), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT77), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n548), .A2(new_n566), .A3(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n560), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT78), .ZN(new_n571));
  INV_X1    g146(.A(new_n560), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT77), .B1(new_n562), .B2(new_n563), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n567), .A2(new_n565), .A3(new_n568), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n571), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G166), .ZN(G303));
  OAI21_X1  g154(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  INV_X1    g156(.A(G49), .ZN(new_n582));
  OAI221_X1 g157(.A(new_n580), .B1(new_n581), .B2(new_n530), .C1(new_n524), .C2(new_n582), .ZN(G288));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n505), .B2(new_n507), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n505), .B2(new_n507), .ZN(new_n589));
  AND2_X1   g164(.A1(G48), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n515), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n542), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n520), .A2(G47), .A3(G543), .A4(new_n523), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n535), .A2(G85), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT79), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n596), .A2(new_n598), .A3(new_n601), .A4(new_n597), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n535), .A2(G92), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT80), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n542), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n548), .A2(G54), .B1(new_n612), .B2(G651), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(G286), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G299), .B(KEYINPUT81), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(G297));
  AOI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n550), .A2(new_n618), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n614), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n461), .A2(new_n464), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n479), .A2(G135), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT82), .Z(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT83), .B1(new_n462), .B2(G111), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G2104), .A3(new_n638), .ZN(new_n639));
  OR3_X1    g214(.A1(new_n462), .A2(KEYINPUT83), .A3(G111), .ZN(new_n640));
  AOI22_X1  g215(.A1(G123), .A2(new_n481), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n631), .A2(new_n632), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n641), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n633), .A2(new_n642), .A3(new_n643), .A4(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n652), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n632), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n636), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n676), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT84), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  OR3_X1    g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n693), .B1(new_n692), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G23), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G288), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(G166), .A2(G16), .ZN(new_n703));
  OR2_X1    g278(.A1(G16), .A2(G22), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n703), .A2(G1971), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT34), .ZN(new_n707));
  INV_X1    g282(.A(G305), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G16), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n710));
  OR2_X1    g285(.A1(G6), .A2(G16), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  OAI21_X1  g288(.A(G1981), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(new_n711), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT32), .ZN(new_n716));
  INV_X1    g291(.A(G1981), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n703), .A2(new_n704), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n706), .A2(new_n707), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n698), .B1(new_n600), .B2(new_n602), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n698), .A2(G24), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT86), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n726), .A2(KEYINPUT86), .A3(new_n727), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n726), .A2(KEYINPUT86), .A3(new_n727), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n732), .A2(G1986), .A3(new_n728), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n479), .A2(G131), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n481), .A2(G119), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n462), .A2(G107), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT85), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n734), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n724), .A2(new_n731), .A3(new_n733), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT87), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n733), .A2(new_n744), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n747), .A2(new_n748), .A3(new_n724), .A4(new_n731), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n706), .A2(new_n720), .A3(new_n723), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT34), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n746), .A2(new_n749), .B1(KEYINPUT34), .B2(new_n752), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT36), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n750), .A2(new_n758), .A3(new_n753), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n750), .A2(new_n753), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT88), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n757), .A2(new_n758), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n763), .A2(new_n755), .A3(KEYINPUT36), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n761), .B2(new_n765), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT30), .B(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(new_n734), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n734), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n734), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT29), .B(G2090), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n772), .B1(new_n774), .B2(new_n775), .C1(new_n644), .C2(new_n734), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n734), .A2(G32), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT92), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT26), .Z(new_n780));
  AOI22_X1  g355(.A1(new_n481), .A2(G129), .B1(G105), .B2(new_n464), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n479), .A2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(new_n734), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n776), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n734), .A2(G33), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(new_n462), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n479), .A2(G139), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2072), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n800), .B(new_n801), .C1(new_n774), .C2(new_n775), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n698), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n698), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G1966), .ZN(new_n805));
  INV_X1    g380(.A(new_n787), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n804), .A2(G1966), .B1(new_n785), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n788), .A2(new_n802), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G27), .A2(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2078), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT24), .ZN(new_n812));
  INV_X1    g387(.A(G34), .ZN(new_n813));
  AOI21_X1  g388(.A(G29), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G160), .B2(new_n734), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2084), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n808), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(G4), .A2(G16), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n615), .B2(G16), .ZN(new_n820));
  INV_X1    g395(.A(G1348), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n698), .A2(G5), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G171), .B2(new_n698), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT93), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1961), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n551), .A2(G16), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G16), .B2(G19), .ZN(new_n828));
  INV_X1    g403(.A(G1341), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n734), .A2(G26), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT28), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n479), .A2(G140), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n481), .A2(G128), .ZN(new_n835));
  OR2_X1    g410(.A1(G104), .A2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT91), .A4(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n833), .B1(new_n842), .B2(G29), .ZN(new_n843));
  INV_X1    g418(.A(G2067), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n830), .A2(new_n831), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n818), .A2(new_n822), .A3(new_n826), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n698), .A2(G20), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT94), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT23), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n571), .A2(new_n577), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(new_n698), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G1956), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n767), .A2(new_n768), .A3(new_n855), .ZN(G311));
  INV_X1    g431(.A(new_n768), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n854), .ZN(G150));
  AOI22_X1  g434(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n502), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT95), .B(G55), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n548), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n535), .A2(G93), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT98), .B(G860), .Z(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n550), .A2(KEYINPUT96), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n547), .A2(new_n871), .A3(new_n549), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n872), .A3(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n550), .A2(KEYINPUT96), .A3(new_n865), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n615), .A2(G559), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT97), .Z(new_n881));
  OAI21_X1  g456(.A(new_n867), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n869), .B1(new_n881), .B2(new_n882), .ZN(G145));
  NAND2_X1  g458(.A1(new_n479), .A2(G142), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  INV_X1    g463(.A(G118), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(G2105), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n481), .B2(G130), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n887), .B1(new_n886), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n630), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n886), .A2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT100), .ZN(new_n897));
  INV_X1    g472(.A(new_n630), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n741), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n741), .B1(new_n895), .B2(new_n899), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n797), .ZN(new_n904));
  NAND3_X1  g479(.A1(G164), .A2(new_n840), .A3(new_n841), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G164), .B1(new_n840), .B2(new_n841), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n842), .A2(new_n500), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n797), .A3(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n784), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n784), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n903), .A2(new_n915), .A3(KEYINPUT101), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT101), .B1(new_n903), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT102), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n913), .A2(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n895), .A2(new_n899), .ZN(new_n921));
  INV_X1    g496(.A(new_n741), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n900), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n903), .A2(new_n915), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n920), .B2(new_n924), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n916), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n919), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G160), .B(G162), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(new_n644), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n916), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n920), .B2(new_n924), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g516(.A(new_n626), .B(new_n875), .Z(new_n942));
  NAND2_X1  g517(.A1(G299), .A2(new_n615), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n851), .A2(new_n614), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT41), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n942), .A2(new_n946), .ZN(new_n950));
  NOR2_X1   g525(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n951));
  OR3_X1    g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n953));
  XNOR2_X1  g528(.A(G290), .B(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(G166), .B(KEYINPUT105), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(G288), .B(G305), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n955), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n951), .B1(new_n949), .B2(new_n950), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n952), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n952), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g543(.A(new_n967), .B1(G868), .B2(new_n866), .ZN(G331));
  INV_X1    g544(.A(new_n961), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n959), .ZN(new_n971));
  XOR2_X1   g546(.A(G301), .B(G286), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n875), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n948), .B2(new_n945), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n946), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n973), .ZN(new_n978));
  INV_X1    g553(.A(new_n945), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT41), .B1(new_n943), .B2(new_n944), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n962), .A3(new_n975), .ZN(new_n982));
  INV_X1    g557(.A(G37), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n977), .A2(new_n982), .A3(new_n986), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(G397));
  XNOR2_X1  g565(.A(new_n842), .B(new_n844), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n500), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n466), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT70), .B1(new_n475), .B2(G2105), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n467), .B(new_n462), .C1(new_n474), .C2(new_n468), .ZN(new_n998));
  OAI211_X1 g573(.A(G40), .B(new_n996), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n991), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n784), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n1000), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n741), .B(new_n743), .Z(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT108), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(KEYINPUT108), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1000), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(new_n725), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1009), .B(new_n1013), .C1(new_n1001), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n495), .B2(new_n499), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT50), .B(G1384), .C1(new_n495), .C2(new_n499), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n999), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G1961), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n999), .B1(KEYINPUT45), .B2(new_n1017), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n993), .A2(new_n1024), .A3(new_n994), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT109), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(KEYINPUT119), .A3(new_n1029), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1022), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1023), .A2(KEYINPUT53), .A3(new_n1026), .A4(new_n995), .ZN(new_n1035));
  AOI21_X1  g610(.A(G301), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1022), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n475), .A2(G2105), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1039));
  INV_X1    g614(.A(G40), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT120), .B(G2078), .ZN(new_n1041));
  NOR4_X1   g616(.A1(new_n466), .A2(new_n1029), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n995), .A2(new_n1038), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1028), .A2(KEYINPUT119), .A3(new_n1029), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT119), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1037), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(G171), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1016), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(G166), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1023), .A2(new_n1027), .A3(new_n1025), .ZN(new_n1055));
  INV_X1    g630(.A(G2090), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1055), .A2(new_n722), .B1(new_n1021), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1054), .B1(new_n1057), .B2(new_n1051), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1040), .B(new_n466), .C1(new_n471), .C2(new_n476), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1039), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1017), .A2(KEYINPUT109), .A3(KEYINPUT45), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1971), .B1(new_n1062), .B2(new_n1027), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G2090), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(new_n1053), .C1(new_n1063), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  OR2_X1    g644(.A1(G288), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(G8), .C1(new_n993), .C2(new_n999), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(G160), .A2(new_n1017), .A3(G40), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(G8), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1070), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n587), .A2(new_n591), .A3(new_n717), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G305), .A2(G1981), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT49), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n993), .B2(new_n999), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT110), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1072), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1076), .A2(KEYINPUT52), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1070), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1058), .A2(new_n1068), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1017), .A2(KEYINPUT45), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1060), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1064), .A2(new_n1100), .A3(new_n1059), .A4(new_n1065), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G286), .A2(G8), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1099), .A2(new_n1107), .A3(new_n1101), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(G286), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1104), .A2(new_n1051), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1106), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(new_n1105), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1096), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1048), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1037), .B(new_n1035), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT54), .B1(new_n1118), .B2(G171), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1034), .A2(new_n1120), .A3(new_n1043), .ZN(new_n1121));
  AOI21_X1  g696(.A(G301), .B1(new_n1046), .B2(KEYINPUT121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT122), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1121), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1048), .A4(new_n1116), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1074), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1055), .B2(G1996), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g708(.A1(KEYINPUT114), .A2(KEYINPUT59), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n551), .A4(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n551), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n560), .B(new_n1139), .C1(new_n562), .C2(new_n563), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n575), .B2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT112), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT112), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1143), .B(new_n1140), .C1(new_n575), .C2(new_n1139), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1021), .A2(G1956), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT56), .B(G2072), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1062), .A2(new_n1027), .A3(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT61), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n551), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1074), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n844), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1021), .B2(G1348), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1150), .A2(new_n1151), .B1(new_n1156), .B2(new_n614), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1156), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n615), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1138), .A2(new_n1149), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1148), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(KEYINPUT117), .A3(new_n1163), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT116), .B(KEYINPUT61), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1161), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1148), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1142), .A2(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1172), .A2(KEYINPUT113), .B1(new_n615), .B2(new_n1154), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT113), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1164), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1171), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1124), .A2(new_n1129), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1181), .A2(new_n1182), .B1(new_n717), .B2(new_n708), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1092), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1180), .A2(new_n1068), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1102), .A2(G8), .A3(G168), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n1096), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1187), .B1(new_n1096), .B2(new_n1186), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1185), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT62), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1113), .A2(new_n1193), .A3(new_n1115), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1118), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1096), .A2(new_n1195), .A3(G301), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1015), .B1(new_n1179), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT124), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1001), .B1(new_n991), .B2(new_n784), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n1202), .B2(new_n1201), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT47), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1000), .A2(new_n725), .A3(new_n600), .A4(new_n602), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT125), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT48), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1009), .A2(new_n1013), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1208), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n741), .A2(new_n743), .ZN(new_n1216));
  OAI22_X1  g791(.A1(new_n1008), .A2(new_n1216), .B1(G2067), .B2(new_n842), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n1218));
  AND3_X1   g793(.A1(new_n1217), .A2(new_n1218), .A3(new_n1000), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1218), .B1(new_n1217), .B2(new_n1000), .ZN(new_n1220));
  NOR3_X1   g795(.A1(new_n1215), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(KEYINPUT126), .B1(new_n1200), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1176), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1127), .A2(new_n1048), .A3(new_n1116), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1225), .B1(new_n1226), .B2(KEYINPUT122), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1198), .B1(new_n1227), .B2(new_n1129), .ZN(new_n1228));
  OAI211_X1 g803(.A(new_n1224), .B(new_n1221), .C1(new_n1228), .C2(new_n1015), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1223), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g805(.A(G319), .ZN(new_n1232));
  NOR3_X1   g806(.A1(G401), .A2(new_n1232), .A3(G227), .ZN(new_n1233));
  OAI21_X1  g807(.A(new_n1233), .B1(new_n695), .B2(new_n696), .ZN(new_n1234));
  AOI21_X1  g808(.A(new_n1234), .B1(new_n936), .B2(new_n939), .ZN(new_n1235));
  AND3_X1   g809(.A1(new_n988), .A2(KEYINPUT127), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g810(.A(KEYINPUT127), .B1(new_n988), .B2(new_n1235), .ZN(new_n1237));
  NOR2_X1   g811(.A1(new_n1236), .A2(new_n1237), .ZN(G308));
  NAND2_X1  g812(.A1(new_n988), .A2(new_n1235), .ZN(G225));
endmodule


