

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595;

  XNOR2_X1 U326 ( .A(n302), .B(KEYINPUT72), .ZN(n303) );
  INV_X1 U327 ( .A(KEYINPUT55), .ZN(n490) );
  INV_X1 U328 ( .A(n382), .ZN(n311) );
  XNOR2_X1 U329 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U330 ( .A(n430), .B(n429), .ZN(n542) );
  XOR2_X1 U331 ( .A(n365), .B(n364), .Z(n294) );
  XOR2_X1 U332 ( .A(KEYINPUT99), .B(n470), .Z(n295) );
  XNOR2_X1 U333 ( .A(n313), .B(n312), .ZN(n409) );
  INV_X1 U334 ( .A(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U335 ( .A(n463), .B(KEYINPUT98), .ZN(n464) );
  XNOR2_X1 U336 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .Z(n356) );
  XNOR2_X1 U338 ( .A(n356), .B(n355), .ZN(n357) );
  INV_X1 U339 ( .A(KEYINPUT94), .ZN(n419) );
  XNOR2_X1 U340 ( .A(n423), .B(n357), .ZN(n359) );
  XNOR2_X1 U341 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U342 ( .A(n304), .B(n303), .ZN(n308) );
  XNOR2_X1 U343 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U344 ( .A(n366), .B(n294), .ZN(n367) );
  XNOR2_X1 U345 ( .A(n422), .B(n311), .ZN(n312) );
  XNOR2_X1 U346 ( .A(n368), .B(n367), .ZN(n371) );
  XNOR2_X1 U347 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U348 ( .A(G218GAT), .ZN(n458) );
  NOR2_X1 U349 ( .A1(n467), .A2(n456), .ZN(n593) );
  XNOR2_X1 U350 ( .A(KEYINPUT93), .B(n471), .ZN(n566) );
  INV_X1 U351 ( .A(G36GAT), .ZN(n483) );
  XNOR2_X1 U352 ( .A(n458), .B(KEYINPUT62), .ZN(n459) );
  XNOR2_X1 U353 ( .A(n498), .B(G190GAT), .ZN(n499) );
  XNOR2_X1 U354 ( .A(n483), .B(KEYINPUT104), .ZN(n484) );
  XNOR2_X1 U355 ( .A(n460), .B(n459), .ZN(G1355GAT) );
  XNOR2_X1 U356 ( .A(n500), .B(n499), .ZN(G1351GAT) );
  XNOR2_X1 U357 ( .A(n485), .B(n484), .ZN(G1329GAT) );
  XOR2_X1 U358 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n297) );
  XNOR2_X1 U359 ( .A(KEYINPUT9), .B(G92GAT), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U361 ( .A(KEYINPUT71), .B(KEYINPUT11), .Z(n299) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G134GAT), .Z(n439) );
  XNOR2_X1 U363 ( .A(n439), .B(n356), .ZN(n298) );
  XNOR2_X1 U364 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U365 ( .A(n301), .B(n300), .Z(n304) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U367 ( .A(G106GAT), .B(G162GAT), .Z(n306) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(KEYINPUT70), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n319) );
  XOR2_X1 U370 ( .A(n319), .B(KEYINPUT64), .Z(n307) );
  XNOR2_X1 U371 ( .A(n308), .B(n307), .ZN(n313) );
  XOR2_X1 U372 ( .A(G36GAT), .B(G190GAT), .Z(n309) );
  XOR2_X1 U373 ( .A(G218GAT), .B(n309), .Z(n422) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n310), .B(KEYINPUT7), .ZN(n382) );
  XNOR2_X1 U376 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n314) );
  XOR2_X1 U377 ( .A(n409), .B(n314), .Z(n478) );
  XOR2_X1 U378 ( .A(KEYINPUT68), .B(G78GAT), .Z(n369) );
  XOR2_X1 U379 ( .A(KEYINPUT24), .B(n369), .Z(n318) );
  XOR2_X1 U380 ( .A(G211GAT), .B(KEYINPUT84), .Z(n316) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n315) );
  XNOR2_X1 U382 ( .A(n316), .B(n315), .ZN(n426) );
  XNOR2_X1 U383 ( .A(G218GAT), .B(n426), .ZN(n317) );
  XNOR2_X1 U384 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U385 ( .A(n319), .B(G22GAT), .Z(n321) );
  NAND2_X1 U386 ( .A1(G228GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U387 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U388 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U389 ( .A(KEYINPUT3), .B(G155GAT), .Z(n325) );
  XNOR2_X1 U390 ( .A(KEYINPUT2), .B(G148GAT), .ZN(n324) );
  XNOR2_X1 U391 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U392 ( .A(G141GAT), .B(n326), .ZN(n454) );
  XOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT85), .Z(n328) );
  XNOR2_X1 U394 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U396 ( .A(n454), .B(n329), .Z(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n486) );
  XOR2_X1 U398 ( .A(KEYINPUT82), .B(KEYINPUT79), .Z(n333) );
  XNOR2_X1 U399 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n332) );
  XNOR2_X1 U400 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U401 ( .A(G99GAT), .B(G134GAT), .Z(n335) );
  XOR2_X1 U402 ( .A(KEYINPUT0), .B(G127GAT), .Z(n443) );
  XNOR2_X1 U403 ( .A(n443), .B(KEYINPUT83), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U405 ( .A(n337), .B(n336), .Z(n339) );
  NAND2_X1 U406 ( .A1(G227GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U408 ( .A(G120GAT), .B(G190GAT), .Z(n341) );
  XNOR2_X1 U409 ( .A(G43GAT), .B(G15GAT), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n351) );
  XOR2_X1 U412 ( .A(KEYINPUT80), .B(KEYINPUT17), .Z(n345) );
  XNOR2_X1 U413 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(n346), .ZN(n429) );
  XOR2_X1 U416 ( .A(G183GAT), .B(G176GAT), .Z(n348) );
  XNOR2_X1 U417 ( .A(KEYINPUT20), .B(G71GAT), .ZN(n347) );
  XNOR2_X1 U418 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U419 ( .A(n429), .B(n349), .Z(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n555) );
  INV_X1 U421 ( .A(n555), .ZN(n545) );
  NAND2_X1 U422 ( .A1(n486), .A2(n545), .ZN(n352) );
  XNOR2_X1 U423 ( .A(n352), .B(KEYINPUT26), .ZN(n467) );
  XOR2_X1 U424 ( .A(G64GAT), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n423) );
  AND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  INV_X1 U428 ( .A(KEYINPUT33), .ZN(n358) );
  NAND2_X1 U429 ( .A1(n359), .A2(n358), .ZN(n362) );
  INV_X1 U430 ( .A(n359), .ZN(n360) );
  NAND2_X1 U431 ( .A1(n360), .A2(KEYINPUT33), .ZN(n361) );
  NAND2_X1 U432 ( .A1(n362), .A2(n361), .ZN(n368) );
  XNOR2_X1 U433 ( .A(G71GAT), .B(KEYINPUT67), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n363), .B(KEYINPUT13), .ZN(n396) );
  XNOR2_X1 U435 ( .A(n396), .B(KEYINPUT69), .ZN(n366) );
  XOR2_X1 U436 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n365) );
  XNOR2_X1 U437 ( .A(G148GAT), .B(G106GAT), .ZN(n364) );
  XOR2_X1 U438 ( .A(G120GAT), .B(G57GAT), .Z(n450) );
  XNOR2_X1 U439 ( .A(n369), .B(n450), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n590) );
  XOR2_X1 U441 ( .A(KEYINPUT41), .B(n590), .Z(n523) );
  XOR2_X1 U442 ( .A(G197GAT), .B(G36GAT), .Z(n373) );
  XNOR2_X1 U443 ( .A(G50GAT), .B(G29GAT), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U445 ( .A(KEYINPUT29), .B(G8GAT), .Z(n375) );
  XNOR2_X1 U446 ( .A(G169GAT), .B(G141GAT), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U448 ( .A(n377), .B(n376), .ZN(n386) );
  XOR2_X1 U449 ( .A(G113GAT), .B(G1GAT), .Z(n451) );
  XNOR2_X1 U450 ( .A(G22GAT), .B(G15GAT), .ZN(n378) );
  XNOR2_X1 U451 ( .A(n378), .B(KEYINPUT66), .ZN(n388) );
  XOR2_X1 U452 ( .A(n451), .B(n388), .Z(n380) );
  NAND2_X1 U453 ( .A1(G229GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U454 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U455 ( .A(n381), .B(KEYINPUT30), .Z(n384) );
  XNOR2_X1 U456 ( .A(n382), .B(KEYINPUT65), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U458 ( .A(n386), .B(n385), .Z(n585) );
  AND2_X1 U459 ( .A1(n523), .A2(n585), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n387), .B(KEYINPUT46), .ZN(n407) );
  XOR2_X1 U461 ( .A(n388), .B(G64GAT), .Z(n390) );
  NAND2_X1 U462 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U463 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U464 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n392) );
  XNOR2_X1 U465 ( .A(KEYINPUT14), .B(KEYINPUT76), .ZN(n391) );
  XNOR2_X1 U466 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U467 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U468 ( .A(G8GAT), .B(G183GAT), .ZN(n395) );
  XNOR2_X1 U469 ( .A(n395), .B(KEYINPUT74), .ZN(n425) );
  XNOR2_X1 U470 ( .A(n396), .B(n425), .ZN(n397) );
  XNOR2_X1 U471 ( .A(n398), .B(n397), .ZN(n406) );
  XOR2_X1 U472 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n400) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U474 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U475 ( .A(G78GAT), .B(G211GAT), .Z(n402) );
  XNOR2_X1 U476 ( .A(G127GAT), .B(G155GAT), .ZN(n401) );
  XNOR2_X1 U477 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U478 ( .A(n404), .B(n403), .Z(n405) );
  XOR2_X1 U479 ( .A(n406), .B(n405), .Z(n577) );
  INV_X1 U480 ( .A(n577), .ZN(n594) );
  NOR2_X1 U481 ( .A1(n407), .A2(n594), .ZN(n408) );
  XNOR2_X1 U482 ( .A(n408), .B(KEYINPUT117), .ZN(n410) );
  NOR2_X1 U483 ( .A1(n410), .A2(n409), .ZN(n411) );
  XOR2_X1 U484 ( .A(KEYINPUT47), .B(n411), .Z(n417) );
  NOR2_X1 U485 ( .A1(n577), .A2(n478), .ZN(n412) );
  XNOR2_X1 U486 ( .A(KEYINPUT45), .B(n412), .ZN(n414) );
  NOR2_X1 U487 ( .A1(n590), .A2(n585), .ZN(n413) );
  AND2_X1 U488 ( .A1(n414), .A2(n413), .ZN(n415) );
  XNOR2_X1 U489 ( .A(n415), .B(KEYINPUT118), .ZN(n416) );
  NOR2_X1 U490 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U491 ( .A(n418), .B(KEYINPUT48), .ZN(n553) );
  NAND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n420) );
  XOR2_X1 U493 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n542), .B(KEYINPUT122), .ZN(n431) );
  NOR2_X1 U497 ( .A1(n553), .A2(n431), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n432), .B(KEYINPUT54), .ZN(n489) );
  XOR2_X1 U499 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n434) );
  XNOR2_X1 U500 ( .A(KEYINPUT89), .B(KEYINPUT91), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U502 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n436) );
  XNOR2_X1 U503 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n435) );
  XNOR2_X1 U504 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U505 ( .A(n438), .B(n437), .Z(n445) );
  XOR2_X1 U506 ( .A(n439), .B(KEYINPUT87), .Z(n441) );
  NAND2_X1 U507 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U508 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U509 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U511 ( .A(KEYINPUT90), .B(KEYINPUT86), .Z(n447) );
  XNOR2_X1 U512 ( .A(G162GAT), .B(G85GAT), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U514 ( .A(n449), .B(n448), .Z(n453) );
  XNOR2_X1 U515 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n471) );
  NAND2_X1 U518 ( .A1(n489), .A2(n566), .ZN(n456) );
  INV_X1 U519 ( .A(n593), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n478), .A2(n457), .ZN(n460) );
  INV_X1 U521 ( .A(n585), .ZN(n570) );
  NOR2_X1 U522 ( .A1(n570), .A2(n590), .ZN(n505) );
  NOR2_X1 U523 ( .A1(n545), .A2(n542), .ZN(n461) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(n461), .Z(n462) );
  NOR2_X1 U525 ( .A1(n486), .A2(n462), .ZN(n465) );
  XOR2_X1 U526 ( .A(n542), .B(KEYINPUT27), .Z(n474) );
  INV_X1 U527 ( .A(n474), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n568) );
  XNOR2_X1 U529 ( .A(n568), .B(KEYINPUT96), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n471), .A2(n295), .ZN(n477) );
  XOR2_X1 U532 ( .A(n486), .B(KEYINPUT28), .Z(n549) );
  INV_X1 U533 ( .A(n549), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n566), .A2(n472), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n554) );
  XOR2_X1 U536 ( .A(KEYINPUT95), .B(n554), .Z(n475) );
  NOR2_X1 U537 ( .A1(n555), .A2(n475), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n504) );
  NOR2_X1 U539 ( .A1(n478), .A2(n504), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n577), .A2(n479), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n539) );
  NAND2_X1 U543 ( .A1(n505), .A2(n539), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT38), .ZN(n520) );
  NOR2_X1 U545 ( .A1(n542), .A2(n520), .ZN(n485) );
  INV_X1 U546 ( .A(n486), .ZN(n487) );
  AND2_X1 U547 ( .A1(n566), .A2(n487), .ZN(n488) );
  AND2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n493) );
  XNOR2_X1 U549 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n491) );
  NOR2_X1 U550 ( .A1(n545), .A2(n494), .ZN(n583) );
  NAND2_X1 U551 ( .A1(n583), .A2(n523), .ZN(n497) );
  XOR2_X1 U552 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(G176GAT), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(G1349GAT) );
  NAND2_X1 U555 ( .A1(n583), .A2(n409), .ZN(n500) );
  XOR2_X1 U556 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n498) );
  INV_X1 U557 ( .A(n409), .ZN(n580) );
  NAND2_X1 U558 ( .A1(n594), .A2(n580), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(KEYINPUT78), .ZN(n502) );
  XNOR2_X1 U560 ( .A(n502), .B(KEYINPUT16), .ZN(n503) );
  NOR2_X1 U561 ( .A1(n504), .A2(n503), .ZN(n524) );
  NAND2_X1 U562 ( .A1(n505), .A2(n524), .ZN(n512) );
  NOR2_X1 U563 ( .A1(n566), .A2(n512), .ZN(n506) );
  XOR2_X1 U564 ( .A(G1GAT), .B(n506), .Z(n507) );
  XNOR2_X1 U565 ( .A(KEYINPUT34), .B(n507), .ZN(G1324GAT) );
  NOR2_X1 U566 ( .A1(n542), .A2(n512), .ZN(n508) );
  XOR2_X1 U567 ( .A(G8GAT), .B(n508), .Z(G1325GAT) );
  NOR2_X1 U568 ( .A1(n545), .A2(n512), .ZN(n510) );
  XNOR2_X1 U569 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U571 ( .A(G15GAT), .B(n511), .ZN(G1326GAT) );
  NOR2_X1 U572 ( .A1(n549), .A2(n512), .ZN(n513) );
  XOR2_X1 U573 ( .A(G22GAT), .B(n513), .Z(G1327GAT) );
  NOR2_X1 U574 ( .A1(n520), .A2(n566), .ZN(n515) );
  XNOR2_X1 U575 ( .A(KEYINPUT101), .B(KEYINPUT39), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U577 ( .A(G29GAT), .B(n516), .Z(G1328GAT) );
  XNOR2_X1 U578 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n518) );
  NOR2_X1 U579 ( .A1(n545), .A2(n520), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G43GAT), .B(n519), .ZN(G1330GAT) );
  NOR2_X1 U582 ( .A1(n549), .A2(n520), .ZN(n521) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(n521), .Z(n522) );
  XNOR2_X1 U584 ( .A(G50GAT), .B(n522), .ZN(G1331GAT) );
  INV_X1 U585 ( .A(n523), .ZN(n573) );
  NOR2_X1 U586 ( .A1(n585), .A2(n573), .ZN(n538) );
  NAND2_X1 U587 ( .A1(n524), .A2(n538), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT108), .ZN(n533) );
  NOR2_X1 U589 ( .A1(n566), .A2(n533), .ZN(n529) );
  XOR2_X1 U590 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n527) );
  XNOR2_X1 U591 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1332GAT) );
  NOR2_X1 U594 ( .A1(n542), .A2(n533), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(n530), .Z(n531) );
  XNOR2_X1 U596 ( .A(G64GAT), .B(n531), .ZN(G1333GAT) );
  NOR2_X1 U597 ( .A1(n545), .A2(n533), .ZN(n532) );
  XOR2_X1 U598 ( .A(G71GAT), .B(n532), .Z(G1334GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n549), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n535) );
  XNOR2_X1 U601 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1335GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n548) );
  NOR2_X1 U605 ( .A1(n566), .A2(n548), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1336GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n548), .ZN(n543) );
  XOR2_X1 U609 ( .A(KEYINPUT114), .B(n543), .Z(n544) );
  XNOR2_X1 U610 ( .A(G92GAT), .B(n544), .ZN(G1337GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n548), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1338GAT) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U615 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U617 ( .A(G106GAT), .B(n552), .Z(G1339GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n554), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n570), .A2(n563), .ZN(n557) );
  XOR2_X1 U621 ( .A(G113GAT), .B(n557), .Z(G1340GAT) );
  NOR2_X1 U622 ( .A1(n573), .A2(n563), .ZN(n559) );
  XNOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(G120GAT), .B(n560), .Z(G1341GAT) );
  NOR2_X1 U626 ( .A1(n577), .A2(n563), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT50), .B(n561), .Z(n562) );
  XNOR2_X1 U628 ( .A(G127GAT), .B(n562), .ZN(G1342GAT) );
  NOR2_X1 U629 ( .A1(n580), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1343GAT) );
  XNOR2_X1 U632 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n572) );
  NOR2_X1 U633 ( .A1(n566), .A2(n553), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT120), .B(n569), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n570), .A2(n579), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1344GAT) );
  NOR2_X1 U638 ( .A1(n579), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G148GAT), .B(n576), .ZN(G1345GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G155GAT), .B(n578), .Z(G1346GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G162GAT), .B(n581), .Z(G1347GAT) );
  NAND2_X1 U646 ( .A1(n583), .A2(n585), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G169GAT), .B(n582), .ZN(G1348GAT) );
  NAND2_X1 U648 ( .A1(n594), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n593), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT61), .Z(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n590), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1353GAT) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(G211GAT), .ZN(G1354GAT) );
endmodule

