//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n223), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n244), .B(new_n250), .Z(G351));
  AOI21_X1  g0051(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(G244), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G274), .A3(new_n255), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OR3_X1    g0062(.A1(new_n257), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n269), .A2(G238), .B1(new_n272), .B2(G107), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1698), .B1(new_n267), .B2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n223), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n252), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT67), .B1(new_n257), .B2(new_n262), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n263), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G200), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT68), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G190), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n218), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n286), .A2(new_n288), .B1(new_n209), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT15), .B(G87), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n209), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n285), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n285), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n208), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G77), .A3(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n294), .B(new_n299), .C1(G77), .C2(new_n295), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n263), .A2(new_n277), .A3(new_n278), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n303), .B2(KEYINPUT68), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n283), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n279), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n300), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n285), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n204), .A2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n286), .ZN(new_n315));
  INV_X1    g0115(.A(new_n292), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n315), .A2(new_n316), .B1(G150), .B2(new_n287), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n297), .A2(G50), .A3(new_n298), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G50), .B2(new_n295), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n269), .A2(G223), .B1(new_n272), .B2(G77), .ZN(new_n322));
  INV_X1    g0122(.A(G222), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n275), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n252), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n262), .B1(G226), .B2(new_n256), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(G179), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n321), .B(new_n328), .C1(new_n308), .C2(new_n327), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n318), .A2(new_n320), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT9), .ZN(new_n331));
  INV_X1    g0131(.A(new_n327), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n331), .B1(G190), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n321), .A2(KEYINPUT9), .B1(G200), .B2(new_n327), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n329), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n312), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n316), .A2(G77), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n313), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT11), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n297), .A2(G68), .A3(new_n298), .ZN(new_n345));
  INV_X1    g0145(.A(G13), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(G1), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(G20), .A3(new_n246), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT12), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n349), .A2(KEYINPUT12), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n345), .B(new_n352), .C1(new_n350), .C2(new_n348), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  OAI211_X1 g0157(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT69), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n267), .A2(new_n268), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n361), .A2(KEYINPUT69), .A3(G232), .A4(G1698), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n274), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n252), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT70), .ZN(new_n367));
  INV_X1    g0167(.A(G274), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n258), .B2(new_n259), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n369), .B2(new_n255), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n367), .A3(new_n255), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n371), .A2(new_n372), .B1(G238), .B2(new_n256), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n357), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n260), .B1(new_n363), .B2(new_n364), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n256), .A2(G238), .ZN(new_n376));
  INV_X1    g0176(.A(new_n372), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n370), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n375), .A2(new_n378), .A3(KEYINPUT13), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n356), .B(G169), .C1(new_n374), .C2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n366), .A2(new_n357), .A3(new_n373), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT13), .B1(new_n375), .B2(new_n378), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G179), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n382), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n356), .B1(new_n385), .B2(G169), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n355), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(G200), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n354), .C1(new_n302), .C2(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n267), .A2(new_n209), .A3(new_n268), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n246), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n222), .A2(new_n246), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n287), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n391), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n272), .B2(new_n209), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n270), .A2(new_n271), .A3(new_n393), .A4(G20), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n400), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n406), .A3(new_n285), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n286), .B1(new_n208), .B2(G20), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n297), .B1(new_n296), .B2(new_n286), .ZN(new_n409));
  INV_X1    g0209(.A(G226), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G1698), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n411), .B1(G223), .B2(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n252), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n256), .A2(G232), .B1(new_n255), .B2(new_n369), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n302), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n260), .B1(new_n412), .B2(new_n413), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n260), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n261), .B1(new_n420), .B2(new_n223), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n280), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n407), .A2(new_n409), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT72), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n407), .A2(new_n426), .A3(new_n423), .A4(new_n409), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n429));
  NAND4_X1  g0229(.A1(new_n407), .A2(new_n409), .A3(new_n423), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n407), .A2(new_n409), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  AOI21_X1  g0233(.A(G169), .B1(new_n415), .B2(new_n416), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n418), .A2(new_n421), .A3(G179), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n432), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n340), .A2(new_n390), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n296), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n208), .A2(G33), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n295), .A2(new_n444), .A3(new_n218), .A4(new_n284), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n445), .B2(new_n442), .ZN(new_n446));
  AOI21_X1  g0246(.A(G20), .B1(G33), .B2(G283), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G33), .B2(new_n224), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(G20), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n285), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(KEYINPUT20), .A3(new_n285), .A4(new_n449), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n361), .A2(KEYINPUT77), .A3(G264), .A4(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n272), .A2(G303), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n361), .A2(G257), .A3(new_n264), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n252), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n254), .A2(G1), .ZN(new_n464));
  AND2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(G270), .A3(new_n260), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n208), .A2(G45), .ZN(new_n469));
  OR2_X1    g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n369), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n306), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n462), .B2(new_n252), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n478), .A2(new_n479), .A3(new_n308), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n455), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n455), .B1(new_n476), .B2(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n302), .B2(new_n476), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT79), .B(KEYINPUT21), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n478), .A2(new_n308), .A3(new_n454), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR4_X1   g0287(.A1(new_n478), .A2(new_n454), .A3(KEYINPUT78), .A4(new_n308), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n481), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n491), .A2(new_n224), .A3(G107), .ZN(new_n492));
  XNOR2_X1  g0292(.A(G97), .B(G107), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n494), .A2(new_n209), .B1(new_n289), .B2(new_n288), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n394), .B2(new_n395), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n285), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n296), .A2(new_n224), .ZN(new_n499));
  INV_X1    g0299(.A(new_n445), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G97), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n472), .A2(new_n225), .A3(new_n252), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n269), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT74), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(new_n264), .C1(new_n270), .C2(new_n271), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT4), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n274), .A2(KEYINPUT74), .A3(KEYINPUT4), .A4(G244), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n504), .B1(new_n512), .B2(new_n252), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G190), .A3(new_n473), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n252), .ZN(new_n515));
  INV_X1    g0315(.A(new_n504), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(new_n473), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n503), .B(new_n514), .C1(new_n517), .C2(new_n280), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n306), .A3(new_n473), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n502), .C1(new_n517), .C2(G169), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n496), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT25), .B1(new_n296), .B2(new_n496), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(new_n496), .B2(new_n445), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n467), .A2(G264), .A3(new_n260), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(new_n473), .ZN(new_n528));
  OAI211_X1 g0328(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(new_n264), .C1(new_n270), .C2(new_n271), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n252), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n280), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G190), .B2(new_n534), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT80), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n496), .A3(G20), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n496), .A2(G20), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT80), .B1(new_n543), .B2(KEYINPUT23), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT22), .ZN(new_n546));
  AOI21_X1  g0346(.A(G20), .B1(new_n267), .B2(new_n268), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(G87), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n209), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(KEYINPUT22), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT24), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n361), .A2(new_n546), .A3(new_n209), .A4(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n545), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n537), .B1(new_n558), .B2(new_n285), .ZN(new_n559));
  AOI211_X1 g0359(.A(KEYINPUT81), .B(new_n313), .C1(new_n552), .C2(new_n557), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n526), .B(new_n536), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n555), .A2(new_n556), .A3(new_n545), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n556), .B1(new_n555), .B2(new_n545), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n285), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT81), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n537), .A3(new_n285), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n525), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n534), .A2(KEYINPUT82), .A3(new_n306), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n528), .A2(G179), .A3(new_n533), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n527), .A2(new_n473), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n252), .B2(new_n532), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(new_n308), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n568), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n561), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n209), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT75), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT75), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n580), .A3(new_n209), .ZN(new_n581));
  INV_X1    g0381(.A(G87), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n224), .A3(new_n496), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n292), .B2(new_n224), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT76), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n585), .C1(new_n292), .C2(new_n224), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n547), .A2(G68), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n584), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(new_n285), .B1(new_n296), .B2(new_n291), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n445), .A2(new_n291), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n369), .A2(new_n464), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n260), .A2(G250), .A3(new_n469), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G238), .B(new_n264), .C1(new_n270), .C2(new_n271), .ZN(new_n599));
  OAI211_X1 g0399(.A(G244), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G116), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n252), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G179), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n252), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n596), .A2(new_n597), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n500), .A2(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n592), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n603), .A2(G190), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(G200), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n595), .A2(new_n609), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n576), .A2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n441), .A2(new_n490), .A3(new_n521), .A4(new_n616), .ZN(G372));
  AND3_X1   g0417(.A1(new_n604), .A2(new_n608), .A3(KEYINPUT83), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT83), .B1(new_n604), .B2(new_n608), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n618), .A2(new_n619), .B1(new_n594), .B2(new_n593), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n567), .A2(new_n575), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n592), .A2(KEYINPUT84), .A3(new_n610), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT84), .B1(new_n592), .B2(new_n610), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n613), .B(new_n612), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n561), .A2(new_n520), .A3(new_n626), .A4(new_n518), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n620), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n615), .B2(new_n520), .ZN(new_n629));
  INV_X1    g0429(.A(new_n520), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n620), .A3(new_n626), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n631), .B2(KEYINPUT26), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n441), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n336), .A2(new_n338), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n311), .A2(new_n389), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n635), .A2(new_n387), .B1(new_n428), .B2(new_n430), .ZN(new_n636));
  INV_X1    g0436(.A(new_n439), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n329), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT85), .Z(G369));
  NAND2_X1  g0442(.A1(new_n347), .A2(new_n209), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G213), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(KEYINPUT27), .B2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n454), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n489), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n622), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT86), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT86), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n653), .A3(new_n650), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n526), .B1(new_n559), .B2(new_n560), .ZN(new_n658));
  INV_X1    g0458(.A(new_n575), .ZN(new_n659));
  INV_X1    g0459(.A(new_n647), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n567), .A2(new_n647), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n576), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT87), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n661), .C1(new_n576), .C2(new_n662), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n658), .A2(new_n659), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n660), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n622), .A2(new_n647), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n670), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(KEYINPUT88), .ZN(new_n675));
  INV_X1    g0475(.A(new_n212), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(G41), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n212), .A2(KEYINPUT88), .A3(new_n253), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n583), .A2(G116), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n680), .A2(new_n208), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n217), .B2(new_n680), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT28), .Z(new_n685));
  NAND4_X1  g0485(.A1(new_n616), .A2(new_n490), .A3(new_n521), .A4(new_n647), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n478), .A2(new_n573), .A3(G179), .A4(new_n603), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n515), .A2(new_n516), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n513), .A2(new_n473), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n534), .A2(new_n306), .A3(new_n607), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n476), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n463), .A2(new_n603), .A3(new_n475), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(KEYINPUT30), .A3(new_n513), .A4(new_n569), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n660), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n686), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n647), .B1(new_n628), .B2(new_n632), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n630), .A2(KEYINPUT26), .A3(new_n620), .A4(new_n626), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT26), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n615), .B2(new_n520), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT29), .B(new_n647), .C1(new_n628), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n701), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n685), .B1(new_n710), .B2(G1), .ZN(G364));
  INV_X1    g0511(.A(new_n655), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n346), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n208), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n680), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n656), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n258), .B1(new_n209), .B2(G169), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT91), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n302), .A2(new_n280), .ZN(new_n726));
  NAND2_X1  g0526(.A1(G20), .A2(G179), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT95), .Z(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n302), .A3(new_n280), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n730), .A2(G326), .B1(G311), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G294), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(G190), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n209), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n733), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n280), .A2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n209), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n272), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n727), .A2(new_n302), .A3(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G322), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n726), .A2(new_n742), .ZN(new_n748));
  INV_X1    g0548(.A(G303), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n727), .A2(new_n280), .A3(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT33), .B(G317), .Z(new_n752));
  OAI221_X1 g0552(.A(new_n747), .B1(new_n748), .B2(new_n749), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n209), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n736), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n745), .B(new_n753), .C1(G329), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n740), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n748), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G87), .ZN(new_n760));
  INV_X1    g0560(.A(new_n746), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n760), .B1(new_n222), .B2(new_n761), .C1(new_n289), .C2(new_n731), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n361), .B1(new_n751), .B2(new_n246), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n729), .A2(new_n202), .B1(new_n743), .B2(new_n496), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n738), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n765), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n725), .B1(new_n758), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT90), .Z(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n725), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT92), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n676), .A2(new_n272), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G355), .B1(new_n442), .B2(new_n676), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n676), .A2(new_n361), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT89), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G45), .B2(new_n216), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n250), .A2(new_n254), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n719), .B(new_n773), .C1(new_n780), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n655), .B2(new_n777), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n720), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n311), .A2(new_n647), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n660), .A2(new_n300), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n283), .B2(new_n304), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n792), .B1(new_n795), .B2(new_n311), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n702), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n796), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n798), .B(new_n647), .C1(new_n628), .C2(new_n632), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n718), .B1(new_n800), .B2(new_n700), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n701), .A2(new_n797), .A3(new_n799), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n724), .A2(new_n774), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n718), .B1(G77), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n798), .A2(new_n775), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n756), .A2(G311), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n751), .A2(new_n744), .B1(new_n743), .B2(new_n582), .ZN(new_n809));
  INV_X1    g0609(.A(new_n729), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G303), .B2(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n761), .A2(new_n734), .B1(new_n731), .B2(new_n442), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n361), .B(new_n812), .C1(G107), .C2(new_n759), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n771), .A2(new_n808), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n810), .A2(G137), .B1(G150), .B2(new_n750), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT97), .B(G143), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n766), .B2(new_n731), .C1(new_n761), .C2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT34), .Z(new_n818));
  NOR2_X1   g0618(.A1(new_n743), .A2(new_n246), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n272), .B(new_n819), .C1(G50), .C2(new_n759), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n755), .C1(new_n222), .C2(new_n738), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n814), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n806), .B(new_n807), .C1(new_n724), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n803), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  INV_X1    g0626(.A(new_n494), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT35), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT35), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n828), .A2(G116), .A3(new_n219), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT36), .Z(new_n831));
  OR3_X1    g0631(.A1(new_n216), .A2(new_n289), .A3(new_n397), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n208), .B(G13), .C1(new_n832), .C2(new_n245), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT98), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n354), .A2(new_n647), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AND4_X1   g0637(.A1(new_n835), .A2(new_n387), .A3(new_n389), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n387), .A2(new_n389), .A3(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n384), .A2(new_n386), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n389), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n835), .B1(new_n841), .B2(new_n836), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n838), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT103), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n513), .A2(new_n569), .A3(new_n478), .A4(new_n603), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n607), .A2(new_n306), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n847), .A2(new_n478), .A3(new_n573), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n687), .A2(new_n846), .B1(new_n848), .B2(new_n691), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n647), .B1(new_n849), .B2(new_n695), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT102), .B1(new_n850), .B2(KEYINPUT31), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT31), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n697), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n686), .A2(new_n845), .A3(new_n855), .ZN(new_n856));
  AND4_X1   g0656(.A1(KEYINPUT40), .A2(new_n843), .A3(new_n856), .A4(new_n798), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n401), .A2(new_n406), .A3(new_n285), .ZN(new_n859));
  INV_X1    g0659(.A(new_n409), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n859), .A2(new_n860), .B1(new_n436), .B2(new_n646), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n424), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n425), .A2(new_n861), .A3(new_n864), .A4(new_n427), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT99), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT100), .B(new_n863), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n432), .A2(new_n646), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n440), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n425), .A2(new_n427), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n874), .A2(KEYINPUT99), .A3(new_n864), .A4(new_n861), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n865), .A2(new_n866), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT100), .B1(new_n877), .B2(new_n863), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n858), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n425), .A2(new_n861), .A3(new_n427), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n867), .B2(new_n868), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n857), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n843), .A2(new_n856), .A3(new_n798), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n875), .A2(new_n876), .B1(KEYINPUT37), .B2(new_n880), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n870), .B1(new_n431), .B2(new_n439), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n888), .A2(new_n858), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n882), .B2(new_n872), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n886), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT104), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n441), .A2(new_n856), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(G330), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n799), .A2(new_n792), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n843), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n901), .A2(new_n892), .B1(new_n439), .B2(new_n646), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT101), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n883), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT100), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n872), .A3(new_n869), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n858), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n858), .B1(new_n888), .B2(new_n889), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n904), .B1(new_n911), .B2(new_n883), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n903), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n889), .B1(new_n877), .B2(new_n881), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT39), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n879), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n883), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT39), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT101), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n387), .A2(new_n660), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n902), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n704), .A2(new_n441), .A3(new_n709), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n924), .A2(new_n640), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n899), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n208), .B2(new_n715), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n899), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n834), .B1(new_n928), .B2(new_n929), .ZN(G367));
  INV_X1    g0730(.A(new_n784), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n780), .B1(new_n212), .B2(new_n291), .C1(new_n236), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n718), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT107), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n624), .A2(new_n625), .A3(new_n647), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(new_n620), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n620), .A3(new_n626), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n743), .A2(new_n289), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G50), .B2(new_n732), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n272), .B1(new_n759), .B2(G58), .ZN(new_n941));
  AOI22_X1  g0741(.A1(G150), .A2(new_n746), .B1(new_n750), .B2(G159), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n816), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n730), .A2(new_n944), .B1(G137), .B2(new_n756), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n943), .B(new_n946), .C1(G68), .C2(new_n770), .ZN(new_n947));
  INV_X1    g0747(.A(new_n743), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(G97), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n749), .B2(new_n761), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G294), .B2(new_n750), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT46), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n748), .A2(new_n952), .A3(new_n442), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n361), .B(new_n953), .C1(G283), .C2(new_n732), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n951), .B(new_n954), .C1(new_n496), .C2(new_n738), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n730), .A2(G311), .B1(G317), .B2(new_n756), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n952), .B1(new_n748), .B2(new_n442), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT108), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n947), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(KEYINPUT47), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT47), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n724), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n934), .B1(new_n777), .B2(new_n938), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT109), .Z(new_n966));
  INV_X1    g0766(.A(new_n666), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n658), .A2(new_n660), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n669), .A2(new_n968), .A3(new_n561), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n665), .B1(new_n969), .B2(new_n661), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n672), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n670), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n521), .B1(new_n503), .B2(new_n647), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n630), .A2(new_n660), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n979), .B(new_n976), .C1(new_n971), .C2(new_n972), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT45), .B1(new_n673), .B2(new_n976), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n671), .B1(new_n664), .B2(new_n666), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n982), .A2(new_n983), .A3(new_n670), .A4(new_n977), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n978), .A2(new_n980), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n668), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n983), .B1(new_n973), .B2(new_n977), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n979), .B1(new_n673), .B2(new_n976), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n973), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n993), .A3(new_n668), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n667), .A2(new_n672), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n982), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n657), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n656), .B1(new_n982), .B2(new_n995), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n710), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n987), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n710), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n679), .B(KEYINPUT41), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n717), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n520), .B1(new_n974), .B2(new_n669), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n647), .ZN(new_n1006));
  XOR2_X1   g0806(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n1007));
  AND3_X1   g0807(.A1(new_n936), .A2(new_n937), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT106), .B1(new_n971), .B2(new_n977), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT106), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n982), .A2(new_n1010), .A3(new_n976), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1011), .A3(KEYINPUT42), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT42), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1006), .B(new_n1008), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1014), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1016), .A2(new_n1012), .B1(new_n647), .B2(new_n1005), .ZN(new_n1017));
  MUX2_X1   g0817(.A(new_n1007), .B(KEYINPUT43), .S(new_n938), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n668), .A2(new_n977), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1015), .B(new_n1020), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n966), .B1(new_n1004), .B2(new_n1024), .ZN(G387));
  NOR2_X1   g0825(.A1(new_n999), .A2(new_n679), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n997), .A2(new_n998), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n710), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n781), .A2(new_n682), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(G107), .B2(new_n212), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n286), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI211_X1 g0832(.A(G45), .B(new_n682), .C1(G68), .C2(G77), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n931), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n240), .A2(new_n254), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n718), .B1(new_n1036), .B2(new_n779), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n667), .A2(new_n777), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n738), .A2(new_n291), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n202), .B2(new_n761), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT110), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n748), .A2(new_n289), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G159), .B2(new_n810), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n361), .A3(new_n949), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G150), .B2(new_n756), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n751), .A2(new_n286), .B1(new_n731), .B2(new_n246), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT111), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n756), .A2(G326), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n361), .B1(new_n948), .B2(G116), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n732), .A2(G303), .B1(G311), .B2(new_n750), .ZN(new_n1051));
  INV_X1    g0851(.A(G317), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n761), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT112), .B(G322), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n730), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n770), .A2(G283), .B1(G294), .B2(new_n759), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT113), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1049), .B(new_n1050), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1048), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1037), .B(new_n1038), .C1(new_n724), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1027), .B2(new_n717), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1028), .A2(new_n1066), .ZN(G393));
  INV_X1    g0867(.A(new_n999), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n990), .A2(new_n993), .A3(new_n668), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n668), .B1(new_n990), .B2(new_n993), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n680), .A3(new_n1000), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n784), .A2(new_n244), .B1(G97), .B2(new_n676), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n780), .A2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n718), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n976), .A2(new_n777), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n361), .B1(new_n743), .B2(new_n582), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G68), .A2(new_n759), .B1(new_n732), .B2(new_n315), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n202), .B2(new_n751), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(new_n756), .C2(new_n944), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n810), .A2(G150), .B1(G159), .B2(new_n746), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G77), .B2(new_n770), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n272), .B1(new_n743), .B2(new_n496), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G283), .A2(new_n759), .B1(new_n732), .B2(G294), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n749), .B2(new_n751), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n756), .C2(new_n1054), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n810), .A2(G317), .B1(G311), .B2(new_n746), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G116), .B2(new_n770), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1082), .A2(new_n1085), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1093), .A2(KEYINPUT115), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n725), .B1(new_n1093), .B2(KEYINPUT115), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1077), .B(new_n1078), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n717), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1072), .A2(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n901), .A2(new_n921), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n913), .A2(new_n919), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n713), .B(new_n796), .C1(new_n686), .C2(new_n698), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n843), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n843), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n310), .B1(new_n305), .B2(new_n794), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n647), .B(new_n1105), .C1(new_n628), .C2(new_n708), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n792), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n884), .B(new_n921), .C1(new_n1104), .C2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1101), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n843), .A2(new_n856), .A3(G330), .A4(new_n798), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n441), .A2(G330), .A3(new_n856), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n924), .A2(new_n1114), .A3(new_n640), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n856), .A2(G330), .A3(new_n798), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1104), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1107), .B1(new_n1102), .B2(new_n843), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(KEYINPUT116), .A3(new_n1118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1104), .B1(new_n700), .B2(new_n796), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1125), .A2(new_n1111), .B1(new_n792), .B2(new_n799), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1116), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n679), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1101), .A2(new_n1109), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1111), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1101), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1122), .A2(KEYINPUT116), .A3(new_n1118), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT116), .B1(new_n1122), .B2(new_n1118), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1127), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1115), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT117), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(KEYINPUT117), .B(new_n1138), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1129), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n920), .A2(new_n775), .ZN(new_n1143));
  INV_X1    g0943(.A(G150), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n748), .A2(KEYINPUT53), .A3(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n272), .B1(new_n732), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT53), .B1(new_n748), .B2(new_n1144), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n810), .A2(G128), .B1(G137), .B2(new_n750), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n202), .B2(new_n743), .C1(new_n821), .C2(new_n761), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(G125), .C2(new_n756), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n770), .A2(G159), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n732), .A2(G97), .B1(G107), .B2(new_n750), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n744), .B2(new_n729), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n819), .B1(G116), .B2(new_n746), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n272), .A3(new_n760), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G294), .C2(new_n756), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n770), .A2(G77), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1153), .A2(new_n1154), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n718), .B1(new_n315), .B2(new_n805), .C1(new_n1161), .C2(new_n725), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1143), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1113), .B2(new_n717), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1142), .A2(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(KEYINPUT119), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n916), .A2(KEYINPUT101), .A3(new_n918), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT101), .B1(new_n916), .B2(new_n918), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n922), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n902), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1166), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n885), .A2(G330), .A3(new_n893), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n330), .A2(new_n646), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT118), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n339), .B(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1177));
  AND2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1172), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n885), .A2(new_n1180), .A3(new_n893), .A4(G330), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1171), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1171), .A2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n717), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1180), .A2(new_n775), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n948), .A2(G58), .B1(new_n746), .B2(G107), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n291), .B2(new_n731), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n272), .A2(new_n253), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n751), .A2(new_n224), .B1(new_n729), .B2(new_n442), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1190), .A2(new_n1042), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n246), .B2(new_n738), .C1(new_n744), .C2(new_n755), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G50), .B1(new_n266), .B2(new_n253), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1194), .A2(new_n1195), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n759), .A2(new_n1147), .B1(G128), .B2(new_n746), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n810), .A2(G125), .B1(G132), .B2(new_n750), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n732), .A2(G137), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n770), .B2(G150), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n266), .B(new_n253), .C1(new_n743), .C2(new_n766), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n756), .B2(G124), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT59), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1197), .B1(new_n1195), .B2(new_n1194), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n724), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n718), .C1(G50), .C2(new_n805), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1188), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT120), .B1(new_n1187), .B2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1183), .B(new_n1182), .C1(new_n923), .C2(new_n1166), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1171), .A2(new_n1184), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n716), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1212), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1116), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1184), .A2(new_n923), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n921), .B1(new_n913), .B2(new_n919), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1182), .B(new_n1183), .C1(new_n1222), .C2(new_n902), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(KEYINPUT57), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n680), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1132), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1115), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1214), .A2(new_n1219), .B1(new_n1225), .B2(new_n1229), .ZN(G375));
  AOI22_X1  g1030(.A1(new_n732), .A2(G107), .B1(G283), .B2(new_n746), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n734), .B2(new_n729), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n939), .A2(new_n361), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n224), .B2(new_n748), .C1(new_n442), .C2(new_n751), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G303), .C2(new_n756), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n746), .A2(G137), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1144), .B2(new_n731), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n810), .A2(G132), .B1(new_n1147), .B2(new_n750), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n766), .B2(new_n748), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(G128), .C2(new_n756), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n361), .B1(new_n743), .B2(new_n222), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT121), .Z(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G50), .B2(new_n770), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1235), .A2(new_n1039), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n718), .B1(G68), .B2(new_n805), .C1(new_n1244), .C2(new_n725), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1104), .B2(new_n774), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1137), .B2(new_n717), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1138), .A2(new_n1003), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1126), .B(new_n1115), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(G381));
  AND2_X1   g1050(.A1(new_n1142), .A2(new_n1164), .ZN(new_n1251));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n825), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1254), .A2(G387), .A3(G381), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1221), .A2(KEYINPUT57), .A3(new_n1223), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1227), .A2(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1226), .A2(new_n1115), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n680), .C1(KEYINPUT57), .C2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1187), .A2(KEYINPUT120), .A3(new_n1213), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1218), .B1(new_n1217), .B2(new_n1212), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1251), .A2(new_n1255), .A3(new_n1259), .A4(new_n1262), .ZN(G407));
  INV_X1    g1063(.A(G343), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(G213), .ZN(new_n1265));
  OR2_X1    g1065(.A1(G378), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(G409));
  NAND2_X1  g1067(.A1(new_n1258), .A2(new_n1003), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1221), .A2(new_n717), .A3(new_n1223), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1213), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1251), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G378), .A2(new_n1262), .A3(new_n1259), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1249), .B1(new_n1138), .B2(KEYINPUT60), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1127), .A4(new_n1116), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n680), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1247), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n825), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G384), .B(new_n1247), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT122), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1273), .A2(new_n1265), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT124), .B1(G387), .B2(new_n1252), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n790), .B1(new_n1028), .B2(new_n1066), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1253), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G390), .B(new_n966), .C1(new_n1004), .C2(new_n1024), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1002), .B1(new_n1000), .B2(new_n710), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1022), .B(new_n1023), .C1(new_n1292), .C2(new_n717), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G390), .B1(new_n1293), .B2(new_n966), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n1286), .A2(new_n1289), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1252), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(new_n1288), .A3(KEYINPUT124), .A4(new_n1290), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1285), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1273), .A2(new_n1265), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1281), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1264), .A2(G213), .A3(G2897), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1279), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT123), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1282), .A2(new_n1307), .A3(new_n1303), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1303), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1301), .A2(new_n1306), .A3(new_n1308), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1299), .A2(new_n1300), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1283), .A2(KEYINPUT62), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1273), .A2(new_n1316), .A3(new_n1265), .A4(new_n1282), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1312), .A2(new_n1315), .A3(new_n1300), .A4(new_n1317), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1295), .A2(KEYINPUT125), .A3(new_n1297), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT125), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1318), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1314), .A2(new_n1323), .ZN(G405));
  AND3_X1   g1124(.A1(new_n1262), .A2(G378), .A3(new_n1259), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G378), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1282), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G375), .A2(new_n1251), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n1272), .A3(new_n1309), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(KEYINPUT126), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1331), .B(new_n1282), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1330), .A2(new_n1321), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1322), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1330), .A2(new_n1321), .A3(KEYINPUT127), .A4(new_n1332), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1335), .A2(new_n1337), .A3(new_n1338), .ZN(G402));
endmodule


