//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT94), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT67), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT2), .A3(G113), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n193), .A2(new_n195), .B1(new_n191), .B2(new_n192), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G116), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT68), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n196), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G107), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT82), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n203), .B(G104), .C1(new_n205), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(G104), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(KEYINPUT3), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT83), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT83), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n216), .A3(new_n211), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(G101), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n208), .A2(new_n216), .A3(new_n211), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n208), .B2(new_n211), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n208), .A2(new_n221), .A3(new_n211), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n214), .A3(KEYINPUT4), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n202), .B(new_n218), .C1(new_n222), .C2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G116), .B(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT5), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n192), .B1(new_n198), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT88), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n206), .A2(KEYINPUT82), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n204), .A2(G107), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n210), .B1(new_n235), .B2(G104), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n237), .A2(new_n223), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n196), .A2(new_n226), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n225), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(G110), .B(G122), .Z(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT90), .B(KEYINPUT6), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n242), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n246), .A3(new_n240), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT89), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT89), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n243), .A2(new_n250), .A3(KEYINPUT6), .A4(new_n247), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n245), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G143), .B(G146), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n255), .A3(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OR3_X1    g078(.A1(new_n264), .A2(KEYINPUT91), .A3(G125), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT91), .B1(new_n264), .B2(G125), .ZN(new_n266));
  INV_X1    g080(.A(G125), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(KEYINPUT0), .A3(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n257), .A2(KEYINPUT0), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT0), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n260), .A2(new_n275), .A3(KEYINPUT64), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(G224), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n252), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(KEYINPUT7), .B2(new_n280), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n242), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n227), .B(KEYINPUT93), .ZN(new_n288));
  INV_X1    g102(.A(new_n229), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n239), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n238), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n238), .B1(new_n232), .B2(new_n239), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n283), .A2(new_n285), .A3(new_n247), .A4(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n190), .B1(new_n282), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n245), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n225), .A2(new_n246), .A3(new_n240), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n246), .B1(new_n225), .B2(new_n240), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n250), .B1(new_n301), .B2(KEYINPUT6), .ZN(new_n302));
  INV_X1    g116(.A(new_n251), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n281), .B(new_n298), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AND4_X1   g118(.A1(new_n297), .A2(new_n304), .A3(new_n190), .A4(new_n295), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n187), .B1(new_n296), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT95), .ZN(new_n307));
  INV_X1    g121(.A(new_n187), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n297), .A3(new_n295), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n189), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(new_n297), .A3(new_n190), .A4(new_n295), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT95), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G472), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT65), .B(G131), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G137), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n319), .B2(G137), .ZN(new_n322));
  INV_X1    g136(.A(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n320), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n320), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n319), .A2(G137), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n264), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n320), .A3(new_n324), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT66), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT66), .A4(new_n320), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G131), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n325), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(new_n277), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n335), .B2(new_n277), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT30), .B(new_n329), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n277), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n329), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT30), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n325), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n333), .A2(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n330), .A2(new_n331), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT69), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n335), .A2(new_n336), .A3(new_n277), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT30), .A4(new_n329), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n340), .A2(new_n202), .A3(new_n344), .A4(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G237), .A2(G953), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G210), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(new_n221), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n202), .B(KEYINPUT71), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n352), .A2(new_n361), .A3(new_n329), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n365));
  INV_X1    g179(.A(new_n361), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(new_n342), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n352), .A2(new_n361), .A3(KEYINPUT28), .A4(new_n329), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n342), .A2(new_n202), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n367), .A2(new_n317), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n360), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n317), .B1(new_n364), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n329), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n366), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n365), .B1(new_n375), .B2(new_n362), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n367), .A2(KEYINPUT73), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n378));
  INV_X1    g192(.A(new_n342), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n361), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n380), .B2(new_n365), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n376), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n382), .B2(new_n372), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n316), .B1(new_n373), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n371), .A2(KEYINPUT72), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n355), .A2(new_n362), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT31), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n355), .A2(KEYINPUT31), .A3(new_n362), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n367), .A2(new_n369), .A3(new_n368), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n360), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n394));
  NOR2_X1   g208(.A1(G472), .A2(G902), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n388), .A2(new_n389), .B1(new_n360), .B2(new_n391), .ZN(new_n397));
  INV_X1    g211(.A(new_n395), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT32), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n384), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n257), .A2(G119), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n199), .A2(G128), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G110), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n402), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT75), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n402), .A3(KEYINPUT75), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT24), .B(G110), .Z(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G140), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(KEYINPUT76), .B2(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT76), .A2(G125), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(G140), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT16), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT16), .B1(new_n415), .B2(G125), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n258), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT16), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(G140), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(KEYINPUT76), .A3(G125), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n426), .A2(G146), .A3(new_n420), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n408), .B(new_n414), .C1(new_n422), .C2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(G125), .B(G140), .Z(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(G146), .ZN(new_n430));
  OAI21_X1  g244(.A(G146), .B1(new_n426), .B2(new_n420), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n413), .B1(new_n411), .B2(new_n412), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n407), .A2(G110), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n401), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT22), .B(G137), .Z(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n434), .A3(new_n401), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G217), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(G234), .B2(new_n297), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G902), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n441), .A2(new_n442), .ZN(new_n450));
  INV_X1    g264(.A(new_n442), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(new_n435), .A3(new_n440), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n297), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT80), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT25), .B1(new_n443), .B2(new_n297), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n449), .B(new_n456), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n448), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n277), .B(new_n218), .C1(new_n222), .C2(new_n224), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n263), .A2(KEYINPUT85), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n263), .A2(KEYINPUT85), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n261), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n238), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT10), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n238), .A2(KEYINPUT10), .A3(new_n264), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n335), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n463), .A2(new_n469), .A3(new_n348), .A4(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n279), .A2(G227), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(G140), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT81), .B(G110), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n264), .B1(new_n223), .B2(new_n237), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n238), .B2(new_n466), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT12), .B1(new_n482), .B2(new_n348), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n484));
  INV_X1    g298(.A(new_n467), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n484), .B(new_n335), .C1(new_n485), .C2(new_n481), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n473), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n473), .A3(new_n486), .A4(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n480), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G469), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n473), .A2(new_n486), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n478), .A4(new_n483), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT87), .B1(new_n487), .B2(new_n479), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n474), .A2(new_n479), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n297), .ZN(new_n501));
  NAND2_X1  g315(.A1(G469), .A2(G902), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT9), .B(G234), .ZN(new_n504));
  OAI21_X1  g318(.A(G221), .B1(new_n504), .B2(G902), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n400), .A2(new_n462), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n318), .ZN(new_n508));
  INV_X1    g322(.A(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n279), .A3(G214), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(new_n253), .ZN(new_n511));
  AOI21_X1  g325(.A(G143), .B1(new_n356), .B2(G214), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n508), .B(KEYINPUT98), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n253), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n356), .A2(G143), .A3(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT98), .B1(new_n517), .B2(new_n508), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT17), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT98), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n515), .A2(new_n516), .A3(new_n318), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n513), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n422), .A2(new_n427), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(G113), .B(G122), .Z(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(G104), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT100), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT18), .A2(G131), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n517), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n416), .B2(new_n418), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT96), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n258), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n430), .A2(KEYINPUT97), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n532), .B(new_n538), .C1(new_n536), .C2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n527), .A2(new_n530), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n529), .B1(new_n527), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n297), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT101), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT101), .B(new_n297), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(G475), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G475), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n535), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT19), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n429), .A2(KEYINPUT19), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n549), .B2(KEYINPUT19), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n258), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n514), .A2(new_n518), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n422), .B1(new_n556), .B2(new_n524), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n529), .B1(new_n558), .B2(new_n540), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n548), .B(new_n297), .C1(new_n559), .C2(new_n541), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n527), .A2(new_n530), .A3(new_n540), .ZN(new_n563));
  INV_X1    g377(.A(new_n540), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n555), .B2(new_n557), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n565), .B2(new_n529), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n566), .A2(KEYINPUT20), .A3(new_n548), .A4(new_n297), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n547), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G128), .B(G143), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT13), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n257), .A2(KEYINPUT13), .A3(G143), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(G134), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n319), .ZN(new_n573));
  XNOR2_X1  g387(.A(G116), .B(G122), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n235), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n235), .A2(new_n574), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n572), .B(new_n573), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n569), .B(new_n319), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT14), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n197), .A2(KEYINPUT14), .A3(G122), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(G107), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n583), .A3(new_n576), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n504), .A2(new_n444), .A3(G953), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n297), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n279), .A2(G952), .ZN(new_n594));
  INV_X1    g408(.A(G234), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n509), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n297), .B(new_n279), .C1(G234), .C2(G237), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT21), .B(G898), .Z(new_n599));
  OAI21_X1  g413(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT102), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n568), .A2(new_n593), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n315), .A2(new_n507), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT103), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G3));
  INV_X1    g420(.A(new_n568), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n588), .A2(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n587), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(G478), .B(new_n297), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT104), .B(G478), .Z(new_n613));
  AND3_X1   g427(.A1(new_n589), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n589), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n312), .A2(new_n601), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n459), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n447), .B1(new_n621), .B2(new_n460), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n397), .B2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n397), .A2(new_n398), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n624), .A2(new_n625), .A3(new_n506), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NOR2_X1   g443(.A1(new_n306), .A2(new_n602), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n568), .A2(new_n592), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n428), .A2(new_n434), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n446), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n459), .B2(new_n461), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n623), .B1(new_n397), .B2(new_n398), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n506), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n315), .A2(new_n603), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  NAND2_X1  g458(.A1(new_n373), .A2(new_n383), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n397), .A2(KEYINPUT32), .A3(new_n398), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n503), .A2(new_n639), .A3(new_n505), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n598), .A2(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n596), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n649), .A2(new_n650), .A3(new_n312), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  AND2_X1   g469(.A1(new_n503), .A2(new_n505), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n652), .B(KEYINPUT39), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT40), .Z(new_n659));
  NAND3_X1  g473(.A1(new_n310), .A2(KEYINPUT38), .A3(new_n311), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT38), .B1(new_n310), .B2(new_n311), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n187), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n360), .B1(new_n355), .B2(new_n362), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n375), .A2(new_n360), .A3(new_n362), .ZN(new_n666));
  OR3_X1    g480(.A1(new_n665), .A2(KEYINPUT106), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT106), .B1(new_n665), .B2(new_n666), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n667), .A2(new_n297), .A3(new_n668), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n647), .A2(new_n648), .B1(new_n669), .B2(new_n316), .ZN(new_n670));
  INV_X1    g484(.A(new_n639), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n568), .A2(new_n593), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n253), .ZN(G45));
  AND3_X1   g490(.A1(new_n568), .A2(new_n616), .A3(new_n652), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n649), .A2(new_n650), .A3(new_n312), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  INV_X1    g493(.A(new_n501), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n500), .B1(new_n499), .B2(new_n297), .ZN(new_n681));
  INV_X1    g495(.A(new_n505), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n649), .A2(new_n622), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n619), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT41), .B(G113), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NOR2_X1   g501(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n505), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n400), .A2(new_n689), .A3(new_n462), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n630), .A3(new_n631), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  AND2_X1   g506(.A1(new_n639), .A2(new_n603), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n649), .A2(new_n312), .A3(new_n683), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  AND3_X1   g509(.A1(new_n312), .A2(new_n673), .A3(new_n683), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n388), .A2(new_n389), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n382), .A2(new_n371), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n395), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n622), .A2(new_n601), .A3(new_n623), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  AND3_X1   g517(.A1(new_n623), .A2(new_n699), .A3(new_n639), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n312), .A3(new_n677), .A4(new_n683), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  NAND2_X1  g520(.A1(new_n396), .A2(new_n399), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n462), .B1(new_n707), .B2(new_n646), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n310), .A2(new_n187), .A3(new_n311), .A4(new_n677), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n506), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n708), .A2(new_n710), .A3(KEYINPUT42), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT42), .B1(new_n708), .B2(new_n710), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G131), .ZN(G33));
  NAND2_X1  g528(.A1(new_n310), .A2(new_n311), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n308), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n708), .A2(new_n656), .A3(new_n653), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G134), .ZN(G36));
  INV_X1    g532(.A(new_n716), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n607), .A2(KEYINPUT108), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n568), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n616), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT43), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n617), .A2(KEYINPUT43), .A3(new_n568), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT109), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n640), .A2(new_n639), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n719), .B1(new_n730), .B2(KEYINPUT44), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n492), .A2(KEYINPUT45), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n492), .A2(new_n733), .A3(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n492), .B2(KEYINPUT45), .ZN(new_n735));
  OAI211_X1 g549(.A(G469), .B(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n502), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT46), .B1(new_n736), .B2(new_n502), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n680), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n682), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n657), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n731), .B(new_n741), .C1(KEYINPUT44), .C2(new_n730), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G137), .ZN(G39));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n744), .B1(new_n739), .B2(new_n682), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n738), .A2(new_n680), .ZN(new_n746));
  OAI211_X1 g560(.A(KEYINPUT47), .B(new_n505), .C1(new_n746), .C2(new_n737), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n709), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n400), .A3(new_n462), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G140), .ZN(G42));
  OR4_X1    g564(.A1(new_n308), .A2(new_n723), .A3(new_n462), .A4(new_n682), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n688), .B(KEYINPUT49), .Z(new_n752));
  OR4_X1    g566(.A1(new_n663), .A2(new_n751), .A3(new_n752), .A4(new_n670), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n618), .A2(new_n631), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n315), .A2(new_n601), .A3(new_n626), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n642), .A2(new_n756), .A3(new_n604), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n503), .A2(new_n639), .A3(new_n505), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n400), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n607), .A2(new_n592), .A3(new_n652), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n716), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n717), .B(new_n763), .C1(new_n711), .C2(new_n712), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n312), .A2(new_n673), .A3(new_n683), .ZN(new_n766));
  OAI22_X1  g580(.A1(new_n684), .A2(new_n619), .B1(new_n700), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n312), .A2(new_n601), .A3(new_n631), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n694), .B1(new_n684), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n308), .B(new_n672), .C1(new_n310), .C2(new_n311), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n503), .A2(new_n505), .A3(new_n652), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n670), .A3(new_n671), .A4(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n654), .A3(new_n678), .A4(new_n705), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n759), .B(new_n312), .C1(new_n653), .C2(new_n677), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT52), .A3(new_n705), .A4(new_n773), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n710), .A2(new_n780), .A3(new_n704), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n780), .B1(new_n710), .B2(new_n704), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n765), .A2(new_n770), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n764), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n642), .A2(new_n756), .A3(new_n604), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n779), .A2(new_n792), .A3(new_n793), .A4(new_n784), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT53), .A4(new_n770), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n785), .B2(new_n786), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n754), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n727), .A2(new_n596), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n622), .A2(new_n623), .A3(new_n699), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n312), .A2(new_n800), .A3(new_n683), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n719), .A2(new_n689), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n800), .A3(new_n708), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT48), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n719), .A2(new_n670), .A3(new_n689), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n462), .A2(new_n596), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n618), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n805), .A2(KEYINPUT48), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(new_n809), .A3(new_n594), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n727), .A2(new_n596), .A3(new_n801), .ZN(new_n812));
  INV_X1    g626(.A(new_n662), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n683), .A2(new_n308), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n813), .A2(new_n660), .B1(new_n814), .B2(KEYINPUT117), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n683), .A2(new_n816), .A3(new_n308), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n812), .A2(KEYINPUT50), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n662), .B2(new_n661), .ZN(new_n821));
  INV_X1    g635(.A(new_n596), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n725), .B1(new_n723), .B2(KEYINPUT43), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n802), .A2(new_n822), .A3(new_n823), .A4(new_n817), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n819), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n804), .A2(new_n800), .A3(new_n704), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n807), .A2(new_n607), .A3(new_n617), .A4(new_n808), .ZN(new_n828));
  AND4_X1   g642(.A1(KEYINPUT51), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n812), .A2(new_n716), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT115), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n688), .A2(new_n682), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n745), .A2(new_n747), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n811), .B1(new_n835), .B2(KEYINPUT118), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n829), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n831), .A2(new_n839), .A3(new_n833), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n831), .B2(new_n833), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n836), .B(new_n838), .C1(new_n843), .C2(KEYINPUT51), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n757), .A2(new_n764), .A3(new_n783), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n690), .A2(new_n620), .B1(new_n696), .B2(new_n701), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n691), .A4(new_n694), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n767), .B2(new_n769), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n850), .A3(KEYINPUT53), .A4(new_n779), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n787), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n799), .A2(new_n803), .A3(new_n844), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n753), .B1(new_n854), .B2(new_n855), .ZN(G75));
  AOI21_X1  g670(.A(new_n297), .B1(new_n787), .B2(new_n851), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT56), .B1(new_n857), .B2(new_n189), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n252), .B(new_n281), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT55), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n858), .A2(new_n861), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n279), .A2(G952), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G51));
  XOR2_X1   g679(.A(new_n502), .B(KEYINPUT57), .Z(new_n866));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n852), .B2(KEYINPUT54), .ZN(new_n868));
  AOI211_X1 g682(.A(KEYINPUT120), .B(new_n754), .C1(new_n787), .C2(new_n851), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n852), .B2(KEYINPUT54), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n787), .A2(new_n851), .A3(KEYINPUT119), .A4(new_n754), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n866), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n499), .ZN(new_n876));
  INV_X1    g690(.A(new_n736), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n857), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n864), .B1(new_n876), .B2(new_n878), .ZN(G54));
  AND2_X1   g693(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n566), .B1(new_n880), .B2(G475), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .A4(new_n566), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n864), .B(new_n881), .C1(new_n884), .C2(new_n885), .ZN(G60));
  NOR2_X1   g700(.A1(new_n608), .A2(new_n610), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n798), .A2(new_n788), .A3(new_n790), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n853), .B1(new_n888), .B2(KEYINPUT54), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n590), .A2(new_n297), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n890), .B(new_n891), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n887), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n864), .ZN(new_n895));
  INV_X1    g709(.A(new_n887), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n892), .C1(new_n870), .C2(new_n874), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(G63));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT60), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n787), .B2(new_n851), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n637), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n902), .B(new_n895), .C1(new_n443), .C2(new_n901), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g718(.A(new_n279), .B1(new_n599), .B2(G224), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n793), .A2(new_n770), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n279), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT123), .ZN(new_n908));
  INV_X1    g722(.A(new_n252), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(G898), .B2(new_n279), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n908), .B(new_n910), .ZN(G69));
  NAND3_X1  g725(.A1(new_n741), .A2(new_n708), .A3(new_n771), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n912), .A2(new_n713), .A3(new_n717), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n777), .A2(new_n705), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n913), .A2(new_n742), .A3(new_n749), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n279), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n340), .A2(new_n344), .A3(new_n354), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n552), .B1(new_n551), .B2(new_n554), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(KEYINPUT124), .B(G900), .Z(new_n924));
  AOI21_X1  g738(.A(new_n919), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT125), .Z(new_n926));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n675), .B2(new_n914), .ZN(new_n928));
  OAI211_X1 g742(.A(KEYINPUT62), .B(new_n915), .C1(new_n664), .C2(new_n674), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n656), .A2(new_n657), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(new_n708), .A3(new_n716), .A4(new_n755), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n930), .A2(new_n742), .A3(new_n749), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n279), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n923), .B(new_n926), .C1(new_n922), .C2(new_n934), .ZN(G72));
  XNOR2_X1  g749(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n316), .A2(new_n297), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT127), .Z(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n933), .B2(new_n906), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n665), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n916), .B2(new_n906), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n364), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n943), .A3(new_n895), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n363), .A2(new_n938), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n665), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n888), .B2(new_n946), .ZN(G57));
endmodule


