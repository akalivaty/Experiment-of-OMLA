//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT74), .A4(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT75), .B(G101), .C1(new_n194), .C2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n196), .A2(G104), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n190), .B2(new_n192), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(KEYINPUT74), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n195), .A2(KEYINPUT74), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n203), .A3(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(new_n207), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT75), .B1(new_n210), .B2(G101), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT76), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n194), .B2(new_n199), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n214), .A3(new_n217), .A4(new_n200), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n220), .B2(G119), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G116), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G119), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT2), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G113), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n230), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n221), .A3(new_n224), .A4(new_n225), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT67), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n237), .B(new_n238), .C1(KEYINPUT4), .C2(new_n215), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n219), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n198), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n206), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n198), .A2(new_n242), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n208), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n220), .A2(G119), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n227), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n226), .B2(new_n249), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n234), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(G110), .B(G122), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n241), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n255), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n239), .B1(new_n212), .B2(new_n218), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(new_n253), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n259), .A3(KEYINPUT6), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(new_n257), .C1(new_n258), .C2(new_n253), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT0), .A3(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  INV_X1    g082(.A(G146), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G143), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n265), .B(new_n266), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G125), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n263), .A2(new_n274), .A3(G128), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n269), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(KEYINPUT65), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n268), .B2(new_n270), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n275), .A2(new_n276), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n273), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G953), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n287), .A2(G224), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n260), .A2(new_n262), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(KEYINPUT80), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n273), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n285), .A2(KEYINPUT80), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  OAI22_X1  g109(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n288), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n255), .B(KEYINPUT8), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n208), .A2(new_n246), .B1(new_n251), .B2(new_n234), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n253), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n288), .A2(new_n295), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n273), .A2(new_n285), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n256), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n291), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI211_X1 g119(.A(KEYINPUT81), .B(G902), .C1(new_n256), .C2(new_n302), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n290), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n253), .B1(new_n219), .B2(new_n240), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(new_n255), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT81), .B1(new_n313), .B2(G902), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n258), .A2(new_n253), .A3(new_n257), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n291), .B(new_n304), .C1(new_n315), .C2(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n308), .A3(new_n290), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n188), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n320));
  NOR2_X1   g134(.A1(G475), .A2(G902), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT86), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G113), .B(G122), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT84), .B(G104), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n326), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n276), .A2(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT82), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT19), .A3(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n334), .A2(KEYINPUT19), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n269), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G143), .B1(new_n343), .B2(G214), .ZN(new_n346));
  OAI21_X1  g160(.A(G131), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G237), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n287), .A3(G214), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n267), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n344), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT16), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n331), .A3(G125), .ZN(new_n355));
  OAI211_X1 g169(.A(G146), .B(new_n355), .C1(new_n334), .C2(new_n354), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n338), .A2(KEYINPUT83), .A3(new_n269), .A4(new_n339), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n342), .A2(new_n353), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n332), .A2(new_n333), .A3(new_n269), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT72), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n336), .A2(G146), .A3(new_n337), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n350), .A2(new_n344), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n350), .B2(new_n344), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n330), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT17), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n347), .A2(new_n369), .A3(new_n352), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n351), .B1(new_n350), .B2(new_n344), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT17), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n355), .B1(new_n334), .B2(new_n354), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n269), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n374), .A4(new_n356), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n330), .A2(KEYINPUT85), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n328), .A2(new_n377), .A3(new_n329), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n367), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n320), .B(new_n323), .C1(new_n368), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n375), .A3(new_n379), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n345), .A2(new_n346), .A3(G131), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n356), .B1(new_n385), .B2(new_n371), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n341), .B2(new_n340), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n387), .A2(new_n357), .B1(new_n362), .B2(new_n366), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n384), .B1(new_n388), .B2(new_n330), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(KEYINPUT87), .A3(new_n320), .A4(new_n323), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n358), .A2(new_n367), .ZN(new_n391));
  INV_X1    g205(.A(new_n330), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n380), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n393), .B2(new_n322), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n383), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n330), .B1(new_n367), .B2(new_n375), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n304), .B1(new_n380), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G475), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n395), .B2(new_n399), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT89), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(G116), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n220), .A2(KEYINPUT89), .A3(G122), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n220), .B2(G122), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n407), .A2(G107), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n267), .A2(G128), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n283), .A2(G143), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT64), .ZN(new_n412));
  INV_X1    g226(.A(G134), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT64), .A2(G134), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n411), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n404), .A2(new_n405), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(new_n220), .B2(G122), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n420), .B2(new_n419), .ZN(new_n422));
  OAI221_X1 g236(.A(new_n408), .B1(new_n417), .B2(new_n418), .C1(new_n422), .C2(new_n196), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n407), .B(G107), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n407), .A2(G107), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n408), .A2(KEYINPUT90), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n267), .A2(KEYINPUT13), .A3(G128), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT91), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n413), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n409), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(new_n429), .A3(KEYINPUT91), .A4(new_n410), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n417), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n426), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  INV_X1    g252(.A(G217), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(G953), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n423), .A2(new_n436), .A3(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G478), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n304), .C1(KEYINPUT15), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n443), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n440), .B1(new_n423), .B2(new_n436), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n304), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n445), .A2(KEYINPUT15), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n287), .A2(G952), .ZN(new_n452));
  INV_X1    g266(.A(G234), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(new_n348), .ZN(new_n454));
  OAI211_X1 g268(.A(G902), .B(G953), .C1(new_n453), .C2(new_n348), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT92), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(G898), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n446), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n400), .A2(new_n401), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n272), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n215), .B2(KEYINPUT4), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n219), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT10), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n275), .A2(new_n284), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n267), .A2(G146), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n280), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n469), .A2(new_n470), .B1(new_n275), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n468), .B1(new_n473), .B2(new_n247), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n246), .A2(new_n208), .ZN(new_n475));
  INV_X1    g289(.A(new_n274), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n269), .A2(G143), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n471), .A3(G128), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n282), .B(new_n284), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(KEYINPUT10), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT11), .ZN(new_n483));
  INV_X1    g297(.A(G137), .ZN(new_n484));
  AND2_X1   g298(.A1(KEYINPUT64), .A2(G134), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT64), .A2(G134), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(G134), .B2(new_n484), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n414), .A2(G137), .A3(new_n415), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n351), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n351), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n489), .B2(new_n487), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n467), .A2(new_n482), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT79), .B1(new_n475), .B2(new_n479), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT78), .B1(new_n275), .B2(new_n284), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n275), .A2(new_n472), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n475), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n479), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n247), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n495), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n504), .A2(KEYINPUT12), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT12), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G110), .B(G140), .ZN(new_n509));
  INV_X1    g323(.A(G227), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n509), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n465), .B1(new_n212), .B2(new_n218), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n481), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n512), .B1(new_n514), .B2(new_n495), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n505), .B1(new_n513), .B2(new_n481), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n508), .A2(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G469), .B1(new_n517), .B2(G902), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n496), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n512), .ZN(new_n520));
  INV_X1    g334(.A(new_n512), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n496), .B(new_n521), .C1(new_n506), .C2(new_n507), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G469), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n304), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n463), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n319), .A2(new_n461), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n374), .A2(new_n356), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n223), .B2(G128), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n283), .A2(KEYINPUT23), .A3(G119), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n534), .C1(G119), .C2(new_n283), .ZN(new_n535));
  XNOR2_X1  g349(.A(G119), .B(G128), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT24), .B(G110), .Z(new_n537));
  AOI22_X1  g351(.A1(new_n535), .A2(G110), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n535), .A2(G110), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT71), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n540), .A2(new_n541), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n541), .B2(new_n540), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n360), .A2(new_n356), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n287), .A2(G221), .A3(G234), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n546), .B(new_n547), .Z(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n539), .B(new_n548), .C1(new_n543), .C2(new_n544), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n530), .B1(new_n552), .B2(new_n304), .ZN(new_n553));
  NAND2_X1  g367(.A1(G217), .A2(G902), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n439), .B2(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT70), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n304), .A3(new_n551), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(KEYINPUT25), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n556), .A2(G902), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT73), .Z(new_n561));
  AND2_X1   g375(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n485), .A2(new_n486), .ZN(new_n566));
  AOI21_X1  g380(.A(G131), .B1(new_n566), .B2(G137), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n490), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n413), .A2(G137), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G131), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n479), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n238), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT67), .B1(new_n232), .B2(new_n234), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(G137), .B1(new_n414), .B2(new_n415), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n488), .B1(new_n577), .B2(new_n483), .ZN(new_n578));
  INV_X1    g392(.A(new_n491), .ZN(new_n579));
  OAI21_X1  g393(.A(G131), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n272), .B1(new_n580), .B2(new_n568), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT68), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n490), .A2(new_n567), .B1(new_n571), .B2(G131), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n237), .A2(new_n238), .B1(new_n584), .B2(new_n479), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n464), .B1(new_n492), .B2(new_n494), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT68), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n574), .A2(new_n575), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT30), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n586), .A2(new_n590), .A3(new_n573), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n586), .B2(new_n573), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT31), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n343), .A2(G210), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT27), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT26), .B(G101), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n588), .A2(new_n593), .A3(new_n594), .A4(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n582), .B1(new_n576), .B2(new_n581), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n237), .A2(new_n238), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n586), .A2(new_n601), .A3(KEYINPUT68), .A4(new_n573), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n602), .A3(new_n598), .ZN(new_n603));
  INV_X1    g417(.A(new_n573), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT30), .B1(new_n581), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n586), .A2(new_n590), .A3(new_n573), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT31), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n589), .B1(new_n581), .B2(new_n604), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n600), .A2(new_n610), .A3(new_n602), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT28), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT28), .B1(new_n585), .B2(new_n586), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n598), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT69), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n599), .A2(new_n608), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n598), .B1(new_n612), .B2(new_n614), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT69), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n565), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT32), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n609), .A2(KEYINPUT69), .A3(new_n617), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n621), .B1(new_n619), .B2(new_n620), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n565), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n624), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n600), .A2(new_n602), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n607), .A2(new_n631), .A3(new_n598), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT29), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n615), .A2(KEYINPUT29), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n613), .B1(new_n611), .B2(KEYINPUT28), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n598), .B1(new_n636), .B2(new_n633), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n628), .A2(new_n630), .B1(G472), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n564), .B1(new_n625), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n319), .A2(new_n461), .A3(KEYINPUT93), .A4(new_n526), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n529), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  NAND2_X1  g457(.A1(new_n526), .A2(new_n563), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n626), .B2(new_n627), .ZN(new_n645));
  INV_X1    g459(.A(G472), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n629), .B1(new_n626), .B2(new_n627), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n317), .A2(new_n308), .A3(new_n290), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n308), .B1(new_n317), .B2(new_n290), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n459), .B(new_n187), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n444), .A2(KEYINPUT33), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n442), .A2(new_n656), .A3(new_n443), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(G478), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n444), .A2(new_n445), .A3(new_n304), .ZN(new_n659));
  NAND2_X1  g473(.A1(G478), .A2(G902), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n400), .B2(new_n401), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n446), .A2(new_n451), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n394), .A2(new_n381), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n399), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n654), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT35), .B(G107), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  OR2_X1    g485(.A1(new_n645), .A2(new_n646), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT94), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n549), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n545), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n561), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n553), .B2(new_n558), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n672), .A2(new_n673), .A3(new_n623), .A4(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n623), .B(new_n677), .C1(new_n645), .C2(new_n646), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n529), .A2(new_n678), .A3(new_n641), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT37), .B(G110), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT95), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(new_n677), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n625), .B2(new_n639), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n187), .B1(new_n650), .B2(new_n651), .ZN(new_n687));
  AOI211_X1 g501(.A(G469), .B(G902), .C1(new_n520), .C2(new_n522), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n496), .A2(new_n516), .A3(new_n521), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n479), .B1(new_n208), .B2(new_n246), .ZN(new_n690));
  OAI22_X1  g504(.A1(new_n690), .A2(new_n502), .B1(new_n473), .B2(new_n247), .ZN(new_n691));
  INV_X1    g505(.A(new_n503), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n505), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT12), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n504), .A2(KEYINPUT12), .A3(new_n505), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n695), .A2(new_n696), .B1(new_n514), .B2(new_n495), .ZN(new_n697));
  OAI211_X1 g511(.A(G469), .B(new_n689), .C1(new_n697), .C2(new_n521), .ZN(new_n698));
  NAND2_X1  g512(.A1(G469), .A2(G902), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n462), .B1(new_n688), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n687), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n686), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n666), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT96), .B(G900), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n454), .B1(new_n456), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT97), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n667), .A2(new_n399), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  NOR2_X1   g526(.A1(new_n650), .A2(new_n651), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT38), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n715), .A2(new_n187), .A3(new_n685), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n707), .B(KEYINPUT39), .Z(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT40), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n666), .B1(new_n400), .B2(new_n401), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n630), .B1(new_n618), .B2(new_n622), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n611), .A2(new_n616), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n603), .A2(new_n607), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n728), .B2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n625), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n716), .A2(new_n720), .A3(new_n722), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  OAI211_X1 g546(.A(new_n661), .B(new_n708), .C1(new_n400), .C2(new_n401), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n703), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  INV_X1    g550(.A(KEYINPUT100), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n638), .A2(G472), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n723), .B(new_n738), .C1(new_n648), .C2(KEYINPUT32), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n695), .A2(new_n696), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n519), .A2(new_n512), .B1(new_n515), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(G469), .B1(new_n741), .B2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n462), .A3(new_n525), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT99), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT99), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n525), .A3(new_n745), .A4(new_n462), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n739), .A2(new_n563), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n748));
  INV_X1    g562(.A(new_n401), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n319), .A3(new_n459), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n737), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n744), .A2(new_n746), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n652), .A2(new_n662), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n640), .A3(new_n755), .A4(KEYINPUT100), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NOR2_X1   g573(.A1(new_n652), .A2(new_n668), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(new_n640), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G116), .ZN(G18));
  INV_X1    g576(.A(KEYINPUT101), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n687), .A2(new_n763), .A3(new_n743), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n742), .A2(new_n462), .A3(new_n525), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT101), .B1(new_n319), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n461), .B(new_n686), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  INV_X1    g582(.A(KEYINPUT102), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n617), .B2(new_n608), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n608), .B(new_n769), .C1(new_n636), .C2(new_n598), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n599), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n565), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n563), .B(new_n773), .C1(new_n645), .C2(new_n646), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n687), .A2(new_n721), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n754), .A2(new_n459), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  OAI211_X1 g592(.A(new_n773), .B(new_n677), .C1(new_n645), .C2(new_n646), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n733), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n764), .B2(new_n766), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  NAND3_X1  g596(.A1(new_n310), .A2(new_n187), .A3(new_n318), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n701), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n640), .A2(new_n734), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT103), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n640), .A2(KEYINPUT103), .A3(new_n734), .A4(new_n784), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT42), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT104), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n625), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT32), .B1(new_n628), .B2(new_n565), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT104), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n639), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n563), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n784), .A2(new_n734), .A3(KEYINPUT42), .ZN(new_n797));
  OAI22_X1  g611(.A1(new_n787), .A2(new_n790), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT105), .B(G131), .Z(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G33));
  NAND4_X1  g614(.A1(new_n784), .A2(new_n739), .A3(new_n563), .A4(new_n710), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT106), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n640), .A2(KEYINPUT106), .A3(new_n710), .A4(new_n784), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  OR2_X1    g620(.A1(new_n517), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n517), .A2(KEYINPUT45), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(G469), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT46), .A3(new_n699), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT107), .Z(new_n811));
  AOI21_X1  g625(.A(KEYINPUT46), .B1(new_n809), .B2(new_n699), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n688), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n462), .A3(new_n717), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT108), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n463), .B1(new_n811), .B2(new_n813), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT108), .A3(new_n717), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n400), .A2(new_n401), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n661), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT43), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT43), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT109), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT109), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n685), .B1(new_n672), .B2(new_n623), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(KEYINPUT44), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n783), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT110), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT44), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n820), .A2(new_n832), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G137), .ZN(G39));
  NOR4_X1   g653(.A1(new_n739), .A2(new_n733), .A3(new_n563), .A4(new_n783), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT47), .B1(new_n814), .B2(new_n462), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n842), .B(new_n463), .C1(new_n811), .C2(new_n813), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G140), .ZN(G42));
  NAND2_X1  g659(.A1(new_n742), .A2(new_n525), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT111), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT49), .Z(new_n848));
  NOR4_X1   g662(.A1(new_n715), .A2(new_n564), .A3(new_n188), .A4(new_n463), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n730), .A2(new_n822), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n841), .A2(new_n843), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n463), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n825), .A2(new_n454), .A3(new_n774), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n830), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n715), .A2(new_n187), .A3(new_n743), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n783), .A2(new_n454), .A3(new_n743), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n823), .A2(new_n824), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n779), .ZN(new_n867));
  INV_X1    g681(.A(new_n730), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n563), .A3(new_n865), .ZN(new_n869));
  INV_X1    g683(.A(new_n821), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n869), .A2(new_n870), .A3(new_n661), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n863), .A2(new_n864), .A3(new_n867), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n858), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n858), .A2(new_n872), .A3(KEYINPUT51), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n452), .B1(new_n869), .B2(new_n662), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n796), .A2(new_n866), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT48), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n764), .A2(new_n766), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n877), .B(new_n879), .C1(new_n880), .C2(new_n857), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT112), .B1(new_n652), .B2(new_n662), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n751), .A2(new_n319), .A3(new_n884), .A4(new_n459), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n649), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n642), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n642), .B2(new_n886), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n870), .A2(new_n704), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n649), .A2(new_n653), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n681), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n767), .A2(new_n761), .A3(new_n777), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n753), .B2(new_n756), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n686), .B(new_n702), .C1(new_n710), .C2(new_n734), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n685), .A2(new_n708), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n730), .A2(new_n702), .A3(new_n722), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n781), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n896), .A2(new_n781), .A3(new_n899), .A4(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n893), .A2(new_n895), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n902), .A2(new_n903), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(KEYINPUT116), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n796), .A2(new_n797), .ZN(new_n909));
  INV_X1    g723(.A(new_n790), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n785), .A2(new_n786), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n779), .A2(new_n733), .A3(new_n783), .A4(new_n701), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT114), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n723), .A2(new_n738), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n677), .B1(new_n916), .B2(new_n793), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n666), .A2(new_n709), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n713), .A2(new_n526), .A3(new_n187), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n918), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n783), .A2(new_n701), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n686), .A2(new_n922), .A3(KEYINPUT114), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n913), .B1(new_n924), .B2(new_n805), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n805), .A3(new_n913), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n912), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n905), .A2(new_n908), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n908), .B1(new_n905), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT54), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n931), .A2(KEYINPUT117), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n753), .A2(new_n756), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT118), .B1(new_n933), .B2(new_n894), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n767), .A2(new_n761), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n757), .A3(new_n936), .A4(new_n777), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n934), .A2(KEYINPUT53), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n642), .A2(new_n886), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT113), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n642), .A2(new_n886), .A3(new_n887), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n940), .A2(new_n681), .A3(new_n941), .A4(new_n891), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n907), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n928), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n889), .A2(new_n892), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n904), .A2(new_n895), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n924), .A2(new_n805), .A3(new_n913), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n798), .B1(new_n947), .B2(new_n925), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n906), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n931), .B(KEYINPUT117), .C1(KEYINPUT54), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n882), .B1(new_n932), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(G952), .A2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n851), .B1(new_n952), .B2(new_n953), .ZN(G75));
  AOI21_X1  g768(.A(new_n304), .B1(new_n944), .B2(new_n949), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(G210), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(KEYINPUT56), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n260), .A2(new_n262), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n289), .ZN(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n287), .A2(G952), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n962), .A2(new_n967), .ZN(G51));
  XNOR2_X1  g782(.A(new_n950), .B(KEYINPUT54), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n699), .B(KEYINPUT57), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n523), .B(KEYINPUT123), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n809), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n955), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n963), .B1(new_n973), .B2(new_n975), .ZN(G54));
  NAND3_X1  g790(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n393), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n393), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n963), .ZN(G60));
  AND2_X1   g794(.A1(new_n655), .A2(new_n657), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n660), .B(KEYINPUT59), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n969), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n964), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n932), .A2(new_n951), .A3(new_n983), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n981), .B2(new_n987), .ZN(G63));
  XNOR2_X1  g802(.A(new_n554), .B(KEYINPUT60), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT53), .B1(new_n905), .B2(new_n928), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n934), .A2(KEYINPUT53), .A3(new_n937), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n904), .A2(new_n941), .A3(new_n945), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n992), .A2(new_n948), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT124), .ZN(new_n996));
  INV_X1    g810(.A(new_n552), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n950), .A2(new_n998), .A3(new_n990), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(new_n950), .B2(new_n990), .ZN(new_n1001));
  AOI211_X1 g815(.A(KEYINPUT124), .B(new_n989), .C1(new_n944), .C2(new_n949), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n675), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1000), .A2(new_n1003), .A3(new_n964), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1000), .A2(new_n1003), .A3(KEYINPUT61), .A4(new_n964), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(G66));
  AOI21_X1  g822(.A(new_n287), .B1(new_n458), .B2(G224), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n893), .A2(new_n895), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n287), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n958), .B1(G898), .B2(new_n287), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(G69));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n896), .A2(new_n781), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n731), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n731), .A2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  INV_X1    g832(.A(new_n890), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n718), .B1(new_n1019), .B2(new_n662), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n640), .A3(new_n784), .ZN(new_n1021));
  AND4_X1   g835(.A1(new_n844), .A2(new_n1016), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(G953), .B1(new_n838), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n605), .A2(new_n606), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n338), .A2(new_n339), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1024), .B(new_n1025), .Z(new_n1026));
  AOI21_X1  g840(.A(new_n287), .B1(G227), .B2(G900), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n798), .A2(new_n805), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT125), .Z(new_n1030));
  NOR3_X1   g844(.A1(new_n796), .A2(new_n687), .A3(new_n721), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n817), .A2(new_n819), .A3(new_n1031), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n1032), .A2(new_n844), .A3(new_n1015), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1030), .A2(new_n1033), .A3(new_n838), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n287), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n510), .A2(G900), .A3(G953), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1028), .B1(new_n1037), .B2(new_n1026), .ZN(G72));
  NAND2_X1  g852(.A1(G472), .A2(G902), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT63), .Z(new_n1040));
  OAI21_X1  g854(.A(new_n1040), .B1(new_n1034), .B2(new_n1010), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n632), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1010), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n838), .A2(new_n1022), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n1040), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n616), .B1(new_n588), .B2(new_n593), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n963), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(new_n632), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n1040), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1049), .A2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1050), .B1(new_n929), .B2(new_n930), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1042), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(KEYINPUT126), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT126), .ZN(new_n1054));
  NAND4_X1  g868(.A1(new_n1042), .A2(new_n1047), .A3(new_n1054), .A4(new_n1051), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1055), .ZN(G57));
endmodule


