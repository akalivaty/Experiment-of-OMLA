//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT71), .B(G902), .Z(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT65), .A2(G953), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT65), .A2(G953), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(G221), .A2(G234), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT75), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OR4_X1    g011(.A1(KEYINPUT75), .A2(new_n192), .A3(new_n193), .A4(new_n196), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n191), .A3(new_n198), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(KEYINPUT76), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT76), .ZN(new_n203));
  INV_X1    g017(.A(new_n201), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(new_n199), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT24), .B(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n209), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n216), .B2(G110), .ZN(new_n217));
  INV_X1    g031(.A(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G125), .ZN(new_n219));
  INV_X1    g033(.A(G125), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n217), .B1(G146), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT73), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G125), .B(G140), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT73), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT16), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n218), .A3(G125), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n225), .A2(G146), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT74), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n223), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n210), .A2(new_n211), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(G110), .B2(new_n216), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n240), .B2(new_n230), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n202), .B(new_n205), .C1(new_n234), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n230), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n236), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n200), .A2(new_n201), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n230), .B(KEYINPUT74), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n244), .B(new_n245), .C1(new_n246), .C2(new_n223), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n247), .A3(new_n188), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n249), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n242), .A2(new_n247), .A3(new_n188), .A4(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n190), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n189), .A2(G902), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n242), .A2(new_n247), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(G137), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n261), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n260), .A2(G137), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n262), .A2(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n239), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n239), .A2(G143), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n277), .A2(new_n206), .B1(KEYINPUT1), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n270), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n261), .A2(new_n265), .A3(new_n263), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT0), .B(G128), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n282), .A2(new_n266), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n258), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT64), .A2(G116), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT64), .A2(G116), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(G119), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n208), .A2(G116), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT2), .B(G113), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n291), .A3(new_n292), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n282), .A2(new_n266), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n284), .A2(new_n286), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n273), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n271), .B2(G128), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n266), .B(new_n269), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n305), .A3(KEYINPUT30), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n288), .A2(new_n298), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n194), .A2(G210), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(new_n314), .A3(new_n312), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n297), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n294), .B1(new_n292), .B2(new_n291), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n301), .A3(new_n305), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n307), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT31), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n321), .A2(new_n301), .A3(KEYINPUT28), .A4(new_n305), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n298), .B1(new_n280), .B2(new_n287), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n316), .A2(new_n317), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n307), .A2(new_n332), .A3(new_n318), .A4(new_n322), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n324), .A2(KEYINPUT67), .A3(new_n331), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(G472), .A2(G902), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(KEYINPUT68), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n343));
  INV_X1    g157(.A(new_n339), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n336), .B2(new_n337), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n343), .B1(new_n345), .B2(KEYINPUT32), .ZN(new_n346));
  INV_X1    g160(.A(G472), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n330), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n328), .A2(new_n322), .A3(KEYINPUT70), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT70), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n298), .B(new_n351), .C1(new_n280), .C2(new_n287), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n353), .A3(new_n326), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n354), .A2(new_n188), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT69), .B1(new_n329), .B2(new_n330), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n321), .B1(new_n301), .B2(new_n305), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n325), .B2(new_n322), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT69), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n318), .A4(new_n327), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n307), .A2(new_n322), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n330), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n356), .A2(new_n360), .A3(new_n348), .A4(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n347), .B1(new_n355), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n345), .B2(KEYINPUT32), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n342), .A2(new_n346), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT72), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n342), .A2(new_n346), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n257), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G122), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n298), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n387), .B2(G101), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(G104), .B2(new_n379), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT78), .B(G107), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n378), .ZN(new_n395));
  AOI21_X1  g209(.A(G101), .B1(new_n377), .B2(G107), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT79), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n385), .A4(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n383), .A2(new_n385), .A3(new_n396), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n398), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n390), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n384), .B1(new_n394), .B2(G104), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n291), .A2(KEYINPUT5), .A3(new_n292), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n413));
  INV_X1    g227(.A(G113), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n297), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n376), .B1(new_n408), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n390), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT80), .B1(new_n406), .B2(new_n391), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n418), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n375), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n419), .A2(KEYINPUT6), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT81), .B(G224), .Z(new_n427));
  INV_X1    g241(.A(G953), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(G125), .B1(new_n279), .B2(new_n273), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n220), .B1(new_n284), .B2(new_n286), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n220), .B1(new_n302), .B2(new_n304), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n300), .A2(G125), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n429), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(new_n376), .C1(new_n408), .C2(new_n418), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n426), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n430), .A2(KEYINPUT7), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n433), .B2(new_n436), .ZN(new_n442));
  AOI211_X1 g256(.A(KEYINPUT7), .B(new_n430), .C1(new_n434), .C2(new_n435), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n402), .A2(new_n407), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n418), .B1(new_n445), .B2(new_n420), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n446), .B2(new_n375), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n375), .B(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(KEYINPUT83), .B(new_n410), .C1(new_n397), .C2(new_n399), .ZN(new_n451));
  INV_X1    g265(.A(new_n417), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n405), .A2(new_n398), .B1(G101), .B2(new_n409), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n417), .B1(new_n454), .B2(KEYINPUT83), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n448), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n452), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n417), .A3(KEYINPUT83), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT84), .A4(new_n450), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n447), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n440), .B1(new_n461), .B2(KEYINPUT85), .ZN(new_n462));
  INV_X1    g276(.A(new_n444), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n425), .A2(new_n463), .A3(new_n456), .A4(new_n459), .ZN(new_n464));
  INV_X1    g278(.A(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n374), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n467), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n373), .A4(new_n440), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n372), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g287(.A1(KEYINPUT65), .A2(G953), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT65), .A2(G953), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n474), .A2(G214), .A3(new_n308), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n275), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n194), .A2(G143), .A3(G214), .A4(new_n308), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(KEYINPUT18), .A2(G131), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n226), .B(new_n239), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G113), .B(G122), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT86), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n377), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(KEYINPUT17), .A3(G131), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n240), .A3(new_n230), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n477), .A2(new_n478), .A3(new_n264), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n264), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n489), .A2(KEYINPUT87), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n488), .A2(new_n240), .A3(new_n495), .A4(new_n230), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n484), .B(new_n487), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n487), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n493), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n484), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n465), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G475), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n498), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n226), .B(KEYINPUT19), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n239), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n490), .B2(new_n491), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n246), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n487), .B1(new_n511), .B2(new_n484), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G475), .A2(G902), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n514), .ZN(new_n516));
  AOI211_X1 g330(.A(KEYINPUT20), .B(new_n516), .C1(new_n507), .C2(new_n512), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n505), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n188), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT9), .B(G234), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n520), .A2(new_n187), .A3(G953), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n275), .A2(G128), .ZN(new_n524));
  OR3_X1    g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n206), .A2(G143), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT90), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n524), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G134), .ZN(new_n531));
  INV_X1    g345(.A(new_n394), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n289), .A2(G122), .A3(new_n290), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G116), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(G122), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n536), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n394), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n260), .A3(new_n524), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(KEYINPUT88), .A3(new_n539), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n531), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n527), .A2(new_n524), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G134), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n543), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n538), .B1(new_n533), .B2(KEYINPUT14), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n533), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n548), .B(new_n539), .C1(new_n379), .C2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n521), .B1(new_n545), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n545), .A2(new_n555), .A3(new_n521), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n519), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n559), .A2(new_n560), .B1(KEYINPUT15), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n563));
  INV_X1    g377(.A(new_n558), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n556), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT93), .B(new_n563), .C1(new_n565), .C2(new_n519), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n560), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n428), .A2(G952), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(G234), .B2(G237), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT21), .B(G898), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT94), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI211_X1 g387(.A(new_n194), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n518), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n473), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G221), .B1(new_n520), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n300), .B(new_n389), .C1(new_n421), .C2(new_n422), .ZN(new_n580));
  INV_X1    g394(.A(new_n299), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n279), .A2(new_n273), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n406), .A2(new_n582), .A3(new_n410), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n454), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n580), .A2(new_n581), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n583), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n454), .A2(new_n582), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n299), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n582), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n411), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n581), .B1(new_n594), .B2(new_n583), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT12), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n587), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n194), .A2(G227), .ZN(new_n598));
  XOR2_X1   g412(.A(G110), .B(G140), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n389), .A2(new_n300), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n402), .B2(new_n407), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n585), .A2(new_n586), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(new_n604), .B2(new_n581), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n299), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n597), .A2(new_n600), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G469), .B1(new_n607), .B2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n587), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n600), .ZN(new_n610));
  INV_X1    g424(.A(new_n600), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n587), .B(new_n611), .C1(new_n592), .C2(new_n596), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G469), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n188), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n579), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n370), .A2(new_n577), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(new_n575), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n473), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT95), .B1(new_n545), .B2(new_n555), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n565), .A2(new_n623), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n564), .A2(new_n556), .B1(new_n621), .B2(new_n622), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n625), .A3(G478), .A4(new_n188), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n561), .B1(new_n565), .B2(new_n519), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n518), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n587), .A2(new_n606), .A3(new_n611), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n590), .A2(new_n591), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n595), .A2(KEYINPUT12), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n581), .A2(new_n604), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n631), .B1(new_n634), .B2(new_n611), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n614), .B1(new_n635), .B2(new_n465), .ZN(new_n636));
  AOI211_X1 g450(.A(G469), .B(new_n519), .C1(new_n610), .C2(new_n612), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n340), .B(new_n578), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n519), .B1(new_n336), .B2(new_n337), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n256), .B1(new_n347), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n630), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n513), .A2(new_n514), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT20), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n513), .A2(new_n506), .A3(new_n514), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(KEYINPUT96), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n515), .B2(new_n517), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n504), .A2(new_n652), .A3(G475), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n652), .B1(new_n504), .B2(G475), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n651), .A2(new_n568), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n620), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n641), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NAND2_X1  g474(.A1(new_n250), .A2(new_n252), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n189), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n205), .A2(new_n202), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT36), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n241), .B2(new_n234), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n234), .A2(new_n241), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n664), .A3(new_n663), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n254), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n578), .B(new_n671), .C1(new_n636), .C2(new_n637), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n338), .A2(new_n188), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n340), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n473), .A3(new_n576), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  NAND2_X1  g493(.A1(new_n469), .A2(new_n472), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n371), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n570), .B1(new_n574), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n651), .A2(new_n655), .A3(new_n568), .A4(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n681), .A2(new_n685), .A3(new_n672), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n367), .A2(new_n369), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XOR2_X1   g503(.A(new_n683), .B(KEYINPUT39), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n616), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT40), .Z(new_n692));
  OR2_X1    g506(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n693));
  INV_X1    g507(.A(new_n361), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n330), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n350), .A2(new_n352), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n330), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n347), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n345), .B2(KEYINPUT32), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n342), .A2(new_n346), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT98), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT98), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n342), .A2(new_n346), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT38), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n680), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n469), .A2(KEYINPUT38), .A3(new_n472), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n518), .A2(new_n568), .A3(new_n371), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n710), .A2(new_n671), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n693), .A2(new_n705), .A3(new_n706), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NOR2_X1   g529(.A1(new_n681), .A2(new_n672), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n518), .A2(new_n628), .A3(new_n684), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n518), .A2(new_n628), .A3(KEYINPUT100), .A4(new_n684), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n687), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  AOI21_X1  g538(.A(new_n614), .B1(new_n613), .B2(new_n188), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n637), .A3(new_n579), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n370), .A2(new_n630), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT41), .B(G113), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT101), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n727), .B(new_n729), .ZN(G15));
  NAND3_X1  g544(.A1(new_n370), .A2(new_n657), .A3(new_n726), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  AND4_X1   g546(.A1(new_n473), .A2(new_n726), .A3(new_n576), .A4(new_n671), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n687), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND2_X1  g549(.A1(new_n324), .A2(new_n333), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n318), .B1(new_n353), .B2(new_n326), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n339), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n674), .A2(new_n256), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n725), .A2(new_n637), .A3(new_n575), .A4(new_n579), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n680), .A4(new_n711), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT102), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND3_X1  g558(.A1(new_n674), .A2(new_n671), .A3(new_n738), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n721), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n726), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n681), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NAND3_X1  g564(.A1(new_n469), .A2(new_n371), .A3(new_n472), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n469), .A2(new_n753), .A3(new_n371), .A4(new_n472), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n616), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n752), .A2(KEYINPUT104), .A3(new_n616), .A4(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n370), .A3(new_n722), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n340), .A2(new_n341), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n257), .B1(new_n763), .B2(new_n365), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n722), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  INV_X1    g581(.A(new_n685), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n759), .A2(new_n370), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n518), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n646), .A2(new_n647), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(KEYINPUT105), .A3(new_n505), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n626), .B2(new_n627), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n774), .A3(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n628), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n777), .B1(new_n783), .B2(new_n518), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n675), .A2(new_n671), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n607), .A2(KEYINPUT45), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n635), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n793), .A3(G469), .ZN(new_n794));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n637), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n579), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n752), .A2(new_n754), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n800), .A2(new_n690), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n789), .A2(new_n790), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NOR2_X1   g619(.A1(new_n800), .A2(KEYINPUT107), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n807), .B(new_n579), .C1(new_n798), .C2(new_n799), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n809));
  NOR3_X1   g623(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n796), .A2(new_n797), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(new_n615), .A3(new_n799), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n807), .B1(new_n813), .B2(new_n579), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n800), .A2(KEYINPUT107), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n687), .A2(new_n801), .A3(new_n256), .A4(new_n721), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NOR2_X1   g634(.A1(new_n725), .A2(new_n637), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT109), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n783), .A2(new_n372), .A3(new_n579), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n775), .A2(new_n825), .A3(new_n256), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n702), .A3(new_n704), .A4(new_n710), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n367), .A2(new_n369), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n566), .A2(new_n562), .A3(new_n567), .A4(new_n684), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n651), .A2(new_n831), .A3(new_n655), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n672), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n754), .A3(new_n752), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n829), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n802), .A2(new_n687), .A3(KEYINPUT110), .A4(new_n833), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n759), .A2(new_n746), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n769), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n680), .A2(new_n711), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n671), .A2(new_n683), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n616), .A3(new_n701), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n723), .A2(new_n688), .A3(new_n749), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n687), .A2(new_n686), .B1(new_n746), .B2(new_n748), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .A3(new_n723), .A4(new_n842), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n568), .A2(new_n773), .A3(new_n505), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n629), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n641), .A2(new_n473), .A3(new_n619), .A4(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(new_n677), .A3(new_n742), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n617), .A3(new_n727), .A4(new_n734), .ZN(new_n853));
  INV_X1    g667(.A(new_n731), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n766), .A2(new_n839), .A3(new_n848), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  INV_X1    g673(.A(new_n734), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n677), .A3(new_n742), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n617), .A3(new_n727), .A4(new_n731), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n769), .A2(new_n837), .A3(new_n838), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n766), .A4(new_n848), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n848), .B2(KEYINPUT111), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n856), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n856), .A2(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n858), .A2(new_n866), .A3(KEYINPUT112), .A4(new_n859), .ZN(new_n874));
  INV_X1    g688(.A(new_n784), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n779), .B2(new_n781), .ZN(new_n876));
  INV_X1    g690(.A(new_n570), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n752), .A2(new_n726), .A3(new_n754), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n764), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n878), .A2(new_n764), .A3(new_n880), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT48), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n876), .A2(new_n877), .A3(new_n739), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n748), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n256), .A2(new_n570), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n705), .A2(new_n879), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n518), .A3(new_n628), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n569), .B(KEYINPUT117), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n518), .A2(new_n628), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n876), .A2(new_n877), .A3(new_n879), .A4(new_n745), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n878), .A2(new_n880), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT116), .B(new_n897), .C1(new_n901), .C2(new_n745), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n747), .A2(new_n371), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n903), .A2(KEYINPUT114), .A3(new_n710), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT114), .B1(new_n903), .B2(new_n710), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n785), .A2(new_n570), .A3(new_n740), .ZN(new_n907));
  OAI211_X1 g721(.A(KEYINPUT115), .B(KEYINPUT50), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n904), .A2(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n910));
  OR2_X1    g724(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n909), .A2(new_n887), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n900), .A2(new_n902), .A3(new_n908), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n822), .A2(new_n578), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n806), .A2(new_n808), .B1(KEYINPUT108), .B2(KEYINPUT47), .ZN(new_n915));
  INV_X1    g729(.A(new_n809), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n814), .A2(new_n815), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n907), .A2(new_n801), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT51), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n894), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n899), .B1(new_n890), .B2(new_n896), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n923), .A2(new_n912), .A3(new_n908), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n914), .B(KEYINPUT113), .Z(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n817), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT51), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n869), .A2(new_n873), .A3(new_n874), .A4(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT119), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(G952), .A2(G953), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n828), .B1(new_n931), .B2(new_n934), .ZN(G75));
  NOR2_X1   g749(.A1(new_n194), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n858), .A2(new_n866), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n519), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n373), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n426), .A2(new_n439), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n437), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(KEYINPUT56), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n939), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n947), .A3(new_n374), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT121), .B1(new_n939), .B2(new_n373), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n945), .B1(new_n951), .B2(new_n943), .ZN(G51));
  XOR2_X1   g766(.A(new_n795), .B(KEYINPUT57), .Z(new_n953));
  INV_X1    g767(.A(new_n867), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n859), .B1(new_n858), .B2(new_n866), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n613), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n939), .A2(new_n794), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n936), .B1(new_n957), .B2(new_n958), .ZN(G54));
  AND2_X1   g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n946), .A2(new_n513), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n513), .B1(new_n946), .B2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n936), .ZN(G60));
  NAND3_X1  g777(.A1(new_n869), .A2(new_n873), .A3(new_n874), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n624), .A2(new_n625), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT59), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n954), .B2(new_n955), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n625), .A3(new_n624), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n936), .B1(new_n968), .B2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n938), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n255), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n936), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n669), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n975), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n977), .B(KEYINPUT61), .C1(new_n978), .C2(new_n975), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  AOI21_X1  g797(.A(new_n428), .B1(new_n572), .B2(new_n427), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT123), .Z(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n855), .B2(new_n195), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n941), .B1(G898), .B2(new_n194), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  INV_X1    g802(.A(G227), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n195), .B1(new_n989), .B2(new_n682), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n288), .A2(new_n306), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(new_n508), .Z(new_n993));
  AND2_X1   g807(.A1(new_n846), .A2(new_n723), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n714), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  INV_X1    g810(.A(new_n370), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n802), .A2(new_n616), .A3(new_n690), .A4(new_n850), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n819), .B(new_n804), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n993), .B1(new_n1000), .B2(new_n195), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n804), .A2(new_n994), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT125), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n800), .A2(new_n690), .A3(new_n840), .A4(new_n764), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n819), .A2(new_n766), .A3(new_n769), .A4(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n194), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n194), .A2(G900), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n993), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n991), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n991), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1012), .B(new_n1001), .C1(new_n1013), .C2(new_n993), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1014), .ZN(G72));
  NOR3_X1   g829(.A1(new_n996), .A2(new_n863), .A3(new_n999), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n695), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n937), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n694), .A2(new_n330), .ZN(new_n1022));
  OR3_X1    g836(.A1(new_n1004), .A2(new_n863), .A3(new_n1006), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n871), .A2(new_n872), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n323), .A2(KEYINPUT126), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(new_n362), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n1018), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT127), .Z(new_n1029));
  NOR2_X1   g843(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1021), .A2(new_n1024), .A3(new_n1030), .ZN(G57));
endmodule


