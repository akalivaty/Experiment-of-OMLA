//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT28), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n209), .B2(KEYINPUT26), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n206), .B(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT66), .B(KEYINPUT26), .Z(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n204), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n205), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n207), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n206), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(G183gat), .B(G190gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(new_n220), .ZN(new_n223));
  AOI211_X1 g022(.A(new_n218), .B(new_n219), .C1(new_n223), .C2(KEYINPUT64), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT25), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n212), .A2(new_n217), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  NOR4_X1   g027(.A1(new_n227), .A2(new_n228), .A3(new_n223), .A4(new_n219), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n216), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT29), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G226gat), .ZN(new_n233));
  INV_X1    g032(.A(G233gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G197gat), .B(G204gat), .ZN(new_n239));
  INV_X1    g038(.A(G211gat), .ZN(new_n240));
  INV_X1    g039(.A(G218gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(KEYINPUT22), .B2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G211gat), .B(G218gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n248), .A3(new_n236), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n230), .B2(new_n236), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n235), .B(new_n245), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G8gat), .B(G36gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G64gat), .B(G92gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OR3_X1    g056(.A1(new_n253), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n247), .A2(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n257), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT30), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G113gat), .B(G120gat), .Z(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n273));
  INV_X1    g072(.A(G148gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G141gat), .ZN(new_n275));
  INV_X1    g074(.A(G141gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(G148gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  OR2_X1    g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(KEYINPUT2), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT70), .B1(new_n274), .B2(G141gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n276), .B2(G148gat), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n274), .A2(KEYINPUT70), .A3(G141gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT72), .B(KEYINPUT3), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n287), .A2(new_n270), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT4), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(KEYINPUT73), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n294), .B(new_n296), .C1(KEYINPUT4), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n295), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n272), .A2(new_n287), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n293), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n299), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT4), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT75), .B1(new_n295), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n297), .B2(new_n307), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n301), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n299), .A4(new_n294), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(G1gat), .B(G29gat), .Z(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT6), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n306), .A2(new_n317), .A3(new_n311), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n312), .A2(KEYINPUT6), .A3(new_n318), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n258), .A2(new_n262), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n230), .A2(new_n270), .ZN(new_n325));
  INV_X1    g124(.A(new_n270), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n326), .B(new_n216), .C1(new_n226), .C2(new_n229), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G227gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(new_n234), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT32), .ZN(new_n334));
  XNOR2_X1  g133(.A(G15gat), .B(G43gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G71gat), .B(G99gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n337), .B1(new_n333), .B2(KEYINPUT32), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT67), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT33), .B1(new_n328), .B2(new_n330), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n337), .ZN(new_n346));
  INV_X1    g145(.A(new_n330), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n325), .B2(new_n327), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT67), .B1(new_n350), .B2(new_n343), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n340), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT34), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g153(.A(KEYINPUT34), .B(new_n340), .C1(new_n345), .C2(new_n351), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n332), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n340), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n342), .B1(new_n341), .B2(new_n344), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n350), .A2(KEYINPUT67), .A3(new_n343), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT34), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n352), .A2(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n331), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n245), .B1(new_n290), .B2(new_n231), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n287), .A2(new_n245), .A3(new_n231), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(new_n291), .A3(G228gat), .A4(G233gat), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n288), .B2(new_n289), .ZN(new_n368));
  INV_X1    g167(.A(G228gat), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n364), .A2(new_n368), .B1(new_n369), .B2(new_n234), .ZN(new_n370));
  INV_X1    g169(.A(G22gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n374));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375));
  INV_X1    g174(.A(G50gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n367), .A2(new_n370), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G22gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n374), .A2(new_n380), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n380), .B1(new_n382), .B2(new_n372), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n372), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT77), .A3(new_n379), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n324), .A2(new_n356), .A3(new_n363), .A4(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n390), .A2(KEYINPUT35), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(KEYINPUT35), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n324), .A2(new_n389), .ZN(new_n393));
  INV_X1    g192(.A(new_n389), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n309), .A2(new_n292), .A3(new_n310), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT39), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n304), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n317), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT40), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT39), .B1(new_n303), .B2(new_n304), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n395), .B2(new_n304), .ZN(new_n401));
  OR3_X1    g200(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n398), .B2(new_n401), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n402), .A2(new_n319), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n262), .A2(new_n258), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n394), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n322), .A2(new_n323), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT37), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n256), .B1(new_n259), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n410), .B2(new_n259), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT38), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n238), .B2(new_n245), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n235), .B1(new_n250), .B2(new_n251), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n245), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT38), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n418), .B(new_n411), .C1(new_n417), .C2(new_n416), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n409), .A2(new_n413), .A3(new_n260), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n393), .B1(new_n407), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n354), .A2(new_n355), .A3(new_n332), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n331), .B1(new_n361), .B2(new_n362), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n356), .A2(new_n363), .A3(KEYINPUT36), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n391), .A2(new_n392), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G113gat), .B(G141gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT80), .B(G197gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT11), .B(G169gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT12), .ZN(new_n434));
  INV_X1    g233(.A(G1gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT16), .ZN(new_n436));
  INV_X1    g235(.A(G15gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G22gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n371), .A2(G15gat), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(G1gat), .B1(new_n438), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g240(.A(G8gat), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n443));
  INV_X1    g242(.A(G8gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G22gat), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n443), .B(new_n444), .C1(G1gat), .C2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n442), .A2(KEYINPUT82), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT82), .B1(new_n442), .B2(new_n446), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G29gat), .ZN(new_n450));
  INV_X1    g249(.A(G36gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT14), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT14), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(G29gat), .B2(G36gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(G29gat), .A2(G36gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457));
  INV_X1    g256(.A(G43gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n376), .ZN(new_n459));
  NAND2_X1  g258(.A1(G43gat), .A2(G50gat), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n460), .ZN(new_n463));
  NOR2_X1   g262(.A1(G43gat), .A2(G50gat), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT15), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n457), .A3(new_n460), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n462), .B(KEYINPUT81), .C1(new_n467), .C2(new_n456), .ZN(new_n468));
  INV_X1    g267(.A(new_n456), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n465), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT17), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n449), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT83), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n442), .A2(new_n446), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n442), .A2(KEYINPUT84), .A3(new_n446), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n468), .A3(new_n471), .A4(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n476), .A2(KEYINPUT18), .A3(new_n479), .A4(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n483), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT84), .B1(new_n442), .B2(new_n446), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n472), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n484), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n478), .B(KEYINPUT13), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n476), .A2(new_n493), .A3(new_n479), .A4(new_n484), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n479), .A3(new_n484), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT18), .B1(new_n495), .B2(KEYINPUT85), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n434), .B(new_n492), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(KEYINPUT85), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT86), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n502), .A3(new_n494), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n491), .A3(KEYINPUT87), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n501), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n497), .B1(new_n507), .B2(new_n434), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n428), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G64gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(G57gat), .ZN(new_n511));
  INV_X1    g310(.A(G57gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(G64gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT9), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  OR2_X1    g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT88), .B1(new_n510), .B2(G57gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n512), .A3(G64gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n518), .B(new_n520), .C1(new_n512), .C2(G64gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n515), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G127gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n486), .A2(new_n487), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n525), .A2(new_n526), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n538));
  INV_X1    g337(.A(G155gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n537), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT89), .B1(G85gat), .B2(G92gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI211_X1 g347(.A(KEYINPUT89), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT90), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT90), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(G92gat), .ZN(new_n554));
  INV_X1    g353(.A(G85gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  INV_X1    g356(.A(G99gat), .ZN(new_n558));
  INV_X1    g357(.A(G106gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT8), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n557), .B1(new_n556), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n550), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n550), .B(new_n564), .C1(new_n561), .C2(new_n562), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n472), .ZN(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n568), .A2(new_n569), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n473), .A2(new_n475), .A3(new_n566), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G190gat), .B(G218gat), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n576), .B(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n544), .A2(new_n580), .A3(KEYINPUT92), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT92), .B1(new_n544), .B2(new_n580), .ZN(new_n582));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n525), .A3(new_n567), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n525), .A4(new_n567), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n517), .A2(new_n524), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n563), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n556), .A2(new_n560), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT91), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n601), .B2(new_n550), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT95), .B(KEYINPUT10), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n593), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n594), .A2(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n568), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n588), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n603), .B1(new_n591), .B2(new_n592), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n587), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n586), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI211_X1 g412(.A(new_n605), .B(new_n603), .C1(new_n591), .C2(new_n592), .ZN(new_n614));
  INV_X1    g413(.A(new_n609), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n587), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n585), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n618), .A3(KEYINPUT96), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT96), .B1(new_n613), .B2(new_n618), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n581), .A2(new_n582), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n509), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n408), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT97), .B(G1gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(G1324gat));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n406), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G8gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(KEYINPUT98), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(KEYINPUT42), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT16), .B(G8gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n635), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(G1325gat));
  AND3_X1   g437(.A1(new_n356), .A2(new_n363), .A3(KEYINPUT36), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT36), .B1(new_n356), .B2(new_n363), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT100), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n425), .A2(new_n642), .A3(new_n426), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G15gat), .B1(new_n624), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n423), .A2(new_n424), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n437), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n624), .B2(new_n647), .ZN(G1326gat));
  NOR3_X1   g447(.A1(new_n428), .A2(new_n389), .A3(new_n508), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n623), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NAND3_X1  g451(.A1(new_n641), .A2(new_n421), .A3(new_n643), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n391), .A2(new_n392), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657));
  INV_X1    g456(.A(new_n580), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT44), .B1(new_n428), .B2(new_n580), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n580), .B1(new_n653), .B2(new_n654), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n656), .B1(new_n662), .B2(new_n657), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n622), .A2(new_n508), .A3(new_n544), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G29gat), .B1(new_n667), .B2(new_n408), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n428), .A2(new_n580), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n665), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(G29gat), .A3(new_n408), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT45), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(G1328gat));
  OAI21_X1  g472(.A(G36gat), .B1(new_n667), .B2(new_n405), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n670), .A2(G36gat), .A3(new_n405), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT46), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(G1329gat));
  INV_X1    g476(.A(new_n646), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n670), .A2(G43gat), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n644), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n680), .A3(new_n666), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n681), .B2(G43gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g482(.A(new_n394), .B(new_n666), .C1(new_n661), .C2(new_n663), .ZN(new_n684));
  NOR4_X1   g483(.A1(new_n622), .A2(G50gat), .A3(new_n544), .A4(new_n580), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n684), .A2(G50gat), .B1(new_n649), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n581), .A2(new_n582), .ZN(new_n688));
  AND4_X1   g487(.A1(new_n508), .A2(new_n655), .A3(new_n688), .A4(new_n622), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n409), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g490(.A(new_n405), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT103), .Z(new_n694));
  NOR2_X1   g493(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1333gat));
  NAND2_X1  g495(.A1(new_n689), .A2(new_n680), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n678), .A2(G71gat), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n697), .A2(G71gat), .B1(new_n689), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g499(.A1(new_n689), .A2(new_n394), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  INV_X1    g501(.A(new_n508), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n621), .A2(new_n703), .A3(new_n544), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n409), .B(new_n704), .C1(new_n661), .C2(new_n663), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G85gat), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n703), .A2(new_n544), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n662), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n662), .A2(KEYINPUT51), .A3(new_n707), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n713), .A3(new_n709), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n622), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n409), .A2(new_n555), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n706), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1336gat));
  INV_X1    g518(.A(new_n715), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n405), .A2(G92gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n664), .A2(new_n406), .A3(new_n704), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n552), .A2(new_n554), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n711), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n622), .A3(new_n721), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(new_n726), .ZN(G1337gat));
  AOI21_X1  g530(.A(G99gat), .B1(new_n720), .B2(new_n646), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n664), .A2(new_n704), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n644), .A2(new_n558), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(G1338gat));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n394), .B(new_n704), .C1(new_n661), .C2(new_n663), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G106gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n389), .A2(new_n621), .A3(G106gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n712), .A2(new_n714), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n728), .A2(new_n740), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n736), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n737), .A2(G106gat), .B1(new_n728), .B2(new_n740), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n746), .B(KEYINPUT106), .C1(new_n739), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1339gat));
  NAND3_X1  g548(.A1(new_n688), .A2(new_n508), .A3(new_n621), .ZN(new_n750));
  INV_X1    g549(.A(new_n544), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n609), .A2(new_n588), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n607), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n616), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n585), .B1(new_n610), .B2(new_n753), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n610), .A2(new_n612), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n585), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT54), .B1(new_n614), .B2(new_n754), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n610), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n753), .B(new_n587), .C1(new_n614), .C2(new_n615), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n586), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n752), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n489), .A2(new_n490), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n479), .B1(new_n476), .B2(new_n484), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n433), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n497), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n658), .A2(new_n760), .A3(new_n765), .A4(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n434), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n505), .A2(new_n506), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n502), .B1(new_n496), .B2(new_n494), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n776), .B2(new_n503), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n765), .B(new_n760), .C1(new_n777), .C2(new_n497), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n770), .B1(new_n619), .B2(new_n620), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n658), .B1(new_n780), .B2(KEYINPUT107), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n772), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n751), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g585(.A(KEYINPUT108), .B(new_n772), .C1(new_n781), .C2(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n750), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n678), .A2(new_n394), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n409), .A3(new_n405), .ZN(new_n791));
  INV_X1    g590(.A(G113gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n792), .A3(new_n508), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n409), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT109), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n796), .A3(new_n409), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n405), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n703), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n793), .B1(new_n800), .B2(new_n792), .ZN(G1340gat));
  INV_X1    g600(.A(G120gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n791), .A2(new_n802), .A3(new_n621), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n622), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n802), .ZN(G1341gat));
  NOR2_X1   g604(.A1(new_n751), .A2(G127gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n795), .A2(new_n405), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G127gat), .B1(new_n791), .B2(new_n751), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n809), .B(KEYINPUT110), .Z(G1342gat));
  INV_X1    g609(.A(G134gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n406), .A2(new_n580), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n798), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT56), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n815), .A3(new_n811), .A4(new_n812), .ZN(new_n816));
  INV_X1    g615(.A(new_n812), .ZN(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n794), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(G1343gat));
  NAND4_X1  g618(.A1(new_n641), .A2(new_n643), .A3(new_n409), .A4(new_n405), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT111), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n788), .B2(new_n394), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n394), .A2(KEYINPUT57), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT55), .B1(new_n761), .B2(new_n610), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n618), .B1(new_n824), .B2(new_n764), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n616), .A2(new_n756), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n758), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n508), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n497), .A2(new_n769), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n613), .A2(new_n618), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT96), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n613), .A2(new_n618), .A3(KEYINPUT96), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n580), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n544), .B1(new_n835), .B2(new_n771), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n750), .B1(new_n836), .B2(KEYINPUT112), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n658), .B1(new_n778), .B2(new_n779), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT112), .B(new_n751), .C1(new_n838), .C2(new_n772), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n823), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT113), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n843), .B(new_n823), .C1(new_n837), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n703), .B(new_n821), .C1(new_n822), .C2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n276), .B1(new_n846), .B2(KEYINPUT116), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(KEYINPUT116), .B2(new_n846), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n788), .A2(new_n394), .ZN(new_n850));
  INV_X1    g649(.A(new_n820), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n703), .A2(new_n276), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT115), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n848), .B(new_n849), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n852), .A2(new_n854), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n821), .B1(new_n822), .B2(new_n845), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT114), .B(new_n821), .C1(new_n822), .C2(new_n845), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n703), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n856), .B1(new_n861), .B2(G141gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n855), .B1(new_n849), .B2(new_n862), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n788), .A2(new_n823), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n751), .B1(new_n838), .B2(new_n772), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n389), .B1(new_n750), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT118), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n867), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n864), .A2(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n788), .A2(KEYINPUT117), .A3(new_n823), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(new_n622), .A3(new_n821), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT59), .B1(new_n873), .B2(new_n274), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n622), .A3(new_n860), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(G148gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n850), .A2(new_n274), .A3(new_n622), .A4(new_n851), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1345gat));
  AND3_X1   g679(.A1(new_n859), .A2(new_n544), .A3(new_n860), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n544), .A2(new_n539), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n881), .A2(new_n539), .B1(new_n852), .B2(new_n882), .ZN(G1346gat));
  NAND3_X1  g682(.A1(new_n859), .A2(new_n658), .A3(new_n860), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G162gat), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n817), .A2(G162gat), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n850), .A2(new_n409), .A3(new_n644), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT119), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n409), .A2(new_n405), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n790), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n703), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(G169gat), .ZN(G1348gat));
  NOR2_X1   g696(.A1(new_n894), .A2(new_n621), .ZN(new_n898));
  XNOR2_X1  g697(.A(KEYINPUT120), .B(G176gat), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n898), .B(new_n899), .ZN(G1349gat));
  AOI21_X1  g699(.A(new_n202), .B1(KEYINPUT121), .B2(G183gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n544), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(G183gat), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n894), .A2(new_n751), .B1(KEYINPUT121), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(G1350gat));
  NAND4_X1  g709(.A1(new_n788), .A2(new_n789), .A3(new_n658), .A4(new_n893), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G190gat), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(KEYINPUT124), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(KEYINPUT124), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n915), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n911), .A2(G190gat), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n917), .A2(KEYINPUT125), .A3(new_n918), .A4(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n918), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n925), .ZN(G1351gat));
  NAND3_X1  g725(.A1(new_n644), .A2(new_n406), .A3(new_n394), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(new_n409), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(new_n788), .ZN(new_n931));
  AOI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n703), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n644), .A2(new_n893), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n872), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n703), .A2(G197gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n621), .A2(G204gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n938));
  OR2_X1    g737(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n931), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(new_n934), .B2(new_n622), .ZN(new_n942));
  AND4_X1   g741(.A1(new_n788), .A2(new_n930), .A3(new_n938), .A4(new_n937), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n931), .A2(new_n240), .A3(new_n544), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n872), .A2(new_n544), .A3(new_n933), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n241), .A3(new_n658), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n934), .A2(new_n658), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n241), .ZN(G1355gat));
endmodule


