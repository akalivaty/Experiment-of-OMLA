//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT65), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n465), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n477), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n476), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n477), .C1(new_n462), .C2(new_n463), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n464), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n488), .A2(G2105), .B1(G102), .B2(new_n467), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  INV_X1    g066(.A(G651), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT6), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G651), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n493), .A2(new_n495), .A3(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G50), .ZN(new_n497));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n493), .A2(new_n495), .A3(new_n500), .A4(new_n502), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT66), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n509), .A2(new_n510), .A3(new_n493), .A4(new_n495), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n497), .B(new_n506), .C1(new_n512), .C2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n518), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n493), .A2(new_n495), .A3(G51), .A4(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n500), .A2(new_n502), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n509), .A2(KEYINPUT67), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n508), .A2(G89), .A3(new_n511), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G168));
  NAND3_X1  g106(.A1(new_n508), .A2(G90), .A3(new_n511), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n503), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n496), .A2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n508), .A2(G81), .A3(new_n511), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n500), .A2(new_n502), .A3(G56), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G651), .B1(new_n496), .B2(G43), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n540), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n541), .A2(new_n545), .A3(new_n540), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND4_X1  g130(.A1(new_n493), .A2(new_n495), .A3(G53), .A4(G543), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n508), .A2(G91), .A3(new_n511), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT69), .B(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n503), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n508), .A2(G89), .A3(new_n511), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n526), .A2(new_n527), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n520), .A2(new_n521), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n564), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n528), .A2(KEYINPUT70), .A3(new_n529), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G286));
  AND2_X1   g146(.A1(new_n508), .A2(new_n511), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G87), .ZN(new_n573));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n492), .B1(new_n503), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(G49), .B2(new_n496), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n572), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n496), .A2(G48), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n503), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n580), .B1(new_n583), .B2(G651), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n583), .A2(new_n580), .A3(G651), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n578), .B(new_n579), .C1(new_n584), .C2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n492), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT72), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(new_n496), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n589), .B1(new_n590), .B2(new_n591), .C1(new_n592), .C2(new_n512), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G171), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n508), .A2(G92), .A3(new_n511), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(KEYINPUT75), .A2(G66), .ZN(new_n601));
  NAND2_X1  g176(.A1(KEYINPUT75), .A2(G66), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n601), .A2(new_n500), .A3(new_n502), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT76), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(G651), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n496), .A2(G54), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n508), .A2(G92), .A3(new_n511), .A4(new_n598), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n600), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n596), .B1(new_n613), .B2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT73), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT73), .B2(new_n595), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(KEYINPUT73), .B2(new_n595), .ZN(G321));
  NAND2_X1  g192(.A1(G299), .A2(new_n594), .ZN(new_n618));
  INV_X1    g193(.A(G286), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n594), .ZN(G280));
  XNOR2_X1  g195(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n613), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND3_X1  g198(.A1(new_n547), .A2(new_n594), .A3(new_n548), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n612), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n594), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g202(.A(new_n464), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n467), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n477), .A2(G111), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n466), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .C1(G99), .C2(G2105), .ZN(new_n636));
  AOI22_X1  g211(.A1(G123), .A2(new_n478), .B1(new_n465), .B2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n639), .ZN(G156));
  INV_X1    g215(.A(G14), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  INV_X1    g221(.A(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OAI21_X1  g224(.A(KEYINPUT14), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT80), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n654), .A2(new_n655), .A3(new_n645), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n644), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n643), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1341), .B(G1348), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n642), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g240(.A1(new_n659), .A2(new_n661), .A3(KEYINPUT81), .A4(new_n663), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n641), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n664), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n687), .B1(KEYINPUT20), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(KEYINPUT20), .C2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT82), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  AOI22_X1  g274(.A1(G119), .A2(new_n478), .B1(new_n465), .B2(G131), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n466), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI221_X1 g278(.A(new_n703), .B1(new_n702), .B2(new_n701), .C1(G107), .C2(new_n477), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT33), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1976), .ZN(new_n714));
  NOR2_X1   g289(.A1(G166), .A2(new_n709), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n709), .B2(G22), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(G6), .ZN(new_n719));
  INV_X1    g294(.A(G305), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n709), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT32), .B(G1981), .ZN(new_n722));
  OAI22_X1  g297(.A1(new_n717), .A2(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n714), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n708), .B1(new_n725), .B2(KEYINPUT34), .ZN(new_n726));
  INV_X1    g301(.A(G24), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT84), .B1(new_n727), .B2(G16), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n727), .A2(KEYINPUT84), .A3(G16), .ZN(new_n729));
  INV_X1    g304(.A(G290), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n709), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT85), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1986), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n726), .B(new_n733), .C1(KEYINPUT34), .C2(new_n725), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G168), .A2(new_n709), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n709), .B2(G21), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n734), .A2(new_n735), .ZN(new_n741));
  INV_X1    g316(.A(G28), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n742), .A2(KEYINPUT89), .A3(KEYINPUT30), .ZN(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT89), .B1(new_n742), .B2(KEYINPUT30), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n477), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G139), .B2(new_n465), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n467), .A2(G103), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n744), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n744), .B2(G33), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n747), .B1(new_n744), .B2(new_n638), .C1(new_n757), .C2(G2072), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT31), .B(G11), .Z(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n744), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n465), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n478), .A2(G128), .ZN(new_n764));
  NOR2_X1   g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(new_n477), .B2(G116), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  NOR2_X1   g344(.A1(G5), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G171), .B2(G16), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(G1961), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n758), .A2(new_n759), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G32), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n465), .A2(G141), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n478), .A2(G129), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n467), .A2(G105), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT26), .Z(new_n781));
  NAND4_X1  g356(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT27), .B(G1996), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n709), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n613), .B2(new_n709), .ZN(new_n788));
  INV_X1    g363(.A(G1348), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n744), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n744), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT92), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT91), .B(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G2072), .B2(new_n757), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n775), .A2(new_n786), .A3(new_n790), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n798), .A2(new_n744), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G160), .B2(new_n744), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G2084), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT88), .ZN(new_n803));
  INV_X1    g378(.A(G299), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT23), .B1(new_n804), .B2(new_n709), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n709), .A2(G20), .ZN(new_n806));
  MUX2_X1   g381(.A(KEYINPUT23), .B(new_n805), .S(new_n806), .Z(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G1956), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(G1956), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G19), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n549), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  NAND4_X1  g387(.A1(new_n803), .A2(new_n808), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n801), .A2(G2084), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT90), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n738), .A2(new_n739), .ZN(new_n816));
  INV_X1    g391(.A(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT93), .B1(new_n817), .B2(G29), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n817), .A2(KEYINPUT93), .A3(G29), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n818), .B(new_n819), .C1(G162), .C2(new_n744), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT29), .Z(new_n821));
  INV_X1    g396(.A(G2090), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n815), .B(new_n823), .C1(new_n822), .C2(new_n821), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n797), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n736), .A2(new_n740), .A3(new_n741), .A4(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NAND3_X1  g402(.A1(new_n500), .A2(new_n502), .A3(G67), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(KEYINPUT94), .A3(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(G651), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n496), .A2(G55), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n508), .A2(G93), .A3(new_n511), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n612), .A2(new_n622), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n541), .A2(new_n545), .ZN(new_n844));
  AND4_X1   g419(.A1(new_n844), .A2(new_n835), .A3(new_n836), .A4(new_n834), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n549), .B2(new_n837), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n843), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n840), .B1(new_n847), .B2(G860), .ZN(G145));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n767), .B(new_n782), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(new_n490), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n490), .ZN(new_n852));
  INV_X1    g427(.A(new_n754), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n477), .A2(G118), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n466), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n859), .B1(new_n858), .B2(new_n857), .C1(G106), .C2(G2105), .ZN(new_n860));
  AOI22_X1  g435(.A1(G130), .A2(new_n478), .B1(new_n465), .B2(G142), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n630), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n705), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n856), .A2(KEYINPUT97), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n854), .A2(new_n864), .A3(new_n855), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n474), .B(new_n638), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G162), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n869), .B(new_n871), .C1(new_n864), .C2(new_n856), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n865), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n865), .B2(new_n868), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n856), .A2(new_n864), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n849), .B(new_n872), .C1(new_n877), .C2(new_n871), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(new_n548), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n837), .B1(new_n880), .B2(new_n546), .ZN(new_n881));
  INV_X1    g456(.A(new_n837), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n844), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n625), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n600), .A2(new_n611), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n607), .B1(new_n603), .B2(new_n604), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n889), .A2(G651), .B1(G54), .B2(new_n496), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(G299), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n612), .A2(new_n804), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  AOI21_X1  g470(.A(G299), .B1(new_n886), .B2(new_n890), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n612), .A2(new_n804), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n892), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n894), .B1(new_n901), .B2(new_n885), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT42), .Z(new_n903));
  XNOR2_X1  g478(.A(G288), .B(G303), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G305), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(G305), .ZN(new_n907));
  OAI21_X1  g482(.A(G290), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n730), .A3(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n903), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(G868), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(G868), .B2(new_n882), .ZN(new_n916));
  MUX2_X1   g491(.A(new_n915), .B(new_n916), .S(KEYINPUT99), .Z(G295));
  MUX2_X1   g492(.A(new_n915), .B(new_n916), .S(KEYINPUT99), .Z(G331));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n919));
  NAND3_X1  g494(.A1(G301), .A2(new_n529), .A3(new_n528), .ZN(new_n920));
  AOI22_X1  g495(.A1(G286), .A2(G171), .B1(new_n920), .B2(KEYINPUT100), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n922));
  AOI211_X1 g497(.A(new_n922), .B(G301), .C1(new_n569), .C2(new_n570), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n884), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND4_X1   g499(.A1(KEYINPUT70), .A2(new_n529), .A3(new_n566), .A4(new_n567), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT70), .B1(new_n528), .B2(new_n529), .ZN(new_n926));
  OAI21_X1  g501(.A(G171), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n920), .A2(KEYINPUT100), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(G286), .A2(KEYINPUT100), .A3(G171), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n846), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI221_X4 g506(.A(new_n919), .B1(new_n898), .B2(new_n899), .C1(new_n924), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n931), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT101), .B1(new_n933), .B2(new_n900), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n924), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n846), .A2(new_n929), .A3(KEYINPUT102), .A4(new_n930), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n893), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n911), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT103), .B1(new_n941), .B2(G37), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n900), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n919), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n933), .A2(KEYINPUT101), .A3(new_n900), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n940), .A2(new_n944), .A3(new_n911), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT104), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n935), .A2(new_n948), .A3(new_n911), .A4(new_n940), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n951));
  INV_X1    g526(.A(new_n893), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n937), .B2(new_n938), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n953), .A2(new_n932), .A3(new_n934), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n951), .B(new_n849), .C1(new_n954), .C2(new_n911), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n942), .A2(new_n950), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n939), .A2(new_n901), .B1(new_n952), .B2(new_n933), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n912), .ZN(new_n960));
  AND4_X1   g535(.A1(KEYINPUT43), .A2(new_n950), .A3(new_n849), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n956), .A2(new_n963), .A3(KEYINPUT43), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n950), .A2(new_n957), .A3(new_n849), .A4(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n962), .B1(new_n968), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n490), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT106), .ZN(new_n974));
  INV_X1    g549(.A(G2067), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n767), .B(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT107), .Z(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(new_n974), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n974), .A2(new_n783), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n973), .A2(G1996), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n783), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n707), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n700), .A4(new_n704), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n767), .A2(G2067), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n974), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n705), .B(new_n985), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n974), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n973), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT48), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n983), .A2(KEYINPUT46), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n983), .A2(KEYINPUT46), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n978), .A2(new_n980), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  NOR3_X1   g573(.A1(new_n988), .A2(new_n994), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT63), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n1001), .B(G1384), .C1(new_n485), .C2(new_n489), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n971), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n972), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n717), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT50), .B1(new_n490), .B2(new_n970), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(G1384), .C1(new_n485), .C2(new_n489), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n972), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(G2090), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(KEYINPUT109), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1014), .B(new_n1015), .C1(new_n1012), .C2(new_n1011), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT110), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n972), .A2(new_n970), .A3(new_n490), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n573), .A2(new_n1022), .A3(G1976), .A4(new_n576), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1020), .A2(G8), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n711), .A2(G1976), .ZN(new_n1025));
  OR3_X1    g600(.A1(new_n1024), .A2(KEYINPUT52), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G305), .A2(G1981), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n585), .A2(new_n584), .ZN(new_n1028));
  INV_X1    g603(.A(G1981), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n579), .A4(new_n578), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1021), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1024), .B2(KEYINPUT52), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1024), .A2(new_n1039), .A3(KEYINPUT52), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1026), .B(new_n1038), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1016), .B1(new_n1010), .B2(G8), .ZN(new_n1043));
  OR3_X1    g618(.A1(new_n1018), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1004), .A2(new_n739), .ZN(new_n1045));
  INV_X1    g620(.A(new_n972), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n490), .A2(new_n970), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1007), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n490), .A2(KEYINPUT50), .A3(new_n970), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G2084), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(KEYINPUT114), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1009), .B2(G2084), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1045), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(G8), .A3(new_n619), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1000), .B1(new_n1044), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1040), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1024), .A2(new_n1039), .A3(KEYINPUT52), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1026), .A4(new_n1038), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1058), .A2(new_n1063), .A3(KEYINPUT63), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1018), .A2(new_n1043), .A3(new_n1056), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT115), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(new_n1063), .A3(KEYINPUT63), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1043), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1055), .A2(G8), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n619), .A3(new_n1017), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1067), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1057), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1058), .A2(new_n1063), .A3(new_n1018), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1038), .A2(new_n1019), .A3(new_n711), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1030), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1036), .B(KEYINPUT113), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1073), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1055), .A2(KEYINPUT123), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1045), .A2(new_n1052), .A3(new_n1054), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G168), .A2(new_n1035), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n530), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1089), .A2(KEYINPUT124), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(KEYINPUT124), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1087), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1069), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1080), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1084), .A2(G168), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1092), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g674(.A(KEYINPUT62), .B1(new_n1069), .B2(new_n1094), .C1(new_n1099), .C2(new_n1087), .ZN(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1003), .A2(new_n1101), .A3(new_n972), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1102), .A2(new_n1103), .B1(G1961), .B2(new_n1050), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1103), .A2(KEYINPUT125), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(KEYINPUT125), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT126), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1102), .A2(new_n1109), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1104), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G301), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1096), .A2(new_n1100), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n971), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1002), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n972), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1003), .A2(KEYINPUT119), .A3(new_n972), .A4(new_n1116), .ZN(new_n1120));
  INV_X1    g695(.A(G1956), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1009), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n558), .A2(new_n1124), .A3(new_n562), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n558), .B2(new_n562), .ZN(new_n1126));
  INV_X1    g701(.A(new_n557), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT117), .B1(new_n1128), .B2(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n804), .A2(KEYINPUT57), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1126), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n558), .A2(new_n1124), .A3(new_n562), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n557), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT118), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1129), .A2(new_n1136), .A3(new_n1139), .A4(new_n1130), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1141), .A2(KEYINPUT120), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(KEYINPUT120), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1123), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1009), .A2(new_n789), .B1(new_n975), .B2(new_n1034), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1141), .A2(new_n1122), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n613), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1123), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1150), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1123), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1149), .B(new_n1152), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT58), .B(G1341), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1004), .A2(G1996), .B1(new_n1034), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n549), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT59), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1145), .A2(KEYINPUT60), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n612), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n613), .A2(KEYINPUT122), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n612), .A2(new_n1164), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(new_n1168), .C1(KEYINPUT60), .C2(new_n1145), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1155), .A2(new_n1152), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1144), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1148), .B1(new_n1158), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n1111), .B2(G301), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1111), .A2(G301), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT54), .B(new_n1174), .C1(new_n1176), .C2(new_n1112), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1111), .A2(G301), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1178), .B(new_n1175), .C1(KEYINPUT127), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1113), .B1(new_n1173), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1044), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1079), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(G290), .A2(G1986), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n973), .B1(new_n991), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n990), .A2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT108), .Z(new_n1190));
  OAI21_X1  g765(.A(new_n999), .B1(new_n1186), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g766(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1193), .A2(KEYINPUT105), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n956), .A2(new_n963), .A3(KEYINPUT43), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1194), .A2(new_n966), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G229), .A2(new_n460), .ZN(new_n1197));
  AOI21_X1  g771(.A(G227), .B1(new_n667), .B2(new_n668), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n878), .A2(new_n1198), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(G308));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n1199), .A3(new_n1197), .ZN(G225));
endmodule


