//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(new_n461), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n461), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n464), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT66), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n477), .B(new_n480), .C1(new_n485), .C2(G136), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n487), .A3(G138), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n461), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(G126), .B2(new_n475), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AND3_X1   g081(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT6), .B1(KEYINPUT67), .B2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(new_n501), .B2(new_n502), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT67), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT68), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n509), .ZN(new_n529));
  OAI21_X1  g104(.A(G543), .B1(new_n507), .B2(new_n508), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT69), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n515), .A2(new_n516), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(new_n533), .A3(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n529), .B1(G51), .B2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n535), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n510), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  OAI21_X1  g115(.A(G64), .B1(new_n501), .B2(new_n502), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(G651), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  AOI211_X1 g120(.A(KEYINPUT70), .B(new_n545), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n539), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(new_n535), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n503), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(G651), .A2(new_n552), .B1(new_n510), .B2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT71), .Z(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n509), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n532), .A2(new_n526), .A3(KEYINPUT72), .A4(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n530), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n517), .A2(new_n569), .A3(G53), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n503), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n566), .A2(new_n571), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(new_n539), .B2(new_n547), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n535), .A2(G52), .B1(G90), .B2(new_n510), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n579), .B(KEYINPUT73), .C1(new_n544), .C2(new_n546), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G301));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n535), .A2(G51), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n529), .ZN(new_n584));
  NAND2_X1  g159(.A1(G168), .A2(KEYINPUT74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  NAND2_X1  g163(.A1(new_n517), .A2(G49), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n509), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n503), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n510), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n517), .A2(G48), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  AND2_X1   g174(.A1(new_n535), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n601), .A2(new_n545), .B1(new_n602), .B2(new_n509), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  AOI21_X1  g180(.A(new_n533), .B1(new_n532), .B2(G543), .ZN(new_n606));
  AOI211_X1 g181(.A(KEYINPUT69), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n607));
  OAI21_X1  g182(.A(G54), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n509), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n532), .A2(new_n526), .A3(KEYINPUT10), .A4(G92), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n503), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G651), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n608), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n618), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g194(.A(new_n618), .B(G301), .S(G868), .Z(G321));
  NOR2_X1   g195(.A1(G299), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n586), .B2(G868), .ZN(G297));
  AOI21_X1  g197(.A(new_n621), .B1(new_n586), .B2(G868), .ZN(G280));
  AND3_X1   g198(.A1(new_n608), .A2(new_n613), .A3(new_n617), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT75), .B(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(G860), .B2(new_n625), .ZN(G148));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n475), .A2(G123), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n461), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n482), .A2(new_n484), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n631), .B1(new_n632), .B2(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(G2100), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT77), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT78), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n643), .A3(new_n645), .ZN(G156));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT80), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT81), .Z(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(KEYINPUT83), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  NOR3_X1   g262(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n687), .B2(new_n690), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n687), .A2(new_n690), .ZN(new_n698));
  INV_X1    g273(.A(new_n691), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n697), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n696), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n697), .A3(new_n692), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(G229));
  XOR2_X1   g283(.A(KEYINPUT84), .B(G29), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G35), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT29), .Z(new_n713));
  INV_X1    g288(.A(G2090), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n710), .A2(G27), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G164), .B2(new_n710), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2078), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT99), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n715), .B(new_n721), .C1(KEYINPUT99), .C2(new_n719), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n709), .A2(G26), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n485), .A2(G140), .ZN(new_n725));
  NOR2_X1   g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT89), .Z(new_n727));
  INV_X1    g302(.A(G116), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n472), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(new_n729), .B1(G128), .B2(new_n475), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n724), .B1(new_n731), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(G2067), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(G33), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI22_X1  g313(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n738), .B1(new_n461), .B2(new_n739), .C1(new_n634), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n736), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT24), .B(G34), .ZN(new_n745));
  AOI22_X1  g320(.A1(G160), .A2(G29), .B1(new_n709), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n485), .A2(G141), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT26), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n750), .B(new_n752), .C1(G129), .C2(new_n475), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n735), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n735), .B2(G32), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n744), .B(new_n748), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n742), .A2(new_n743), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n734), .B(new_n759), .C1(KEYINPUT90), .C2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G16), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G19), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n555), .B2(new_n763), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1341), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NOR2_X1   g342(.A1(G5), .A2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  INV_X1    g344(.A(G171), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n763), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n757), .A2(new_n758), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(KEYINPUT90), .B2(new_n761), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n763), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n624), .B2(new_n763), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n722), .A2(new_n762), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n763), .A2(G21), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G168), .B2(new_n763), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT92), .B(G1966), .Z(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT96), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n771), .A2(new_n767), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n783), .A2(new_n785), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G11), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n735), .B1(new_n792), .B2(G28), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT94), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n794), .A2(KEYINPUT94), .B1(new_n792), .B2(G28), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n636), .B2(new_n709), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT98), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n763), .A2(G20), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT23), .Z(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G299), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  INV_X1    g380(.A(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n781), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G6), .A2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G305), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n763), .A2(G22), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n763), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n814), .B1(new_n816), .B2(G1971), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G1971), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g393(.A1(G16), .A2(G23), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT86), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n821));
  NAND2_X1  g396(.A1(G288), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n510), .A2(G87), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n823), .A2(KEYINPUT87), .A3(new_n589), .A4(new_n590), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n825), .B2(new_n763), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT33), .B(G1976), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n818), .A2(KEYINPUT34), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT34), .B1(new_n818), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n710), .A2(G25), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n485), .A2(G131), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n833));
  INV_X1    g408(.A(G107), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(G2105), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G119), .B2(new_n475), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n831), .B1(new_n838), .B2(new_n710), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G1991), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT85), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n604), .A2(G16), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G16), .B2(G24), .ZN(new_n844));
  INV_X1    g419(.A(G1986), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n829), .A2(new_n830), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n809), .A2(new_n852), .ZN(G150));
  INV_X1    g428(.A(G150), .ZN(G311));
  AOI22_X1  g429(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n545), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n531), .B2(new_n534), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n509), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(G55), .B1(new_n606), .B2(new_n607), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  INV_X1    g438(.A(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n856), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT103), .B(G860), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  INV_X1    g444(.A(new_n856), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n858), .A2(KEYINPUT101), .A3(new_n860), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n554), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n554), .B1(new_n866), .B2(KEYINPUT102), .ZN(new_n878));
  AOI211_X1 g453(.A(new_n874), .B(new_n856), .C1(new_n861), .C2(new_n865), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT38), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n624), .A2(G559), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT39), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n867), .B1(new_n884), .B2(KEYINPUT39), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n869), .B1(new_n887), .B2(new_n888), .ZN(G145));
  AND2_X1   g464(.A1(new_n725), .A2(new_n730), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n755), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n754), .A2(new_n731), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n838), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n837), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n498), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n493), .A2(KEYINPUT105), .A3(new_n497), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(new_n741), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n741), .ZN(new_n902));
  OAI21_X1  g477(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G118), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n903), .A2(new_n904), .B1(new_n906), .B2(G2105), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n905), .A2(new_n907), .B1(new_n475), .B2(G130), .ZN(new_n908));
  INV_X1    g483(.A(G142), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n634), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n639), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n901), .A2(new_n902), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n901), .B2(new_n902), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n896), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n900), .B(new_n741), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n911), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n918), .A2(new_n894), .A3(new_n895), .A4(new_n913), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n636), .B(G160), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G162), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n916), .B2(new_n919), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(G395));
  XNOR2_X1  g503(.A(G166), .B(new_n604), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n825), .B(G305), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT42), .Z(new_n932));
  XNOR2_X1  g507(.A(new_n881), .B(new_n627), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n624), .A2(new_n934), .A3(G299), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n566), .A2(new_n571), .A3(new_n575), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n936), .B2(new_n618), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT108), .B1(new_n936), .B2(new_n618), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n624), .A2(new_n940), .A3(G299), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n935), .B2(new_n937), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n934), .B1(new_n624), .B2(G299), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n936), .A2(KEYINPUT109), .A3(new_n618), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n942), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n938), .A2(KEYINPUT41), .A3(new_n942), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n944), .B1(new_n933), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n944), .B(new_n957), .C1(new_n933), .C2(new_n954), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n932), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n932), .ZN(new_n960));
  OAI21_X1  g535(.A(G868), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g537(.A(new_n961), .B1(G868), .B2(new_n866), .ZN(G331));
  NAND3_X1  g538(.A1(new_n578), .A2(new_n580), .A3(G168), .ZN(new_n964));
  NAND3_X1  g539(.A1(G171), .A2(new_n584), .A3(new_n585), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n878), .A2(new_n879), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n873), .A2(new_n874), .A3(new_n554), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n964), .A2(new_n965), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n877), .A3(new_n880), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(KEYINPUT41), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n938), .A3(new_n942), .ZN(new_n973));
  INV_X1    g548(.A(new_n931), .ZN(new_n974));
  INV_X1    g549(.A(new_n950), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n973), .B(new_n974), .C1(new_n975), .C2(new_n972), .ZN(new_n976));
  AND4_X1   g551(.A1(new_n952), .A2(new_n969), .A3(new_n953), .A4(new_n971), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n943), .B1(new_n969), .B2(new_n971), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n931), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n979), .A3(new_n923), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n952), .A2(new_n969), .A3(new_n953), .A4(new_n971), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n969), .A2(new_n971), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n982), .B(new_n974), .C1(new_n983), .C2(new_n943), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n923), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n981), .B(KEYINPUT44), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n987), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n976), .A2(new_n979), .A3(new_n923), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n898), .A2(new_n995), .A3(new_n899), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n466), .A2(new_n469), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT114), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1000), .A2(G1996), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n755), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n890), .A2(new_n733), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n731), .A2(G2067), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n755), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1004), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  OR3_X1    g586(.A1(new_n1011), .A2(new_n841), .A3(new_n837), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1002), .B1(new_n1012), .B2(new_n1005), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1003), .B(KEYINPUT46), .Z(new_n1014));
  OAI21_X1  g589(.A(new_n1001), .B1(new_n754), .B2(new_n1007), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT47), .Z(new_n1017));
  XNOR2_X1  g592(.A(new_n837), .B(new_n841), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1011), .B1(new_n1001), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1000), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G290), .A2(G1986), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1013), .B(new_n1017), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n498), .A2(new_n995), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1384), .B1(new_n493), .B2(new_n497), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n999), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n714), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n898), .A2(KEYINPUT45), .A3(new_n995), .A4(new_n899), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n997), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1032), .A2(new_n999), .A3(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1031), .B(KEYINPUT119), .C1(new_n1034), .C2(G1971), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n999), .B1(new_n1027), .B2(KEYINPUT45), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1971), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1026), .A2(new_n1029), .A3(G2090), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1035), .A2(G8), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n521), .A2(new_n522), .A3(G8), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1031), .B1(new_n1034), .B2(G1971), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(G8), .A4(new_n1047), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1047), .B(G8), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n825), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n999), .B2(new_n1027), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n822), .A2(new_n824), .A3(KEYINPUT116), .A4(G1976), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  OR2_X1    g638(.A1(G305), .A2(G1981), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G305), .A2(G1981), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1064), .B(new_n1065), .C1(new_n1067), .C2(KEYINPUT49), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1060), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT117), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1074), .A2(KEYINPUT117), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1025), .A2(new_n997), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n784), .B1(new_n1078), .B2(new_n1037), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n747), .A3(new_n999), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(G286), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1049), .A2(new_n1055), .A3(new_n1077), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1047), .B1(new_n1050), .B2(G8), .ZN(new_n1089));
  NOR4_X1   g664(.A1(new_n1089), .A2(new_n1087), .A3(G286), .A4(new_n1084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n1055), .A3(new_n1077), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1049), .A2(new_n1055), .A3(new_n1077), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G168), .A2(new_n1059), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1094), .B2(KEYINPUT123), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1084), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1096), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1059), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1094), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1038), .A2(new_n1032), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1030), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n767), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1105), .A2(G2078), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1038), .B(new_n1110), .C1(new_n997), .C2(new_n1025), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G301), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1101), .A2(new_n1114), .A3(new_n1102), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1093), .A2(new_n1104), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1055), .ZN(new_n1117));
  INV_X1    g692(.A(G288), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1071), .A2(new_n1057), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1064), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1117), .A2(new_n1077), .B1(new_n1060), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1092), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n996), .A2(new_n997), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n999), .A3(new_n1032), .A4(new_n1110), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1107), .A2(new_n1109), .A3(G301), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1112), .B2(G301), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1126), .A2(new_n1127), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1112), .B2(G301), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1107), .A2(new_n1109), .A3(new_n1124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1130), .A2(KEYINPUT124), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1128), .A2(new_n1093), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1034), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1108), .A2(new_n806), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n566), .A2(new_n575), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT121), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n571), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(KEYINPUT121), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n936), .A2(KEYINPUT57), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1141), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(new_n1140), .A3(new_n1149), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(KEYINPUT122), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1149), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT61), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1034), .A2(new_n1008), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n999), .A2(new_n1027), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n554), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n1030), .A2(G1348), .B1(G2067), .B2(new_n1159), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(KEYINPUT60), .A3(new_n618), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1164), .B(new_n624), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1167), .A2(KEYINPUT60), .B1(KEYINPUT59), .B2(new_n1162), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1151), .A2(KEYINPUT61), .A3(new_n1152), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1157), .A2(new_n1166), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1164), .A2(new_n624), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1154), .B1(new_n1152), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1135), .A2(new_n1136), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1122), .B1(new_n1137), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n604), .A2(new_n845), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1020), .B1(new_n1021), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1019), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1024), .B1(new_n1174), .B2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g753(.A1(G227), .A2(new_n459), .ZN(new_n1180));
  OAI21_X1  g754(.A(new_n1180), .B1(new_n662), .B2(new_n663), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n703), .B1(new_n696), .B2(new_n701), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n705), .A2(new_n706), .A3(new_n702), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g758(.A(new_n1184), .B1(new_n925), .B2(new_n924), .ZN(new_n1185));
  INV_X1    g759(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g760(.A(KEYINPUT126), .B1(new_n991), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n1188));
  AOI211_X1 g762(.A(new_n1188), .B(new_n1185), .C1(new_n989), .C2(new_n990), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1189), .ZN(G308));
  NAND2_X1  g764(.A1(new_n991), .A2(new_n1186), .ZN(G225));
endmodule


