//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT70), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  AND4_X1   g044(.A1(new_n463), .A2(new_n465), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(G2104), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n469), .A2(new_n474), .A3(KEYINPUT68), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT68), .B1(new_n469), .B2(new_n474), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g054(.A(KEYINPUT69), .B(G125), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n473), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(G160));
  NAND4_X1  g060(.A1(new_n465), .A2(new_n468), .A3(G2105), .A4(new_n469), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(new_n489));
  MUX2_X1   g064(.A(G100), .B(G112), .S(G2105), .Z(new_n490));
  AOI22_X1  g065(.A1(new_n470), .A2(G136), .B1(G2104), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n489), .A2(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(new_n463), .A2(G102), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2105), .ZN(new_n494));
  AOI211_X1 g069(.A(KEYINPUT73), .B(new_n464), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n496));
  INV_X1    g071(.A(G102), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n498), .B2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n495), .A2(new_n499), .B1(new_n486), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n465), .A2(new_n468), .A3(new_n463), .A4(new_n469), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n505), .B1(new_n475), .B2(new_n476), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT74), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n531), .A2(new_n508), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n528), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n510), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n527), .A2(G52), .B1(G90), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n527), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  AND2_X1   g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n541), .A2(G81), .B1(new_n551), .B2(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n523), .A2(G53), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n549), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n508), .A2(KEYINPUT79), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(G78), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n510), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT77), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G91), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n572), .A2(KEYINPUT78), .A3(G91), .A4(new_n573), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n563), .A2(new_n570), .A3(new_n576), .A4(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n528), .A2(new_n535), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND3_X1  g155(.A1(new_n572), .A2(G87), .A3(new_n573), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n516), .B1(new_n549), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(G49), .B2(new_n523), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G288));
  NAND3_X1  g160(.A1(new_n572), .A2(G86), .A3(new_n573), .ZN(new_n586));
  OAI21_X1  g161(.A(G61), .B1(new_n547), .B2(new_n548), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(KEYINPUT80), .A3(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n523), .A2(G48), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n586), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n516), .B1(new_n510), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G47), .B2(new_n527), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n572), .A2(G92), .A3(new_n573), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n566), .A2(new_n567), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT81), .B(G66), .Z(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT82), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(G299), .B(KEYINPUT83), .Z(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n610), .B(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G860), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(G559), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT84), .ZN(G148));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n554), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n611), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(new_n626), .B2(new_n623), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT85), .ZN(G323));
  XOR2_X1   g203(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n629));
  XNOR2_X1  g204(.A(G323), .B(new_n629), .ZN(G282));
  NOR2_X1   g205(.A1(new_n475), .A2(new_n476), .ZN(new_n631));
  INV_X1    g206(.A(new_n471), .ZN(new_n632));
  OAI21_X1  g207(.A(KEYINPUT12), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT68), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n467), .A2(G2104), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n469), .A2(new_n474), .A3(KEYINPUT68), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT12), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(new_n471), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2100), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  AND2_X1   g222(.A1(G111), .A2(G2105), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(G99), .B2(new_n463), .ZN(new_n649));
  OAI22_X1  g224(.A1(new_n486), .A2(new_n647), .B1(new_n649), .B2(new_n464), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n470), .B2(G135), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT87), .B(KEYINPUT14), .Z(new_n660));
  XOR2_X1   g235(.A(G2427), .B(G2430), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n662), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  INV_X1    g251(.A(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .A3(new_n670), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n670), .B1(new_n677), .B2(KEYINPUT17), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n674), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n671), .A2(new_n674), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(new_n681), .B2(KEYINPUT17), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n676), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2096), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(G227));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT89), .Z(new_n689));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  INV_X1    g268(.A(new_n688), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n686), .A2(new_n687), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n691), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT91), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT91), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G24), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT92), .Z(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G290), .B2(new_n708), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  NOR2_X1   g288(.A1(G25), .A2(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n470), .A2(G131), .ZN(new_n715));
  INV_X1    g290(.A(G119), .ZN(new_n716));
  AND2_X1   g291(.A1(G107), .A2(G2105), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G95), .B2(new_n463), .ZN(new_n718));
  OAI22_X1  g293(.A1(new_n486), .A2(new_n716), .B1(new_n718), .B2(new_n464), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT90), .Z(new_n723));
  OR2_X1    g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n723), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n713), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G6), .B(G305), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT32), .B(G1981), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n708), .A2(G22), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G166), .B2(new_n708), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT94), .B(G1971), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G23), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g311(.A1(G288), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT93), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT33), .B(G1976), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n734), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT95), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n734), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT34), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n726), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n744), .A2(KEYINPUT34), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT36), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n749), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n705), .A2(G5), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G171), .B2(new_n705), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1961), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n708), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n554), .B2(new_n708), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1341), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n651), .A2(G29), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT103), .B(G28), .Z(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT30), .B2(new_n763), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT31), .B(G11), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n758), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G27), .A2(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G164), .B2(G29), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(G2078), .ZN(new_n771));
  INV_X1    g346(.A(G29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  INV_X1    g349(.A(G128), .ZN(new_n775));
  AND2_X1   g350(.A1(G116), .A2(G2105), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G104), .B2(new_n463), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n486), .A2(new_n775), .B1(new_n777), .B2(new_n464), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n470), .B2(G140), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(new_n772), .ZN(new_n780));
  INV_X1    g355(.A(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n770), .A2(G2078), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G21), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G168), .B2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT102), .Z(new_n787));
  AOI211_X1 g362(.A(new_n771), .B(new_n784), .C1(new_n787), .C2(G1966), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(new_n772), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G160), .B2(new_n772), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G2084), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n709), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT107), .B(KEYINPUT23), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G299), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n705), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n768), .A2(new_n788), .A3(new_n793), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G2084), .B2(new_n792), .ZN(new_n802));
  INV_X1    g377(.A(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT105), .B1(new_n803), .B2(G29), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n803), .A2(KEYINPUT105), .A3(G29), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n804), .B(new_n805), .C1(G162), .C2(new_n772), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT106), .B(KEYINPUT29), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G2090), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n611), .A2(G16), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G4), .B2(G16), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n810), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n787), .A2(KEYINPUT104), .A3(G1966), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT104), .B1(new_n787), .B2(G1966), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n815), .A2(new_n816), .B1(new_n809), .B2(new_n808), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n471), .A2(G103), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT25), .Z(new_n820));
  INV_X1    g395(.A(G139), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n502), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n639), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n463), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n824), .B2(KEYINPUT96), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(KEYINPUT96), .B2(new_n824), .ZN(new_n826));
  MUX2_X1   g401(.A(G33), .B(new_n826), .S(G29), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2072), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT101), .B1(G29), .B2(G32), .ZN(new_n830));
  NAND3_X1  g405(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT99), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT26), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n471), .A2(G105), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G129), .ZN(new_n838));
  INV_X1    g413(.A(G141), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n838), .A2(new_n486), .B1(new_n502), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G29), .ZN(new_n843));
  MUX2_X1   g418(.A(KEYINPUT101), .B(new_n830), .S(new_n843), .Z(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT27), .B(G1996), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n813), .A2(new_n811), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AND4_X1   g424(.A1(new_n802), .A2(new_n818), .A3(new_n829), .A4(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n755), .A2(new_n850), .ZN(G311));
  NAND2_X1  g426(.A1(new_n755), .A2(new_n850), .ZN(G150));
  NAND2_X1  g427(.A1(new_n527), .A2(G55), .ZN(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n549), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n541), .A2(G93), .B1(new_n856), .B2(G651), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  OR2_X1    g435(.A1(new_n553), .A2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n553), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n619), .A2(new_n625), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n620), .B1(new_n866), .B2(KEYINPUT39), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT108), .ZN(G145));
  XNOR2_X1  g445(.A(G160), .B(new_n651), .ZN(new_n871));
  INV_X1    g446(.A(G162), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT110), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n826), .A2(new_n841), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n826), .B2(new_n842), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n642), .B(new_n720), .ZN(new_n880));
  MUX2_X1   g455(.A(G106), .B(G118), .S(G2105), .Z(new_n881));
  AOI22_X1  g456(.A1(new_n487), .A2(G130), .B1(G2104), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G142), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n502), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n884), .ZN(new_n886));
  XNOR2_X1  g461(.A(G164), .B(new_n779), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n878), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(G160), .B(new_n651), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G162), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n873), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n876), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n873), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n902), .A2(new_n894), .A3(KEYINPUT109), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT109), .B1(new_n902), .B2(new_n894), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n900), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g481(.A1(new_n858), .A2(new_n623), .ZN(new_n907));
  XOR2_X1   g482(.A(KEYINPUT112), .B(KEYINPUT42), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n739), .B(new_n599), .ZN(new_n909));
  OR2_X1    g484(.A1(G303), .A2(G305), .ZN(new_n910));
  NAND2_X1  g485(.A1(G303), .A2(G305), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n739), .A2(new_n599), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n739), .A2(new_n599), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n914), .A2(new_n915), .B1(new_n911), .B2(new_n910), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n908), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(new_n912), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n911), .A4(new_n910), .ZN(new_n919));
  INV_X1    g494(.A(new_n908), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n626), .A2(new_n862), .A3(new_n861), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n797), .A2(new_n604), .A3(new_n609), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n610), .A2(G299), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n611), .A2(new_n625), .A3(new_n863), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n626), .B(new_n863), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n930), .A3(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n924), .A2(new_n933), .A3(new_n930), .A4(new_n925), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n926), .A2(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n922), .B(new_n928), .C1(new_n929), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n923), .A2(new_n927), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n940), .A2(new_n934), .A3(new_n932), .A4(new_n935), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n941), .A2(KEYINPUT114), .A3(new_n922), .A4(new_n928), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n928), .B1(new_n929), .B2(new_n936), .ZN(new_n944));
  INV_X1    g519(.A(new_n922), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n944), .A2(KEYINPUT113), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n907), .B1(new_n948), .B2(new_n623), .ZN(G295));
  OAI21_X1  g524(.A(new_n907), .B1(new_n948), .B2(new_n623), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n913), .A2(new_n916), .A3(KEYINPUT115), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n918), .B2(new_n919), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G301), .A2(G286), .ZN(new_n956));
  NAND3_X1  g531(.A1(G168), .A2(new_n540), .A3(new_n542), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n863), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n956), .A2(new_n861), .A3(new_n957), .A4(new_n862), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n931), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n931), .A2(new_n962), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n935), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n961), .A2(new_n926), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n955), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n936), .A2(new_n961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n918), .A2(new_n919), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n968), .B(new_n969), .C1(new_n926), .C2(new_n961), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n901), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g547(.A(new_n968), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n955), .B1(new_n973), .B2(new_n966), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n901), .A4(new_n970), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n951), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n975), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n974), .A2(KEYINPUT43), .A3(new_n901), .A4(new_n970), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT44), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(G397));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G164), .B2(G1384), .ZN(new_n983));
  INV_X1    g558(.A(new_n501), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n504), .A2(new_n506), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT117), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT45), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n480), .A2(new_n481), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT69), .B1(new_n639), .B2(G125), .ZN(new_n990));
  OAI21_X1  g565(.A(G2105), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n991), .A2(G40), .A3(new_n472), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n841), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(G1996), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT119), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n988), .A2(new_n992), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1996), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n779), .B(new_n781), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n998), .A2(new_n842), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n720), .B(new_n722), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n996), .B(new_n1000), .C1(new_n997), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1986), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n599), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT118), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n1003), .B2(new_n599), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1002), .B1(new_n993), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G303), .A2(G8), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n991), .A2(G40), .A3(new_n472), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G164), .B2(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G164), .B2(G1384), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n504), .A2(new_n506), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n1018), .C1(new_n1019), .C2(new_n501), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1017), .A2(new_n483), .A3(G40), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1971), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1015), .A2(new_n809), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1010), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G305), .A2(G1981), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n516), .B1(new_n587), .B2(new_n588), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(new_n591), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n541), .A2(G86), .B1(new_n523), .B2(G48), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1026), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n592), .A3(new_n593), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G1981), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n986), .A2(new_n991), .A3(G40), .A4(new_n472), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1033), .A2(G8), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n737), .A2(G1976), .A3(new_n738), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1039), .A3(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1037), .A2(new_n1039), .A3(G8), .A4(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1038), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(new_n809), .A3(new_n992), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1010), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(G8), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1025), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1966), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1021), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(new_n992), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(G2084), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1056), .B2(G286), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1058));
  INV_X1    g633(.A(G2084), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1015), .A2(new_n1059), .B1(new_n1021), .B2(new_n1053), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n1060), .B2(G168), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1024), .B1(new_n1060), .B2(G168), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1052), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n1065));
  INV_X1    g640(.A(G1961), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1055), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1021), .B2(G2078), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1021), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(G301), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1068), .A2(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n483), .A2(new_n1020), .A3(G40), .A4(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1067), .B(new_n1069), .C1(new_n988), .C2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1065), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1065), .B1(new_n1077), .B2(G171), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1073), .A2(G301), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1069), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1015), .A2(G1961), .B1(new_n988), .B2(new_n1076), .ZN(new_n1085));
  OAI21_X1  g660(.A(G171), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n1080), .A2(new_n1086), .A3(KEYINPUT54), .A4(new_n1082), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1064), .B(new_n1079), .C1(new_n1083), .C2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(G299), .B(KEYINPUT57), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1015), .A2(G1956), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT56), .B(G2072), .Z(new_n1091));
  NOR2_X1   g666(.A1(new_n1021), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1037), .A2(G2067), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1055), .B2(new_n811), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n619), .B2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1021), .A2(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1055), .A2(new_n799), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G299), .B(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n992), .A2(new_n781), .A3(new_n986), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(KEYINPUT60), .C1(new_n1015), .C2(G1348), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT124), .B1(new_n1104), .B2(new_n611), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1095), .A2(new_n1106), .A3(new_n619), .A4(KEYINPUT60), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n611), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1095), .A2(KEYINPUT60), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT125), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT61), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1093), .A2(new_n1101), .A3(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1037), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1037), .A2(KEYINPUT123), .A3(new_n1116), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1119), .B(new_n1120), .C1(G1996), .C2(new_n1021), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n554), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1124), .A3(new_n554), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1113), .A2(new_n1115), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1127), .B(new_n1128), .C1(KEYINPUT60), .C2(new_n1095), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1111), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1088), .B1(new_n1102), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1062), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT62), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1058), .A2(new_n1063), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n1052), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1051), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1038), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G288), .A2(G1976), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT120), .Z(new_n1145));
  OAI22_X1  g720(.A1(new_n1143), .A2(new_n1145), .B1(G1981), .B2(G305), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1037), .A2(G8), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1045), .A2(new_n1142), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G286), .A2(new_n1024), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1056), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT121), .B1(new_n1060), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1150), .B(new_n1151), .C1(new_n1158), .C2(new_n1052), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1157), .A2(new_n1045), .A3(new_n1051), .A4(new_n1025), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1151), .B1(new_n1161), .B2(new_n1150), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1141), .B(new_n1149), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1008), .B1(new_n1131), .B2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n715), .A2(new_n719), .A3(new_n722), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n996), .A2(new_n1000), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n779), .A2(new_n781), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT127), .B1(new_n1168), .B2(new_n993), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n998), .A2(KEYINPUT46), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n998), .A2(KEYINPUT46), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n993), .B1(new_n994), .B2(new_n999), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1006), .A2(new_n997), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT48), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1174), .B1(new_n1002), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1178), .B(new_n997), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1169), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1164), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g756(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n905), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n978), .A2(new_n979), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n1184), .A2(new_n1185), .ZN(G308));
  OR2_X1    g760(.A1(new_n1184), .A2(new_n1185), .ZN(G225));
endmodule


