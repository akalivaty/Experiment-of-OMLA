

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774;

  XNOR2_X1 U378 ( .A(n476), .B(n475), .ZN(n543) );
  XNOR2_X1 U379 ( .A(G107), .B(G116), .ZN(n515) );
  XNOR2_X1 U380 ( .A(G125), .B(G146), .ZN(n531) );
  NAND2_X1 U381 ( .A1(n357), .A2(n627), .ZN(n447) );
  XNOR2_X2 U382 ( .A(n587), .B(n586), .ZN(n627) );
  NOR2_X2 U383 ( .A1(n626), .A2(n625), .ZN(n357) );
  OR2_X2 U384 ( .A1(n578), .A2(n630), .ZN(n580) );
  XNOR2_X2 U385 ( .A(n543), .B(n542), .ZN(n749) );
  XNOR2_X1 U386 ( .A(n765), .B(G146), .ZN(n526) );
  XNOR2_X1 U387 ( .A(n600), .B(n455), .ZN(n717) );
  AND2_X1 U388 ( .A1(n717), .A2(n588), .ZN(n408) );
  AND2_X1 U389 ( .A1(n418), .A2(n416), .ZN(n358) );
  XNOR2_X2 U390 ( .A(n404), .B(n374), .ZN(n402) );
  XNOR2_X2 U391 ( .A(n386), .B(KEYINPUT94), .ZN(n629) );
  AND2_X2 U392 ( .A1(n415), .A2(n639), .ZN(n438) );
  OR2_X2 U393 ( .A1(n646), .A2(G902), .ZN(n528) );
  INV_X1 U394 ( .A(n705), .ZN(n579) );
  NAND2_X2 U395 ( .A1(n444), .A2(n442), .ZN(n386) );
  AND2_X2 U396 ( .A1(n446), .A2(n445), .ZN(n444) );
  NAND2_X2 U397 ( .A1(n564), .A2(n707), .ZN(n630) );
  XNOR2_X2 U398 ( .A(n407), .B(n592), .ZN(n733) );
  XNOR2_X2 U399 ( .A(n748), .B(n522), .ZN(n544) );
  XNOR2_X2 U400 ( .A(n413), .B(n521), .ZN(n748) );
  XNOR2_X2 U401 ( .A(n514), .B(n479), .ZN(n765) );
  XNOR2_X2 U402 ( .A(n532), .B(n478), .ZN(n514) );
  XNOR2_X1 U403 ( .A(n563), .B(KEYINPUT6), .ZN(n578) );
  INV_X1 U404 ( .A(G104), .ZN(n414) );
  XNOR2_X1 U405 ( .A(KEYINPUT67), .B(G101), .ZN(n522) );
  NOR2_X1 U406 ( .A1(n740), .A2(G953), .ZN(n741) );
  AND2_X1 U407 ( .A1(n421), .A2(n419), .ZN(n418) );
  AND2_X1 U408 ( .A1(n603), .A2(n602), .ZN(n696) );
  XNOR2_X1 U409 ( .A(n596), .B(n597), .ZN(n773) );
  XNOR2_X1 U410 ( .A(n403), .B(n372), .ZN(n774) );
  AND2_X1 U411 ( .A1(n606), .A2(n605), .ZN(n688) );
  NAND2_X1 U412 ( .A1(n402), .A2(n691), .ZN(n403) );
  NAND2_X1 U413 ( .A1(n605), .A2(n443), .ZN(n442) );
  NOR2_X1 U414 ( .A1(n693), .A2(n691), .ZN(n721) );
  NOR2_X1 U415 ( .A1(n580), .A2(n579), .ZN(n412) );
  XNOR2_X1 U416 ( .A(KEYINPUT101), .B(n609), .ZN(n693) );
  INV_X1 U417 ( .A(n710), .ZN(n631) );
  INV_X1 U418 ( .A(n578), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U420 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U421 ( .A(n456), .B(G119), .ZN(n476) );
  XNOR2_X1 U422 ( .A(n414), .B(KEYINPUT89), .ZN(n413) );
  XNOR2_X1 U423 ( .A(G140), .B(G137), .ZN(n523) );
  NAND2_X1 U424 ( .A1(n444), .A2(n442), .ZN(n387) );
  NAND2_X1 U425 ( .A1(n418), .A2(n416), .ZN(n360) );
  BUF_X1 U426 ( .A(n717), .Z(n361) );
  BUF_X1 U427 ( .A(n543), .Z(n362) );
  BUF_X1 U428 ( .A(n700), .Z(n363) );
  XNOR2_X2 U429 ( .A(n553), .B(n552), .ZN(n604) );
  NAND2_X1 U430 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U431 ( .A(n636), .ZN(n382) );
  OR2_X1 U432 ( .A1(n679), .A2(n694), .ZN(n383) );
  INV_X1 U433 ( .A(G237), .ZN(n482) );
  XNOR2_X1 U434 ( .A(n486), .B(KEYINPUT15), .ZN(n642) );
  XNOR2_X1 U435 ( .A(G902), .B(KEYINPUT88), .ZN(n486) );
  XNOR2_X1 U436 ( .A(KEYINPUT4), .B(G131), .ZN(n479) );
  XNOR2_X1 U437 ( .A(n492), .B(n434), .ZN(n513) );
  INV_X1 U438 ( .A(KEYINPUT8), .ZN(n434) );
  XNOR2_X1 U439 ( .A(n436), .B(n545), .ZN(n671) );
  XNOR2_X1 U440 ( .A(n749), .B(n544), .ZN(n436) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n638) );
  XNOR2_X1 U442 ( .A(n549), .B(n548), .ZN(n551) );
  XNOR2_X1 U443 ( .A(n547), .B(KEYINPUT91), .ZN(n548) );
  NOR2_X1 U444 ( .A1(G953), .A2(G237), .ZN(n505) );
  NOR2_X1 U445 ( .A1(n420), .A2(n364), .ZN(n419) );
  NOR2_X1 U446 ( .A1(n458), .A2(n457), .ZN(n420) );
  INV_X1 U447 ( .A(KEYINPUT77), .ZN(n454) );
  XNOR2_X1 U448 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n500) );
  XNOR2_X1 U449 ( .A(n531), .B(KEYINPUT10), .ZN(n763) );
  INV_X1 U450 ( .A(KEYINPUT33), .ZN(n411) );
  OR2_X1 U451 ( .A1(n560), .A2(n719), .ZN(n561) );
  XNOR2_X1 U452 ( .A(G113), .B(KEYINPUT71), .ZN(n475) );
  XNOR2_X1 U453 ( .A(n763), .B(n392), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n489), .B(KEYINPUT23), .ZN(n392) );
  XNOR2_X1 U455 ( .A(G128), .B(G110), .ZN(n489) );
  XOR2_X1 U456 ( .A(KEYINPUT7), .B(G122), .Z(n516) );
  INV_X1 U457 ( .A(G134), .ZN(n478) );
  NOR2_X1 U458 ( .A1(n719), .A2(n406), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n573), .B(n572), .ZN(n574) );
  NOR2_X1 U460 ( .A1(n591), .A2(n571), .ZN(n573) );
  XNOR2_X1 U461 ( .A(n577), .B(KEYINPUT32), .ZN(n625) );
  XNOR2_X1 U462 ( .A(n511), .B(n428), .ZN(n607) );
  XNOR2_X1 U463 ( .A(n512), .B(n429), .ZN(n428) );
  INV_X1 U464 ( .A(G475), .ZN(n429) );
  NAND2_X1 U465 ( .A1(n558), .A2(n371), .ZN(n445) );
  NOR2_X1 U466 ( .A1(n558), .A2(n371), .ZN(n443) );
  NOR2_X1 U467 ( .A1(n595), .A2(n594), .ZN(n606) );
  XNOR2_X1 U468 ( .A(n388), .B(KEYINPUT28), .ZN(n595) );
  NAND2_X1 U469 ( .A1(n631), .A2(n593), .ZN(n388) );
  INV_X1 U470 ( .A(KEYINPUT64), .ZN(n463) );
  INV_X1 U471 ( .A(KEYINPUT102), .ZN(n380) );
  NOR2_X1 U472 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U473 ( .A1(G237), .A2(G234), .ZN(n462) );
  INV_X1 U474 ( .A(G902), .ZN(n483) );
  XOR2_X1 U475 ( .A(KEYINPUT4), .B(KEYINPUT18), .Z(n538) );
  XNOR2_X1 U476 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n533) );
  XNOR2_X1 U477 ( .A(n440), .B(n439), .ZN(n700) );
  INV_X1 U478 ( .A(KEYINPUT45), .ZN(n439) );
  INV_X1 U479 ( .A(n716), .ZN(n406) );
  INV_X1 U480 ( .A(KEYINPUT38), .ZN(n455) );
  AND2_X1 U481 ( .A1(n575), .A2(n369), .ZN(n593) );
  XOR2_X1 U482 ( .A(G137), .B(KEYINPUT5), .Z(n471) );
  INV_X1 U483 ( .A(KEYINPUT74), .ZN(n472) );
  NAND2_X1 U484 ( .A1(n417), .A2(KEYINPUT80), .ZN(n416) );
  INV_X1 U485 ( .A(G953), .ZN(n753) );
  INV_X1 U486 ( .A(KEYINPUT65), .ZN(n453) );
  XNOR2_X1 U487 ( .A(n763), .B(n508), .ZN(n509) );
  XNOR2_X1 U488 ( .A(n394), .B(KEYINPUT43), .ZN(n393) );
  OR2_X1 U489 ( .A1(n574), .A2(n430), .ZN(n394) );
  INV_X1 U490 ( .A(KEYINPUT34), .ZN(n581) );
  INV_X1 U491 ( .A(KEYINPUT22), .ZN(n397) );
  NAND2_X1 U492 ( .A1(n387), .A2(n562), .ZN(n396) );
  XNOR2_X1 U493 ( .A(n561), .B(KEYINPUT103), .ZN(n562) );
  XNOR2_X1 U494 ( .A(KEYINPUT16), .B(G122), .ZN(n541) );
  XNOR2_X1 U495 ( .A(n493), .B(n389), .ZN(n744) );
  XNOR2_X1 U496 ( .A(n391), .B(n390), .ZN(n389) );
  XNOR2_X1 U497 ( .A(n490), .B(n491), .ZN(n390) );
  XNOR2_X1 U498 ( .A(n435), .B(n433), .ZN(n658) );
  NAND2_X1 U499 ( .A1(n513), .A2(G217), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n663), .B(KEYINPUT59), .ZN(n664) );
  XNOR2_X1 U501 ( .A(n526), .B(n400), .ZN(n646) );
  XNOR2_X1 U502 ( .A(n544), .B(n525), .ZN(n400) );
  OR2_X1 U503 ( .A1(n766), .A2(G952), .ZN(n742) );
  OR2_X1 U504 ( .A1(n735), .A2(n461), .ZN(n736) );
  NAND2_X1 U505 ( .A1(n460), .A2(n606), .ZN(n596) );
  INV_X1 U506 ( .A(n733), .ZN(n460) );
  INV_X1 U507 ( .A(n625), .ZN(n624) );
  XNOR2_X1 U508 ( .A(n401), .B(KEYINPUT31), .ZN(n694) );
  INV_X1 U509 ( .A(KEYINPUT100), .ZN(n425) );
  NOR2_X2 U510 ( .A1(n635), .A2(n634), .ZN(n679) );
  AND2_X1 U511 ( .A1(n402), .A2(n693), .ZN(n364) );
  BUF_X1 U512 ( .A(n551), .Z(n600) );
  NAND2_X1 U513 ( .A1(n393), .A2(n432), .ZN(n458) );
  INV_X1 U514 ( .A(n607), .ZN(n427) );
  XOR2_X1 U515 ( .A(KEYINPUT73), .B(n611), .Z(n365) );
  AND2_X1 U516 ( .A1(n624), .A2(n378), .ZN(n366) );
  AND2_X1 U517 ( .A1(n705), .A2(n628), .ZN(n367) );
  NOR2_X1 U518 ( .A1(n576), .A2(n359), .ZN(n368) );
  NOR2_X1 U519 ( .A1(n570), .A2(n560), .ZN(n369) );
  AND2_X1 U520 ( .A1(n579), .A2(n565), .ZN(n370) );
  XOR2_X1 U521 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n371) );
  XOR2_X1 U522 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n372) );
  XNOR2_X1 U523 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n373) );
  NAND2_X1 U524 ( .A1(n546), .A2(G214), .ZN(n716) );
  XNOR2_X1 U525 ( .A(n590), .B(KEYINPUT39), .ZN(n374) );
  OR2_X1 U526 ( .A1(n642), .A2(n641), .ZN(n375) );
  AND2_X1 U527 ( .A1(n623), .A2(KEYINPUT68), .ZN(n376) );
  XOR2_X1 U528 ( .A(n622), .B(KEYINPUT82), .Z(n377) );
  INV_X1 U529 ( .A(n378), .ZN(n379) );
  NAND2_X1 U530 ( .A1(n378), .A2(KEYINPUT68), .ZN(n626) );
  XNOR2_X2 U531 ( .A(n395), .B(KEYINPUT104), .ZN(n378) );
  XNOR2_X1 U532 ( .A(n379), .B(n566), .ZN(G12) );
  BUF_X1 U533 ( .A(n671), .Z(n384) );
  NAND2_X1 U534 ( .A1(n551), .A2(n716), .ZN(n553) );
  INV_X1 U535 ( .A(n559), .ZN(n608) );
  NAND2_X1 U536 ( .A1(n559), .A2(n427), .ZN(n426) );
  XNOR2_X1 U537 ( .A(n520), .B(G478), .ZN(n559) );
  INV_X1 U538 ( .A(n604), .ZN(n605) );
  NAND2_X1 U539 ( .A1(n600), .A2(n716), .ZN(n431) );
  NAND2_X1 U540 ( .A1(n579), .A2(n716), .ZN(n430) );
  AND2_X1 U541 ( .A1(n704), .A2(n632), .ZN(n588) );
  XNOR2_X1 U542 ( .A(n519), .B(n514), .ZN(n435) );
  INV_X1 U543 ( .A(n600), .ZN(n432) );
  NAND2_X1 U544 ( .A1(n717), .A2(n405), .ZN(n407) );
  NAND2_X1 U545 ( .A1(n361), .A2(n716), .ZN(n720) );
  AND2_X2 U546 ( .A1(n452), .A2(n699), .ZN(n385) );
  AND2_X2 U547 ( .A1(n452), .A2(n699), .ZN(n743) );
  XNOR2_X1 U548 ( .A(n412), .B(n411), .ZN(n725) );
  NAND2_X1 U549 ( .A1(n629), .A2(n725), .ZN(n582) );
  NAND2_X1 U550 ( .A1(n409), .A2(n370), .ZN(n395) );
  XNOR2_X2 U551 ( .A(n396), .B(n397), .ZN(n409) );
  AND2_X1 U552 ( .A1(n409), .A2(n368), .ZN(n577) );
  NAND2_X1 U553 ( .A1(n399), .A2(n398), .ZN(n441) );
  OR2_X2 U554 ( .A1(n627), .A2(KEYINPUT68), .ZN(n398) );
  NAND2_X1 U555 ( .A1(n627), .A2(n376), .ZN(n399) );
  NAND2_X1 U556 ( .A1(n387), .A2(n367), .ZN(n401) );
  NAND2_X1 U557 ( .A1(n408), .A2(n589), .ZN(n404) );
  NAND2_X1 U558 ( .A1(n409), .A2(n578), .ZN(n410) );
  XNOR2_X1 U559 ( .A(n410), .B(KEYINPUT84), .ZN(n568) );
  XNOR2_X2 U560 ( .A(n497), .B(n496), .ZN(n564) );
  NAND2_X1 U561 ( .A1(n441), .A2(n366), .ZN(n437) );
  NAND2_X1 U562 ( .A1(n774), .A2(n773), .ZN(n599) );
  XNOR2_X2 U563 ( .A(n481), .B(G472), .ZN(n563) );
  XNOR2_X1 U564 ( .A(n459), .B(n377), .ZN(n424) );
  NAND2_X1 U565 ( .A1(n447), .A2(KEYINPUT44), .ZN(n415) );
  INV_X1 U566 ( .A(n424), .ZN(n417) );
  NAND2_X1 U567 ( .A1(n424), .A2(n422), .ZN(n421) );
  NOR2_X1 U568 ( .A1(n423), .A2(KEYINPUT80), .ZN(n422) );
  INV_X1 U569 ( .A(n458), .ZN(n423) );
  XNOR2_X2 U570 ( .A(n426), .B(n425), .ZN(n691) );
  NOR2_X1 U571 ( .A1(n574), .A2(n431), .ZN(n601) );
  NAND2_X1 U572 ( .A1(n438), .A2(n437), .ZN(n440) );
  NAND2_X1 U573 ( .A1(n604), .A2(n371), .ZN(n446) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n663) );
  XNOR2_X2 U575 ( .A(n449), .B(n453), .ZN(n452) );
  NAND2_X1 U576 ( .A1(n450), .A2(n375), .ZN(n449) );
  XNOR2_X1 U577 ( .A(n451), .B(n454), .ZN(n450) );
  NAND2_X1 U578 ( .A1(n640), .A2(n358), .ZN(n451) );
  XNOR2_X2 U579 ( .A(G116), .B(KEYINPUT3), .ZN(n456) );
  INV_X1 U580 ( .A(KEYINPUT80), .ZN(n457) );
  NAND2_X1 U581 ( .A1(n621), .A2(n620), .ZN(n459) );
  INV_X1 U582 ( .A(n658), .ZN(n659) );
  XOR2_X1 U583 ( .A(n734), .B(KEYINPUT121), .Z(n461) );
  XNOR2_X1 U584 ( .A(n522), .B(n472), .ZN(n473) );
  INV_X1 U585 ( .A(n531), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n593), .A2(n359), .ZN(n571) );
  XNOR2_X1 U587 ( .A(n474), .B(n473), .ZN(n477) );
  INV_X1 U588 ( .A(KEYINPUT106), .ZN(n572) );
  XNOR2_X1 U589 ( .A(n495), .B(KEYINPUT25), .ZN(n496) );
  INV_X1 U590 ( .A(KEYINPUT83), .ZN(n590) );
  INV_X1 U591 ( .A(KEYINPUT122), .ZN(n738) );
  XNOR2_X1 U592 ( .A(n462), .B(KEYINPUT14), .ZN(n464) );
  NAND2_X1 U593 ( .A1(G952), .A2(n464), .ZN(n731) );
  NOR2_X1 U594 ( .A1(n731), .A2(G953), .ZN(n556) );
  XNOR2_X2 U595 ( .A(n463), .B(G953), .ZN(n766) );
  NAND2_X1 U596 ( .A1(G902), .A2(n464), .ZN(n465) );
  XOR2_X1 U597 ( .A(KEYINPUT92), .B(n465), .Z(n554) );
  INV_X1 U598 ( .A(n554), .ZN(n466) );
  NOR2_X1 U599 ( .A1(n766), .A2(n466), .ZN(n467) );
  XNOR2_X1 U600 ( .A(n467), .B(KEYINPUT105), .ZN(n468) );
  NOR2_X1 U601 ( .A1(G900), .A2(n468), .ZN(n469) );
  NOR2_X1 U602 ( .A1(n556), .A2(n469), .ZN(n570) );
  NAND2_X1 U603 ( .A1(n505), .A2(G210), .ZN(n470) );
  XNOR2_X1 U604 ( .A(n471), .B(n470), .ZN(n474) );
  XNOR2_X1 U605 ( .A(n362), .B(n477), .ZN(n480) );
  XNOR2_X2 U606 ( .A(G143), .B(G128), .ZN(n532) );
  XNOR2_X1 U607 ( .A(n480), .B(n526), .ZN(n653) );
  NAND2_X1 U608 ( .A1(n653), .A2(n483), .ZN(n481) );
  NAND2_X1 U609 ( .A1(n483), .A2(n482), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n563), .A2(n716), .ZN(n484) );
  XNOR2_X1 U611 ( .A(KEYINPUT30), .B(n484), .ZN(n485) );
  NOR2_X1 U612 ( .A1(n570), .A2(n485), .ZN(n589) );
  NAND2_X1 U613 ( .A1(n642), .A2(G234), .ZN(n487) );
  XNOR2_X1 U614 ( .A(n487), .B(KEYINPUT20), .ZN(n494) );
  NAND2_X1 U615 ( .A1(n494), .A2(G221), .ZN(n488) );
  XNOR2_X1 U616 ( .A(n488), .B(KEYINPUT21), .ZN(n560) );
  INV_X1 U617 ( .A(n560), .ZN(n707) );
  XOR2_X1 U618 ( .A(KEYINPUT24), .B(G119), .Z(n490) );
  INV_X1 U619 ( .A(n523), .ZN(n491) );
  NAND2_X1 U620 ( .A1(n766), .A2(G234), .ZN(n492) );
  NAND2_X1 U621 ( .A1(n513), .A2(G221), .ZN(n493) );
  NOR2_X1 U622 ( .A1(n744), .A2(G902), .ZN(n497) );
  NAND2_X1 U623 ( .A1(G217), .A2(n494), .ZN(n495) );
  INV_X1 U624 ( .A(n630), .ZN(n704) );
  AND2_X1 U625 ( .A1(n589), .A2(n704), .ZN(n530) );
  XNOR2_X1 U626 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n512) );
  XOR2_X1 U627 ( .A(G113), .B(G104), .Z(n499) );
  XNOR2_X1 U628 ( .A(G143), .B(G122), .ZN(n498) );
  XNOR2_X1 U629 ( .A(n499), .B(n498), .ZN(n504) );
  INV_X1 U630 ( .A(n500), .ZN(n502) );
  XNOR2_X1 U631 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n501) );
  XNOR2_X1 U632 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U633 ( .A(n504), .B(n503), .Z(n510) );
  XOR2_X1 U634 ( .A(G131), .B(G140), .Z(n507) );
  NAND2_X1 U635 ( .A1(n505), .A2(G214), .ZN(n506) );
  XNOR2_X1 U636 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U637 ( .A1(G902), .A2(n663), .ZN(n511) );
  XNOR2_X1 U638 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U639 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n517) );
  XNOR2_X1 U640 ( .A(n518), .B(n517), .ZN(n519) );
  NOR2_X1 U641 ( .A1(G902), .A2(n658), .ZN(n520) );
  NAND2_X1 U642 ( .A1(n427), .A2(n608), .ZN(n583) );
  XNOR2_X1 U643 ( .A(G107), .B(G110), .ZN(n521) );
  XNOR2_X1 U644 ( .A(n523), .B(KEYINPUT95), .ZN(n762) );
  NAND2_X1 U645 ( .A1(n766), .A2(G227), .ZN(n524) );
  XNOR2_X1 U646 ( .A(n762), .B(n524), .ZN(n525) );
  XNOR2_X1 U647 ( .A(KEYINPUT70), .B(G469), .ZN(n527) );
  XNOR2_X2 U648 ( .A(n528), .B(n527), .ZN(n632) );
  INV_X1 U649 ( .A(n632), .ZN(n594) );
  NOR2_X1 U650 ( .A1(n583), .A2(n594), .ZN(n529) );
  NAND2_X1 U651 ( .A1(n530), .A2(n529), .ZN(n550) );
  INV_X1 U652 ( .A(n532), .ZN(n534) );
  XNOR2_X1 U653 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U654 ( .A(n536), .B(n535), .ZN(n540) );
  NAND2_X1 U655 ( .A1(n766), .A2(G224), .ZN(n537) );
  XNOR2_X1 U656 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U657 ( .A(n540), .B(n539), .ZN(n545) );
  XNOR2_X1 U658 ( .A(n541), .B(KEYINPUT72), .ZN(n542) );
  NAND2_X1 U659 ( .A1(n671), .A2(n642), .ZN(n549) );
  NAND2_X1 U660 ( .A1(n546), .A2(G210), .ZN(n547) );
  NOR2_X1 U661 ( .A1(n550), .A2(n432), .ZN(n615) );
  XOR2_X1 U662 ( .A(G143), .B(n615), .Z(G45) );
  XNOR2_X1 U663 ( .A(G110), .B(KEYINPUT115), .ZN(n566) );
  INV_X1 U664 ( .A(KEYINPUT19), .ZN(n552) );
  NOR2_X1 U665 ( .A1(G898), .A2(n753), .ZN(n751) );
  NAND2_X1 U666 ( .A1(n751), .A2(n554), .ZN(n555) );
  XNOR2_X1 U667 ( .A(n555), .B(KEYINPUT93), .ZN(n557) );
  NOR2_X1 U668 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U669 ( .A1(n559), .A2(n607), .ZN(n719) );
  XNOR2_X2 U670 ( .A(n632), .B(KEYINPUT1), .ZN(n705) );
  INV_X1 U671 ( .A(n563), .ZN(n710) );
  INV_X1 U672 ( .A(n564), .ZN(n575) );
  NOR2_X1 U673 ( .A1(n631), .A2(n564), .ZN(n565) );
  XNOR2_X1 U674 ( .A(G101), .B(KEYINPUT112), .ZN(n569) );
  NAND2_X1 U675 ( .A1(n579), .A2(n564), .ZN(n567) );
  NOR2_X1 U676 ( .A1(n568), .A2(n567), .ZN(n637) );
  XOR2_X1 U677 ( .A(n569), .B(n637), .Z(G3) );
  INV_X1 U678 ( .A(n691), .ZN(n591) );
  XOR2_X1 U679 ( .A(G140), .B(n423), .Z(G42) );
  XOR2_X1 U680 ( .A(KEYINPUT87), .B(n705), .Z(n602) );
  NAND2_X1 U681 ( .A1(n602), .A2(n575), .ZN(n576) );
  XNOR2_X1 U682 ( .A(n624), .B(G119), .ZN(G21) );
  XNOR2_X1 U683 ( .A(n582), .B(n581), .ZN(n585) );
  XNOR2_X1 U684 ( .A(n583), .B(KEYINPUT75), .ZN(n584) );
  NAND2_X1 U685 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U686 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n586) );
  XNOR2_X1 U687 ( .A(n627), .B(G122), .ZN(G24) );
  XOR2_X1 U688 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n597) );
  XOR2_X1 U689 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n592) );
  INV_X1 U690 ( .A(KEYINPUT46), .ZN(n598) );
  XNOR2_X1 U691 ( .A(n599), .B(n598), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n601), .B(n373), .ZN(n603) );
  INV_X1 U693 ( .A(n696), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U695 ( .A(n721), .B(KEYINPUT76), .ZN(n636) );
  NOR2_X1 U696 ( .A1(n636), .A2(KEYINPUT47), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n688), .A2(n610), .ZN(n611) );
  NAND2_X1 U698 ( .A1(n612), .A2(n365), .ZN(n619) );
  INV_X1 U699 ( .A(n721), .ZN(n613) );
  NAND2_X1 U700 ( .A1(n688), .A2(n613), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n614), .A2(KEYINPUT47), .ZN(n617) );
  INV_X1 U702 ( .A(n615), .ZN(n616) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U704 ( .A(KEYINPUT48), .B(KEYINPUT69), .Z(n622) );
  INV_X1 U705 ( .A(KEYINPUT44), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n710), .A2(n630), .ZN(n628) );
  INV_X1 U707 ( .A(n629), .ZN(n635) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n700), .A2(n642), .ZN(n640) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n358), .A2(KEYINPUT2), .ZN(n643) );
  XOR2_X1 U714 ( .A(KEYINPUT78), .B(n643), .Z(n644) );
  INV_X1 U715 ( .A(n363), .ZN(n754) );
  NAND2_X1 U716 ( .A1(n644), .A2(n754), .ZN(n699) );
  NAND2_X1 U717 ( .A1(n743), .A2(G469), .ZN(n648) );
  XNOR2_X1 U718 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n649), .A2(n742), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U722 ( .A1(n743), .A2(G472), .ZN(n655) );
  XNOR2_X1 U723 ( .A(KEYINPUT86), .B(KEYINPUT111), .ZN(n651) );
  XOR2_X1 U724 ( .A(n651), .B(KEYINPUT62), .Z(n652) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n656), .A2(n742), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U728 ( .A1(n385), .A2(G478), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n661), .A2(n742), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U732 ( .A1(n743), .A2(G475), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n666), .A2(n742), .ZN(n668) );
  XOR2_X1 U735 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(G60) );
  NAND2_X1 U737 ( .A1(n385), .A2(G210), .ZN(n673) );
  XNOR2_X1 U738 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n669), .B(KEYINPUT55), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n384), .B(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n674), .A2(n742), .ZN(n676) );
  XNOR2_X1 U743 ( .A(KEYINPUT81), .B(KEYINPUT56), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(G51) );
  XOR2_X1 U745 ( .A(G104), .B(KEYINPUT113), .Z(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n691), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n678), .B(n677), .ZN(G6) );
  XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT26), .ZN(n683) );
  XOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n681) );
  NAND2_X1 U750 ( .A1(n679), .A2(n693), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(G9) );
  XOR2_X1 U753 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n685) );
  NAND2_X1 U754 ( .A1(n688), .A2(n693), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(n687) );
  XOR2_X1 U756 ( .A(G128), .B(KEYINPUT29), .Z(n686) );
  XNOR2_X1 U757 ( .A(n687), .B(n686), .ZN(G30) );
  NAND2_X1 U758 ( .A1(n688), .A2(n691), .ZN(n689) );
  XNOR2_X1 U759 ( .A(n689), .B(KEYINPUT118), .ZN(n690) );
  XNOR2_X1 U760 ( .A(G146), .B(n690), .ZN(G48) );
  NAND2_X1 U761 ( .A1(n691), .A2(n694), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(G113), .ZN(G15) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(G116), .ZN(G18) );
  XOR2_X1 U765 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n698) );
  XNOR2_X1 U766 ( .A(G125), .B(n696), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n698), .B(n697), .ZN(G27) );
  XOR2_X1 U768 ( .A(G134), .B(n364), .Z(G36) );
  INV_X1 U769 ( .A(n699), .ZN(n703) );
  NOR2_X1 U770 ( .A1(n360), .A2(n363), .ZN(n701) );
  NOR2_X1 U771 ( .A1(n701), .A2(KEYINPUT2), .ZN(n702) );
  NOR2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n737) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U774 ( .A(n706), .B(KEYINPUT50), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n707), .A2(n564), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n708), .B(KEYINPUT49), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U779 ( .A1(n713), .A2(n367), .ZN(n714) );
  XOR2_X1 U780 ( .A(KEYINPUT51), .B(n714), .Z(n715) );
  NOR2_X1 U781 ( .A1(n733), .A2(n715), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n361), .A2(n716), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U786 ( .A(n724), .B(KEYINPUT120), .ZN(n726) );
  INV_X1 U787 ( .A(n725), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n726), .A2(n732), .ZN(n727) );
  NOR2_X1 U789 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U790 ( .A(n729), .B(KEYINPUT52), .ZN(n730) );
  NOR2_X1 U791 ( .A1(n731), .A2(n730), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U793 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n741), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U796 ( .A(n742), .ZN(n747) );
  NAND2_X1 U797 ( .A1(n385), .A2(G217), .ZN(n745) );
  XNOR2_X1 U798 ( .A(n744), .B(n745), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(G66) );
  XOR2_X1 U800 ( .A(n748), .B(G101), .Z(n750) );
  XNOR2_X1 U801 ( .A(n749), .B(n750), .ZN(n752) );
  NOR2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n761) );
  NAND2_X1 U803 ( .A1(n754), .A2(n753), .ZN(n758) );
  NAND2_X1 U804 ( .A1(G953), .A2(G224), .ZN(n755) );
  XNOR2_X1 U805 ( .A(KEYINPUT61), .B(n755), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n756), .A2(G898), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U808 ( .A(n759), .B(KEYINPUT126), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(G69) );
  XNOR2_X1 U810 ( .A(n763), .B(n762), .ZN(n764) );
  XOR2_X1 U811 ( .A(n765), .B(n764), .Z(n768) );
  XNOR2_X1 U812 ( .A(n360), .B(n768), .ZN(n767) );
  NAND2_X1 U813 ( .A1(n767), .A2(n766), .ZN(n772) );
  XNOR2_X1 U814 ( .A(n768), .B(G227), .ZN(n769) );
  NAND2_X1 U815 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U816 ( .A1(n770), .A2(G953), .ZN(n771) );
  NAND2_X1 U817 ( .A1(n772), .A2(n771), .ZN(G72) );
  XNOR2_X1 U818 ( .A(G137), .B(n773), .ZN(G39) );
  XNOR2_X1 U819 ( .A(n774), .B(G131), .ZN(G33) );
endmodule

