

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U322 ( .A(n297), .B(n290), .ZN(n298) );
  INV_X1 U323 ( .A(KEYINPUT47), .ZN(n372) );
  XOR2_X1 U324 ( .A(n368), .B(n397), .Z(n570) );
  XOR2_X1 U325 ( .A(n305), .B(n304), .Z(n567) );
  AND2_X1 U326 ( .A1(G231GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U327 ( .A(n348), .B(n347), .Z(n559) );
  XNOR2_X1 U328 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n349) );
  XNOR2_X1 U329 ( .A(n350), .B(n349), .ZN(n371) );
  INV_X1 U330 ( .A(KEYINPUT67), .ZN(n353) );
  XNOR2_X1 U331 ( .A(n354), .B(n353), .ZN(n355) );
  NOR2_X1 U332 ( .A1(n380), .A2(n379), .ZN(n381) );
  INV_X1 U333 ( .A(KEYINPUT79), .ZN(n324) );
  XNOR2_X1 U334 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U335 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U336 ( .A(n325), .B(n324), .ZN(n326) );
  OR2_X1 U337 ( .A1(n457), .A2(n483), .ZN(n415) );
  XNOR2_X1 U338 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U339 ( .A(n415), .B(KEYINPUT117), .ZN(n558) );
  XNOR2_X1 U340 ( .A(KEYINPUT83), .B(n570), .ZN(n553) );
  INV_X1 U341 ( .A(G127GAT), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U343 ( .A(n453), .B(KEYINPUT50), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(G64GAT), .B(G57GAT), .Z(n292) );
  XNOR2_X1 U346 ( .A(G183GAT), .B(G155GAT), .ZN(n291) );
  XNOR2_X1 U347 ( .A(n292), .B(n291), .ZN(n305) );
  XOR2_X1 U348 ( .A(G71GAT), .B(KEYINPUT13), .Z(n308) );
  XOR2_X1 U349 ( .A(G1GAT), .B(G127GAT), .Z(n385) );
  XOR2_X1 U350 ( .A(n308), .B(n385), .Z(n294) );
  XNOR2_X1 U351 ( .A(G211GAT), .B(G78GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n299) );
  XOR2_X1 U353 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n296) );
  XNOR2_X1 U354 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U356 ( .A(n300), .B(KEYINPUT15), .Z(n303) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(G15GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n301), .B(KEYINPUT73), .ZN(n341) );
  XNOR2_X1 U359 ( .A(n341), .B(KEYINPUT12), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n307) );
  XNOR2_X1 U362 ( .A(KEYINPUT78), .B(KEYINPUT33), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n329) );
  XOR2_X1 U364 ( .A(n308), .B(G92GAT), .Z(n310) );
  XOR2_X1 U365 ( .A(G176GAT), .B(G64GAT), .Z(n406) );
  XNOR2_X1 U366 ( .A(G85GAT), .B(n406), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n312) );
  INV_X1 U368 ( .A(KEYINPUT75), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n322) );
  XNOR2_X1 U370 ( .A(G120GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n313), .B(G57GAT), .ZN(n388) );
  INV_X1 U372 ( .A(n388), .ZN(n315) );
  XOR2_X1 U373 ( .A(KEYINPUT76), .B(G78GAT), .Z(n439) );
  INV_X1 U374 ( .A(n439), .ZN(n314) );
  NAND2_X1 U375 ( .A1(n315), .A2(n314), .ZN(n317) );
  NAND2_X1 U376 ( .A1(n388), .A2(n439), .ZN(n316) );
  NAND2_X1 U377 ( .A1(n317), .A2(n316), .ZN(n319) );
  AND2_X1 U378 ( .A1(G230GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n320), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n327) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n323), .B(KEYINPUT77), .ZN(n356) );
  XNOR2_X1 U384 ( .A(n356), .B(KEYINPUT74), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n584) );
  XOR2_X1 U386 ( .A(n584), .B(KEYINPUT41), .Z(n519) );
  INV_X1 U387 ( .A(n519), .ZN(n564) );
  XOR2_X1 U388 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n331) );
  XNOR2_X1 U389 ( .A(KEYINPUT71), .B(KEYINPUT68), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n348) );
  XOR2_X1 U391 ( .A(G141GAT), .B(G197GAT), .Z(n333) );
  XNOR2_X1 U392 ( .A(G29GAT), .B(G36GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U394 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n335) );
  XNOR2_X1 U395 ( .A(G113GAT), .B(G1GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U397 ( .A(n337), .B(n336), .Z(n346) );
  XOR2_X1 U398 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n339) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G43GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(KEYINPUT7), .B(n340), .Z(n362) );
  XOR2_X1 U402 ( .A(G169GAT), .B(G8GAT), .Z(n410) );
  XOR2_X1 U403 ( .A(n410), .B(n341), .Z(n343) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n362), .B(n344), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  NOR2_X1 U408 ( .A1(n564), .A2(n559), .ZN(n350) );
  INV_X1 U409 ( .A(n567), .ZN(n587) );
  XOR2_X1 U410 ( .A(KEYINPUT81), .B(KEYINPUT10), .Z(n352) );
  XNOR2_X1 U411 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n358) );
  NAND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n364) );
  XOR2_X1 U415 ( .A(KEYINPUT82), .B(G92GAT), .Z(n360) );
  XNOR2_X1 U416 ( .A(G190GAT), .B(G218GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U418 ( .A(G36GAT), .B(n361), .Z(n403) );
  XNOR2_X1 U419 ( .A(n362), .B(n403), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT80), .B(G85GAT), .Z(n366) );
  XNOR2_X1 U422 ( .A(G134GAT), .B(G162GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(G29GAT), .B(n367), .Z(n397) );
  INV_X1 U425 ( .A(n570), .ZN(n369) );
  NOR2_X1 U426 ( .A1(n587), .A2(n369), .ZN(n370) );
  AND2_X1 U427 ( .A1(n371), .A2(n370), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n380) );
  XOR2_X1 U429 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n375) );
  XNOR2_X1 U430 ( .A(KEYINPUT36), .B(n553), .ZN(n589) );
  NAND2_X1 U431 ( .A1(n589), .A2(n587), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n376) );
  NOR2_X1 U433 ( .A1(n584), .A2(n376), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n377), .B(KEYINPUT116), .ZN(n378) );
  INV_X1 U435 ( .A(n559), .ZN(n580) );
  AND2_X1 U436 ( .A1(n378), .A2(n559), .ZN(n379) );
  XNOR2_X1 U437 ( .A(KEYINPUT48), .B(n381), .ZN(n457) );
  XOR2_X1 U438 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n383) );
  XNOR2_X1 U439 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U441 ( .A(n384), .B(KEYINPUT5), .Z(n387) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT6), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U444 ( .A(G113GAT), .B(KEYINPUT0), .Z(n427) );
  XOR2_X1 U445 ( .A(n388), .B(n427), .Z(n390) );
  NAND2_X1 U446 ( .A1(G225GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n399) );
  XNOR2_X1 U449 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n393), .B(KEYINPUT93), .ZN(n394) );
  XOR2_X1 U451 ( .A(n394), .B(KEYINPUT2), .Z(n396) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(G155GAT), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n446) );
  XNOR2_X1 U454 ( .A(n446), .B(n397), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n481) );
  XOR2_X1 U456 ( .A(KEYINPUT96), .B(n481), .Z(n537) );
  XOR2_X1 U457 ( .A(KEYINPUT21), .B(G211GAT), .Z(n401) );
  XNOR2_X1 U458 ( .A(KEYINPUT91), .B(G204GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U460 ( .A(G197GAT), .B(n402), .Z(n450) );
  XNOR2_X1 U461 ( .A(n450), .B(n403), .ZN(n414) );
  XOR2_X1 U462 ( .A(G183GAT), .B(KEYINPUT18), .Z(n405) );
  XNOR2_X1 U463 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n426) );
  XOR2_X1 U465 ( .A(n406), .B(n426), .Z(n408) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U468 ( .A(n409), .B(KEYINPUT98), .Z(n412) );
  XNOR2_X1 U469 ( .A(n410), .B(KEYINPUT97), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U471 ( .A(n414), .B(n413), .Z(n539) );
  XNOR2_X1 U472 ( .A(n539), .B(KEYINPUT27), .ZN(n477) );
  NAND2_X1 U473 ( .A1(n537), .A2(n477), .ZN(n483) );
  XOR2_X1 U474 ( .A(G176GAT), .B(KEYINPUT20), .Z(n417) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(KEYINPUT90), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n435) );
  XOR2_X1 U477 ( .A(G190GAT), .B(G134GAT), .Z(n419) );
  XNOR2_X1 U478 ( .A(G43GAT), .B(G99GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U480 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n421) );
  XNOR2_X1 U481 ( .A(G127GAT), .B(G120GAT), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n423), .B(n422), .Z(n433) );
  XOR2_X1 U484 ( .A(G71GAT), .B(KEYINPUT65), .Z(n425) );
  XNOR2_X1 U485 ( .A(G15GAT), .B(KEYINPUT89), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U487 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n542) );
  INV_X1 U493 ( .A(n542), .ZN(n529) );
  XOR2_X1 U494 ( .A(G148GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U495 ( .A(G22GAT), .B(G106GAT), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U497 ( .A(n438), .B(G218GAT), .Z(n441) );
  XNOR2_X1 U498 ( .A(G50GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U500 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n443) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U503 ( .A(n445), .B(n444), .Z(n448) );
  XNOR2_X1 U504 ( .A(n446), .B(KEYINPUT23), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n475) );
  XOR2_X1 U507 ( .A(KEYINPUT28), .B(n475), .Z(n531) );
  INV_X1 U508 ( .A(n531), .ZN(n544) );
  NOR2_X1 U509 ( .A1(n529), .A2(n544), .ZN(n451) );
  NAND2_X1 U510 ( .A1(n558), .A2(n451), .ZN(n452) );
  XOR2_X1 U511 ( .A(KEYINPUT118), .B(n452), .Z(n554) );
  INV_X1 U512 ( .A(n554), .ZN(n550) );
  NOR2_X1 U513 ( .A1(n567), .A2(n550), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(n454), .ZN(G1342GAT) );
  XNOR2_X1 U515 ( .A(KEYINPUT123), .B(n539), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT54), .ZN(n459) );
  INV_X1 U518 ( .A(n537), .ZN(n522) );
  NAND2_X1 U519 ( .A1(n459), .A2(n522), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT64), .ZN(n579) );
  NOR2_X1 U521 ( .A1(n579), .A2(n475), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT55), .ZN(n462) );
  NOR2_X2 U523 ( .A1(n529), .A2(n462), .ZN(n574) );
  NAND2_X1 U524 ( .A1(n574), .A2(n519), .ZN(n465) );
  XOR2_X1 U525 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n463) );
  XNOR2_X1 U526 ( .A(n463), .B(G176GAT), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  NAND2_X1 U528 ( .A1(n574), .A2(n553), .ZN(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n467) );
  INV_X1 U530 ( .A(G190GAT), .ZN(n466) );
  NOR2_X1 U531 ( .A1(n559), .A2(n584), .ZN(n502) );
  NOR2_X1 U532 ( .A1(n567), .A2(n553), .ZN(n471) );
  XNOR2_X1 U533 ( .A(KEYINPUT16), .B(KEYINPUT86), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n471), .B(n470), .ZN(n487) );
  XOR2_X1 U535 ( .A(KEYINPUT99), .B(KEYINPUT25), .Z(n474) );
  INV_X1 U536 ( .A(n539), .ZN(n527) );
  NOR2_X1 U537 ( .A1(n529), .A2(n527), .ZN(n472) );
  NOR2_X1 U538 ( .A1(n475), .A2(n472), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n475), .A2(n529), .ZN(n476) );
  XOR2_X1 U541 ( .A(n476), .B(KEYINPUT26), .Z(n577) );
  NAND2_X1 U542 ( .A1(n477), .A2(n577), .ZN(n478) );
  NAND2_X1 U543 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U544 ( .A(KEYINPUT100), .B(n480), .ZN(n482) );
  NAND2_X1 U545 ( .A1(n482), .A2(n481), .ZN(n486) );
  NOR2_X1 U546 ( .A1(n544), .A2(n483), .ZN(n484) );
  NAND2_X1 U547 ( .A1(n529), .A2(n484), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n499) );
  NAND2_X1 U549 ( .A1(n487), .A2(n499), .ZN(n520) );
  INV_X1 U550 ( .A(n520), .ZN(n488) );
  NAND2_X1 U551 ( .A1(n502), .A2(n488), .ZN(n496) );
  NOR2_X1 U552 ( .A1(n522), .A2(n496), .ZN(n490) );
  XNOR2_X1 U553 ( .A(KEYINPUT101), .B(KEYINPUT34), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U555 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U556 ( .A1(n527), .A2(n496), .ZN(n492) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(n492), .Z(n493) );
  XNOR2_X1 U558 ( .A(G8GAT), .B(n493), .ZN(G1325GAT) );
  NOR2_X1 U559 ( .A1(n529), .A2(n496), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U561 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n531), .A2(n496), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(G1327GAT) );
  NAND2_X1 U565 ( .A1(n589), .A2(n499), .ZN(n500) );
  NOR2_X1 U566 ( .A1(n587), .A2(n500), .ZN(n501) );
  XNOR2_X1 U567 ( .A(KEYINPUT37), .B(n501), .ZN(n536) );
  INV_X1 U568 ( .A(n536), .ZN(n503) );
  NAND2_X1 U569 ( .A1(n503), .A2(n502), .ZN(n505) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n517), .A2(n522), .ZN(n510) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n507) );
  XNOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(KEYINPUT104), .B(n508), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  NOR2_X1 U578 ( .A1(n527), .A2(n517), .ZN(n511) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(n511), .Z(n512) );
  XNOR2_X1 U580 ( .A(G36GAT), .B(n512), .ZN(G1329GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n514) );
  XNOR2_X1 U582 ( .A(G43GAT), .B(KEYINPUT110), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(n516) );
  NOR2_X1 U584 ( .A1(n529), .A2(n517), .ZN(n515) );
  XOR2_X1 U585 ( .A(n516), .B(n515), .Z(G1330GAT) );
  NOR2_X1 U586 ( .A1(n517), .A2(n531), .ZN(n518) );
  XOR2_X1 U587 ( .A(G50GAT), .B(n518), .Z(G1331GAT) );
  NAND2_X1 U588 ( .A1(n559), .A2(n519), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n535), .A2(n520), .ZN(n521) );
  XOR2_X1 U590 ( .A(KEYINPUT112), .B(n521), .Z(n532) );
  NOR2_X1 U591 ( .A1(n522), .A2(n532), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n524) );
  XNOR2_X1 U593 ( .A(G57GAT), .B(KEYINPUT113), .ZN(n523) );
  XNOR2_X1 U594 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1332GAT) );
  NOR2_X1 U596 ( .A1(n527), .A2(n532), .ZN(n528) );
  XOR2_X1 U597 ( .A(G64GAT), .B(n528), .Z(G1333GAT) );
  NOR2_X1 U598 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U599 ( .A(G71GAT), .B(n530), .Z(G1334GAT) );
  NOR2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(G1335GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n537), .A2(n545), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G85GAT), .B(n538), .ZN(G1336GAT) );
  NAND2_X1 U606 ( .A1(n539), .A2(n545), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n540), .B(KEYINPUT114), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G92GAT), .B(n541), .ZN(G1337GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n545), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT44), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G106GAT), .B(n547), .ZN(G1339GAT) );
  XNOR2_X1 U614 ( .A(G113GAT), .B(KEYINPUT119), .ZN(n549) );
  NOR2_X1 U615 ( .A1(n559), .A2(n550), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1340GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n564), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1341GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G134GAT), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n577), .ZN(n569) );
  NOR2_X1 U625 ( .A1(n559), .A2(n569), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n564), .A2(n569), .ZN(n565) );
  XOR2_X1 U632 ( .A(n566), .B(n565), .Z(G1345GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n569), .ZN(n568) );
  XOR2_X1 U634 ( .A(G155GAT), .B(n568), .Z(G1346GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n571), .Z(G1347GAT) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n580), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1348GAT) );
  XOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U641 ( .A1(n574), .A2(n587), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  INV_X1 U644 ( .A(n577), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n590), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n590), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

