//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n190), .A2(KEYINPUT65), .A3(G137), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT65), .B1(new_n190), .B2(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n192), .B2(G134), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n190), .A2(KEYINPUT65), .A3(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n191), .A2(new_n202), .A3(new_n193), .A4(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(new_n200), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(KEYINPUT66), .A3(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT0), .B(G128), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  MUX2_X1   g028(.A(new_n208), .B(new_n209), .S(new_n214), .Z(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n207), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n192), .A2(KEYINPUT67), .A3(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n190), .A2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT67), .B1(new_n192), .B2(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n211), .A3(new_n213), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n212), .A3(G143), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n210), .B(G146), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n221), .B(new_n227), .C1(G131), .C2(new_n204), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n234), .A2(KEYINPUT69), .A3(G116), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G119), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n233), .B(new_n235), .C1(new_n236), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n234), .B2(G116), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(new_n238), .A3(G119), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(G116), .B2(new_n234), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT70), .A3(new_n233), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n244), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n233), .B1(new_n248), .B2(new_n235), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT72), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n252));
  AOI211_X1 g066(.A(new_n252), .B(new_n249), .C1(new_n242), .C2(new_n246), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n216), .B(new_n228), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(G101), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n256), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n216), .A2(new_n228), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n199), .A2(new_n265), .A3(new_n227), .A4(new_n221), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n216), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n263), .A2(KEYINPUT30), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n247), .A2(new_n250), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT71), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n206), .A2(new_n207), .A3(new_n215), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n266), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n228), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n270), .A4(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n188), .B(new_n262), .C1(new_n271), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n260), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n254), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n267), .A2(new_n270), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(new_n254), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n279), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n274), .A2(new_n270), .A3(new_n275), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n261), .B1(new_n290), .B2(new_n276), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n287), .B1(new_n291), .B2(new_n188), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n262), .B1(new_n271), .B2(new_n277), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n187), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n282), .A2(new_n284), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n188), .A2(new_n291), .B1(new_n299), .B2(new_n279), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT73), .B1(new_n293), .B2(KEYINPUT31), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n291), .A2(new_n287), .A3(new_n188), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n304), .A3(KEYINPUT77), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n295), .A2(new_n297), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G472), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n216), .A2(new_n228), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n270), .A2(new_n252), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n249), .B1(new_n242), .B2(new_n246), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n254), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n280), .B1(new_n315), .B2(new_n254), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(KEYINPUT29), .A3(new_n260), .A4(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT75), .B(G902), .Z(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(KEYINPUT76), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT76), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n254), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n290), .B2(new_n276), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n260), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n299), .A2(new_n279), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT29), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n310), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n309), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT9), .B(G234), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G221), .B1(new_n337), .B2(G902), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n338), .B(KEYINPUT83), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G140), .ZN(new_n341));
  INV_X1    g155(.A(G227), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G953), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n341), .B(new_n343), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G104), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n346), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  INV_X1    g162(.A(G107), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(G107), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G101), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(G101), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n347), .A2(new_n350), .A3(new_n356), .A4(new_n351), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n215), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n349), .A2(G104), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n346), .A2(G107), .ZN(new_n361));
  OAI21_X1  g175(.A(G101), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n227), .A2(KEYINPUT10), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n357), .A2(new_n362), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n227), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(KEYINPUT84), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT84), .B1(new_n369), .B2(new_n370), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n359), .B(new_n367), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n206), .A2(new_n207), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT86), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n375), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n368), .B(new_n227), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT12), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT12), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n345), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n375), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n369), .A2(new_n370), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n371), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n390), .A3(new_n359), .A4(new_n367), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n374), .A2(new_n378), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n344), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(KEYINPUT87), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT87), .B1(new_n384), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(G469), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  INV_X1    g212(.A(G902), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n392), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n345), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n381), .B2(new_n382), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n378), .A2(new_n379), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT12), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT88), .A3(new_n380), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(new_n391), .A3(new_n408), .A4(new_n344), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n323), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n400), .B1(new_n410), .B2(new_n398), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n340), .B1(new_n397), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT82), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT24), .B(G110), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT80), .ZN(new_n416));
  XNOR2_X1  g230(.A(G119), .B(G128), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT23), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(G119), .B2(new_n222), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n234), .A2(KEYINPUT23), .A3(G128), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(G119), .B2(new_n222), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n416), .A2(new_n417), .B1(G110), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G125), .B(G140), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT16), .ZN(new_n424));
  INV_X1    g238(.A(G125), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n425), .A2(KEYINPUT16), .A3(G140), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(G146), .A3(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n212), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n422), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n212), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n427), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n416), .A2(new_n417), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n421), .A2(G110), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT22), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(G137), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n431), .A2(new_n441), .A3(new_n437), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OR4_X1    g260(.A1(new_n414), .A2(new_n446), .A3(KEYINPUT25), .A4(new_n323), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT78), .B(G217), .ZN(new_n448));
  INV_X1    g262(.A(G234), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n323), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT79), .ZN(new_n451));
  OAI22_X1  g265(.A1(new_n446), .A2(new_n323), .B1(new_n414), .B2(KEYINPUT25), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(G902), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n413), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT96), .B1(new_n210), .B2(G128), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n222), .A3(G143), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n210), .A2(G128), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n190), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G116), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n238), .A2(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G107), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n349), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT97), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT13), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n464), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n473), .B1(new_n464), .B2(new_n475), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n465), .A2(new_n474), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI221_X1 g293(.A(new_n466), .B1(new_n471), .B2(new_n472), .C1(new_n479), .C2(new_n190), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n238), .A2(KEYINPUT14), .A3(G122), .ZN(new_n481));
  OAI211_X1 g295(.A(G107), .B(new_n481), .C1(new_n470), .C2(KEYINPUT14), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n464), .A2(new_n465), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n471), .B1(new_n486), .B2(new_n466), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT99), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT99), .B1(new_n484), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n480), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n336), .A2(new_n258), .A3(new_n448), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n480), .B(new_n493), .C1(new_n488), .C2(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n460), .B1(new_n495), .B2(new_n324), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n323), .B(new_n459), .C1(new_n492), .C2(new_n494), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT100), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT100), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n496), .B2(new_n497), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n434), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n257), .A2(new_n258), .A3(G214), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(G143), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(new_n198), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n505), .B(new_n198), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n503), .B(new_n507), .C1(new_n508), .C2(KEYINPUT17), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n346), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(KEYINPUT18), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n505), .B1(new_n513), .B2(new_n198), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n423), .B(new_n212), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n423), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n423), .A2(new_n518), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n212), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n428), .A2(new_n429), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT95), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n428), .A2(new_n524), .A3(new_n429), .A4(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n508), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n526), .A2(new_n516), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n517), .B1(new_n527), .B2(new_n511), .ZN(new_n528));
  INV_X1    g342(.A(G475), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(KEYINPUT20), .A3(new_n529), .A4(new_n399), .ZN(new_n530));
  INV_X1    g344(.A(new_n517), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n511), .B1(new_n509), .B2(new_n516), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n399), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G475), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n511), .B1(new_n526), .B2(new_n516), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n529), .B(new_n399), .C1(new_n535), .C2(new_n531), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G952), .ZN(new_n540));
  AOI211_X1 g354(.A(G953), .B(new_n540), .C1(G234), .C2(G237), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n258), .B(new_n324), .C1(G234), .C2(G237), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT21), .B(G898), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n502), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT89), .B(KEYINPUT5), .Z(new_n547));
  OAI21_X1  g361(.A(KEYINPUT90), .B1(new_n547), .B2(new_n235), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT89), .B(KEYINPUT5), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n550), .A3(G116), .A4(new_n234), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(G113), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n245), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n549), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n247), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n363), .B(KEYINPUT85), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n358), .A2(new_n354), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n313), .ZN(new_n558));
  XOR2_X1   g372(.A(G110), .B(G122), .Z(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  OAI221_X1 g375(.A(new_n561), .B1(new_n557), .B2(new_n313), .C1(new_n555), .C2(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT6), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT6), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n565), .A3(new_n559), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT91), .A4(KEYINPUT6), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  MUX2_X1   g383(.A(new_n227), .B(new_n215), .S(G125), .Z(new_n570));
  INV_X1    g384(.A(G224), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G953), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n570), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n572), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n570), .A2(KEYINPUT92), .A3(KEYINPUT7), .A4(new_n573), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n578), .A2(new_n562), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n555), .A2(new_n368), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n552), .B1(KEYINPUT5), .B2(new_n245), .ZN(new_n583));
  INV_X1    g397(.A(new_n247), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n368), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n559), .B(KEYINPUT8), .Z(new_n586));
  AND3_X1   g400(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n399), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT93), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n575), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n574), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n567), .B2(new_n568), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n591), .B1(new_n595), .B2(new_n588), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G214), .B1(G237), .B2(G902), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT94), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n600));
  INV_X1    g414(.A(new_n598), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n600), .B(new_n601), .C1(new_n593), .C2(new_n596), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n546), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n335), .A2(new_n457), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  AOI21_X1  g420(.A(new_n310), .B1(new_n303), .B2(new_n324), .ZN(new_n607));
  NOR4_X1   g421(.A1(new_n413), .A2(new_n607), .A3(new_n306), .A4(new_n456), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT101), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n601), .B1(new_n593), .B2(new_n596), .ZN(new_n610));
  INV_X1    g424(.A(new_n545), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n490), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n495), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n492), .A2(new_n614), .A3(KEYINPUT33), .A4(new_n494), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n324), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G478), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n495), .A2(new_n458), .A3(new_n324), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n539), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n609), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  INV_X1    g440(.A(new_n539), .ZN(new_n627));
  AND4_X1   g441(.A1(new_n610), .A2(new_n627), .A3(new_n502), .A4(new_n611), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n609), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  OAI21_X1  g445(.A(G472), .B1(new_n295), .B2(new_n323), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n297), .B2(new_n295), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n442), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n438), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n454), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n453), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n412), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n603), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT37), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G110), .ZN(G12));
  INV_X1    g455(.A(new_n542), .ZN(new_n642));
  OR3_X1    g456(.A1(new_n642), .A2(KEYINPUT103), .A3(G900), .ZN(new_n643));
  INV_X1    g457(.A(new_n541), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT103), .B1(new_n642), .B2(G900), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n502), .A2(new_n627), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n638), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n335), .A2(new_n610), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n597), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT38), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n329), .A2(new_n279), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n399), .B1(new_n316), .B2(new_n260), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n653), .B1(new_n309), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n646), .B(KEYINPUT39), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n412), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n637), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n502), .A2(new_n598), .A3(new_n539), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n657), .A2(new_n662), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  INV_X1    g480(.A(new_n622), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n646), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n413), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n335), .A2(new_n610), .A3(new_n637), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT105), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n212), .ZN(G48));
  INV_X1    g486(.A(new_n456), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n410), .A2(new_n398), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n410), .A2(new_n398), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n338), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT106), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n674), .A2(new_n679), .A3(new_n675), .A4(new_n338), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n335), .A2(new_n673), .A3(new_n623), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n335), .A2(new_n673), .A3(new_n628), .A4(new_n681), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  AND3_X1   g500(.A1(new_n678), .A2(new_n610), .A3(new_n680), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n335), .A2(new_n546), .A3(new_n637), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  NAND2_X1  g503(.A1(new_n290), .A2(new_n276), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n188), .B1(new_n690), .B2(new_n262), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n260), .B1(new_n319), .B2(new_n321), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT74), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n254), .B2(new_n280), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n320), .A2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n694), .B(new_n280), .C1(new_n315), .C2(new_n254), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n279), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n698), .B(new_n699), .C1(new_n188), .C2(new_n291), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n693), .A2(new_n278), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n701), .A2(new_n702), .A3(new_n296), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n701), .B2(new_n296), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n607), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n664), .A2(new_n597), .A3(new_n611), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n681), .A4(new_n673), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  INV_X1    g522(.A(new_n646), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n622), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n687), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n703), .A2(new_n704), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n632), .A4(new_n637), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n701), .A2(new_n296), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT108), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n701), .A2(new_n702), .A3(new_n296), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n632), .A3(new_n637), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n711), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT110), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  NAND3_X1  g536(.A1(new_n384), .A2(G469), .A3(new_n393), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n411), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n338), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n593), .A2(new_n598), .A3(new_n596), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n335), .A2(new_n673), .A3(new_n710), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n334), .A2(new_n304), .A3(new_n298), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(new_n673), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n710), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n729), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n728), .A2(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT111), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n198), .ZN(G33));
  INV_X1    g550(.A(new_n647), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n335), .A2(new_n673), .A3(new_n737), .A4(new_n727), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  INV_X1    g553(.A(new_n726), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n619), .A2(new_n620), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n539), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT43), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n633), .A3(new_n637), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT44), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n384), .A2(KEYINPUT45), .A3(new_n393), .ZN(new_n746));
  INV_X1    g560(.A(new_n396), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n394), .ZN(new_n748));
  OAI211_X1 g562(.A(G469), .B(new_n746), .C1(new_n748), .C2(KEYINPUT45), .ZN(new_n749));
  INV_X1    g563(.A(new_n400), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT46), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n398), .B2(new_n410), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n677), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n755), .A2(new_n756), .A3(new_n658), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT112), .B1(new_n754), .B2(new_n659), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n740), .B(new_n745), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  XNOR2_X1  g574(.A(new_n754), .B(KEYINPUT47), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n333), .B1(new_n305), .B2(new_n308), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n673), .A2(new_n726), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n710), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  NAND2_X1  g579(.A1(new_n653), .A2(new_n673), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n601), .B(new_n766), .C1(KEYINPUT49), .C2(new_n676), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n309), .A2(new_n656), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n676), .A2(KEYINPUT49), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n340), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n742), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n705), .A2(new_n673), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n743), .A2(new_n541), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n676), .A2(new_n339), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n740), .B(new_n774), .C1(new_n761), .C2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n773), .A2(new_n681), .A3(new_n740), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n713), .B1(new_n705), .B2(new_n637), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n681), .A2(new_n541), .A3(new_n740), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n768), .A3(new_n456), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n627), .A3(new_n741), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n653), .A2(new_n601), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n681), .A3(new_n772), .A4(new_n773), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT50), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT51), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n687), .A2(new_n710), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n779), .B2(new_n778), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n664), .A2(new_n597), .ZN(new_n792));
  INV_X1    g606(.A(new_n725), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n637), .A2(new_n709), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n768), .A2(new_n792), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n649), .A3(new_n670), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n670), .A2(new_n649), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n791), .A4(new_n795), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n682), .A2(new_n685), .A3(new_n688), .A4(new_n707), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n627), .A2(new_n498), .A3(new_n646), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n309), .B2(new_n334), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n740), .A2(new_n412), .A3(new_n637), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n762), .A2(new_n808), .A3(new_n803), .A4(new_n805), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n731), .A2(new_n733), .ZN(new_n814));
  INV_X1    g628(.A(new_n727), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n762), .A2(new_n815), .A3(new_n456), .A4(new_n668), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n816), .B2(KEYINPUT42), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n732), .B1(new_n714), .B2(new_n719), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n762), .A2(new_n815), .A3(new_n456), .A4(new_n647), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n639), .ZN(new_n821));
  INV_X1    g635(.A(new_n599), .ZN(new_n822));
  INV_X1    g636(.A(new_n602), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n627), .A2(new_n498), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(KEYINPUT113), .C1(new_n621), .C2(new_n627), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n667), .B2(KEYINPUT113), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n608), .A2(new_n824), .A3(new_n611), .A4(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n605), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n817), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n813), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT53), .B1(new_n801), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n732), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n779), .B2(new_n778), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n603), .B1(new_n309), .B2(new_n334), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n639), .B1(new_n835), .B2(new_n457), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n836), .A3(new_n738), .A4(new_n828), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n734), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n682), .A2(new_n685), .A3(new_n688), .A4(new_n707), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT114), .B1(new_n804), .B2(new_n806), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n810), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n838), .A2(new_n797), .A3(new_n842), .A4(new_n800), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n832), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n831), .A2(KEYINPUT53), .A3(new_n797), .A4(new_n800), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n797), .A2(new_n800), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n605), .A2(new_n821), .A3(new_n828), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(new_n819), .A3(new_n818), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n817), .A3(new_n802), .A4(new_n812), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n774), .A2(new_n687), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n782), .A2(new_n667), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(G952), .A3(new_n258), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n777), .A2(new_n731), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT48), .Z(new_n860));
  NOR4_X1   g674(.A1(new_n789), .A2(new_n855), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n771), .B1(new_n861), .B2(new_n862), .ZN(G75));
  XNOR2_X1  g677(.A(new_n569), .B(new_n574), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT116), .Z(new_n865));
  NAND2_X1  g679(.A1(new_n847), .A2(new_n852), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n323), .A3(new_n591), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT55), .ZN(new_n874));
  INV_X1    g688(.A(new_n865), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n540), .A2(G953), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT117), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n872), .A2(new_n877), .A3(new_n879), .ZN(G51));
  INV_X1    g694(.A(new_n879), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n402), .A2(new_n409), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n853), .B1(new_n847), .B2(new_n852), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n855), .B2(KEYINPUT118), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n400), .B(KEYINPUT57), .Z(new_n886));
  OAI21_X1  g700(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n866), .A2(new_n323), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(new_n749), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n881), .B1(new_n887), .B2(new_n889), .ZN(G54));
  INV_X1    g704(.A(new_n528), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .A4(new_n323), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n891), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n895));
  OAI221_X1 g709(.A(new_n879), .B1(new_n891), .B2(new_n892), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(G60));
  NAND2_X1  g711(.A1(new_n616), .A2(new_n617), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n846), .B2(new_n854), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n899), .B(new_n902), .C1(new_n904), .C2(new_n884), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n846), .B2(new_n854), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n906), .A2(KEYINPUT120), .A3(new_n899), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n847), .A2(new_n852), .A3(new_n853), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n909), .B2(new_n883), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n898), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n879), .B(new_n905), .C1(new_n907), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n866), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n635), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n879), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n446), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n920), .C1(KEYINPUT121), .C2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT121), .B(new_n879), .C1(new_n916), .C2(new_n917), .ZN(new_n923));
  INV_X1    g737(.A(new_n920), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT61), .B(new_n923), .C1(new_n924), .C2(new_n918), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n544), .B2(new_n571), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n839), .A2(new_n849), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n567), .B(new_n568), .C1(G898), .C2(new_n258), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  XNOR2_X1  g745(.A(new_n269), .B(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n519), .A2(new_n520), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT123), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n791), .A2(new_n649), .A3(new_n670), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n665), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n660), .A2(new_n726), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n335), .A2(new_n673), .A3(new_n827), .A4(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n940), .A2(new_n759), .A3(new_n764), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n943), .B2(new_n258), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n734), .A2(new_n819), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n792), .B(new_n731), .C1(new_n757), .C2(new_n758), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(new_n937), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n948), .A3(new_n759), .A4(new_n764), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n258), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n258), .A2(G900), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT124), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n944), .B1(new_n934), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(G900), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n342), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  INV_X1    g773(.A(new_n928), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n949), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT126), .B(new_n959), .C1(new_n949), .C2(new_n960), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n279), .A3(new_n329), .A4(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n959), .B1(new_n943), .B2(new_n960), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n881), .B1(new_n966), .B2(new_n654), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n330), .B(KEYINPUT127), .Z(new_n968));
  OAI211_X1 g782(.A(new_n866), .B(new_n959), .C1(new_n291), .C2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(G57));
endmodule


