//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n906, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943;
  INV_X1    g000(.A(G226gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(new_n208), .B2(new_n207), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT24), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT25), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(new_n208), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT64), .B(new_n205), .C1(new_n207), .C2(new_n208), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n216), .A2(KEYINPUT25), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n212), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G190gat), .Z(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(KEYINPUT66), .A3(new_n222), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n219), .B1(new_n227), .B2(KEYINPUT67), .ZN(new_n228));
  INV_X1    g027(.A(new_n226), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT66), .B1(new_n221), .B2(new_n222), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n212), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n214), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT28), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT26), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n205), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n239), .B(new_n211), .C1(new_n238), .C2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n204), .B1(new_n234), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n233), .ZN(new_n245));
  INV_X1    g044(.A(new_n214), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n243), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT29), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n244), .B1(new_n249), .B2(new_n204), .ZN(new_n250));
  XOR2_X1   g049(.A(G211gat), .B(G218gat), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT72), .ZN(new_n252));
  XNOR2_X1  g051(.A(G197gat), .B(G204gat), .ZN(new_n253));
  INV_X1    g052(.A(G211gat), .ZN(new_n254));
  INV_X1    g053(.A(G218gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(KEYINPUT22), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n252), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n234), .B2(new_n243), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n202), .B2(new_n203), .ZN(new_n265));
  INV_X1    g064(.A(new_n258), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n244), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n259), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n262), .B1(new_n259), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT73), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n262), .ZN(new_n273));
  INV_X1    g072(.A(new_n267), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n265), .B2(new_n244), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(new_n277), .C1(new_n269), .C2(new_n268), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n279));
  AOI22_X1  g078(.A1(new_n272), .A2(new_n278), .B1(new_n268), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G113gat), .ZN(new_n281));
  INV_X1    g080(.A(G120gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285));
  OAI221_X1 g084(.A(new_n283), .B1(new_n281), .B2(new_n282), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n247), .A2(new_n288), .A3(new_n248), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n284), .A2(new_n285), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n283), .B1(new_n281), .B2(new_n282), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(new_n287), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n234), .B2(new_n243), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G227gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(new_n203), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT34), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n297), .A3(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT32), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT33), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G15gat), .B(G43gat), .Z(new_n308));
  XNOR2_X1  g107(.A(G71gat), .B(G99gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n310), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n304), .B(KEYINPUT32), .C1(new_n306), .C2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n303), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n301), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n311), .A2(new_n313), .A3(new_n303), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n311), .A2(new_n313), .A3(new_n303), .ZN(new_n319));
  OAI22_X1  g118(.A1(new_n319), .A2(new_n314), .B1(new_n300), .B2(new_n301), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT2), .B1(new_n322), .B2(new_n323), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  XOR2_X1   g130(.A(G141gat), .B(G148gat), .Z(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT77), .B(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n336), .B2(new_n322), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n332), .C1(new_n324), .C2(new_n325), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n288), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n292), .A2(new_n287), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n292), .A2(new_n287), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n335), .B(new_n338), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n293), .B1(KEYINPUT3), .B2(new_n339), .ZN(new_n348));
  INV_X1    g147(.A(new_n339), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n346), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(KEYINPUT4), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n293), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n352), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT78), .B1(new_n352), .B2(new_n356), .ZN(new_n358));
  OAI211_X1 g157(.A(KEYINPUT5), .B(new_n347), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n352), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n353), .A2(KEYINPUT79), .A3(new_n355), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n343), .A2(new_n367), .A3(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n359), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  INV_X1    g173(.A(new_n363), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n347), .A2(KEYINPUT5), .ZN(new_n376));
  INV_X1    g175(.A(new_n358), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n352), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n379), .B2(new_n370), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n359), .A2(new_n381), .A3(new_n363), .A4(new_n371), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n373), .A2(new_n374), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n380), .A2(new_n374), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n266), .B1(new_n351), .B2(new_n263), .ZN(new_n386));
  INV_X1    g185(.A(new_n251), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n257), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n387), .B2(new_n257), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n349), .B1(new_n389), .B2(new_n350), .ZN(new_n390));
  INV_X1    g189(.A(G228gat), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n386), .A2(new_n390), .B1(new_n391), .B2(new_n203), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT81), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n386), .A2(new_n391), .A3(new_n203), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT82), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n350), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n258), .A2(KEYINPUT82), .A3(KEYINPUT29), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n339), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G22gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  MUX2_X1   g204(.A(new_n401), .B(new_n402), .S(new_n405), .Z(new_n406));
  XNOR2_X1  g205(.A(new_n400), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n280), .A2(new_n321), .A3(new_n385), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT35), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n268), .A2(new_n279), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n411), .B(new_n276), .C1(new_n269), .C2(new_n268), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n407), .B(new_n412), .C1(new_n318), .C2(new_n320), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n363), .B(KEYINPUT84), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n379), .B2(new_n370), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n373), .A2(new_n374), .A3(new_n382), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT35), .B1(new_n417), .B2(new_n384), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g219(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n321), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n318), .A2(new_n320), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n268), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT37), .B1(new_n274), .B2(new_n275), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n262), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n271), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n430), .B2(KEYINPUT38), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n276), .B1(new_n428), .B2(new_n262), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT38), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT87), .B(KEYINPUT37), .C1(new_n274), .C2(new_n275), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n432), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n431), .A2(new_n437), .A3(new_n384), .A4(new_n417), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n348), .A2(new_n351), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n366), .A2(new_n439), .A3(new_n368), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n346), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n440), .A2(new_n346), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT39), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT85), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n414), .B(new_n442), .C1(new_n443), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT40), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n416), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n447), .B2(new_n448), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n407), .B1(new_n453), .B2(new_n412), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n272), .A2(new_n278), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n385), .A2(new_n456), .A3(new_n411), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n407), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n425), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n420), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G134gat), .B(G162gat), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n467));
  OR2_X1    g266(.A1(G43gat), .A2(G50gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469));
  NAND2_X1  g268(.A1(G43gat), .A2(G50gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT89), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n470), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  INV_X1    g273(.A(G29gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(G36gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n475), .B2(KEYINPUT14), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(G29gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n468), .A2(new_n482), .A3(new_n469), .A4(new_n470), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n472), .A2(new_n474), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(new_n476), .C1(new_n480), .C2(new_n478), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n494));
  INV_X1    g293(.A(G92gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT8), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n497), .A2(KEYINPUT100), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT100), .B1(new_n497), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT101), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G99gat), .ZN(new_n506));
  INV_X1    g305(.A(G106gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT101), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n498), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n484), .A2(KEYINPUT17), .A3(new_n486), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT100), .ZN(new_n514));
  AND2_X1   g313(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n515), .A2(new_n516), .A3(G92gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n499), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n497), .A2(KEYINPUT100), .A3(new_n499), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n511), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n493), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n489), .A2(new_n512), .A3(new_n513), .A4(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n484), .A2(new_n486), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n512), .B2(new_n523), .ZN(new_n526));
  NAND3_X1  g325(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n526), .A2(KEYINPUT102), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT102), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n522), .B1(new_n521), .B2(new_n493), .ZN(new_n531));
  AOI211_X1 g330(.A(new_n492), .B(new_n511), .C1(new_n519), .C2(new_n520), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n487), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n530), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n524), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G190gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT102), .B1(new_n526), .B2(new_n528), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n530), .A3(new_n527), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G190gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n524), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n467), .B1(new_n542), .B2(new_n255), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n536), .A2(G218gat), .A3(new_n541), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n466), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n540), .B1(new_n539), .B2(new_n524), .ZN(new_n546));
  INV_X1    g345(.A(new_n524), .ZN(new_n547));
  AOI211_X1 g346(.A(G190gat), .B(new_n547), .C1(new_n537), .C2(new_n538), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n255), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(new_n544), .A3(KEYINPUT97), .A4(new_n466), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n464), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(G57gat), .A2(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G57gat), .A2(G64gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(G71gat), .ZN(new_n557));
  INV_X1    g356(.A(G78gat), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n557), .B(new_n558), .C1(KEYINPUT94), .C2(KEYINPUT9), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n555), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT94), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT92), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G71gat), .B2(G78gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n565), .A2(new_n567), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n553), .A3(new_n554), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n564), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G127gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G15gat), .B(G22gat), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(G1gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(G1gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT90), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n579), .B2(G1gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(G8gat), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(G8gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n580), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n570), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT93), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n591), .A2(new_n592), .B1(new_n563), .B2(new_n560), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n589), .B1(KEYINPUT21), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n578), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n595), .B(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n549), .A2(new_n544), .A3(KEYINPUT97), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n465), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n463), .A3(new_n550), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n593), .B1(new_n531), .B2(new_n532), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n512), .A2(new_n573), .A3(new_n523), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(KEYINPUT10), .B(new_n593), .C1(new_n531), .C2(new_n532), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n605), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n614), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n552), .A2(new_n600), .A3(new_n603), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n583), .B(new_n587), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n513), .A3(new_n489), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n589), .A2(new_n487), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT18), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n626), .A2(KEYINPUT18), .A3(new_n627), .A4(new_n628), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n525), .A2(new_n588), .A3(new_n586), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n627), .B(KEYINPUT13), .Z(new_n635));
  AOI21_X1  g434(.A(KEYINPUT91), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT91), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  AOI211_X1 g437(.A(new_n637), .B(new_n638), .C1(new_n628), .C2(new_n633), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n631), .B(new_n632), .C1(new_n636), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G197gat), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT11), .B(G169gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n640), .A2(KEYINPUT88), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n640), .B2(KEYINPUT88), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n624), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n460), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n385), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT104), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(G1gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  NAND3_X1  g455(.A1(new_n460), .A2(new_n412), .A3(new_n651), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(G8gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n425), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n652), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n321), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n652), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n652), .A2(new_n408), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  AND3_X1   g471(.A1(new_n602), .A2(new_n463), .A3(new_n550), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n463), .B1(new_n602), .B2(new_n550), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n420), .B2(new_n459), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n600), .A2(new_n650), .A3(new_n622), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(G29gat), .A3(new_n385), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT45), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  INV_X1    g480(.A(new_n675), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n425), .A2(new_n455), .A3(new_n458), .ZN(new_n683));
  AOI22_X1  g482(.A1(KEYINPUT35), .A2(new_n409), .B1(new_n413), .B2(new_n418), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n681), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT44), .B1(new_n676), .B2(new_n681), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n677), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n385), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n680), .A2(new_n691), .ZN(G1328gat));
  NAND2_X1  g491(.A1(new_n685), .A2(new_n686), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n681), .A3(KEYINPUT44), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n412), .A4(new_n677), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n477), .B1(new_n695), .B2(KEYINPUT107), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n689), .A2(new_n697), .A3(new_n412), .A4(new_n677), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n412), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n678), .A2(G36gat), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n690), .B2(new_n425), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n678), .A2(G43gat), .A3(new_n667), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n689), .A2(new_n664), .A3(new_n677), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(G43gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(KEYINPUT47), .B2(new_n713), .ZN(G1330gat));
  NOR3_X1   g513(.A1(new_n678), .A2(G50gat), .A3(new_n408), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n407), .A3(new_n677), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(G50gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g517(.A(new_n594), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n578), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n578), .A2(new_n719), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n599), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n599), .B1(new_n720), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n673), .A2(new_n674), .A3(new_n724), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n460), .A2(new_n650), .A3(new_n725), .A4(new_n622), .ZN(new_n726));
  INV_X1    g525(.A(new_n385), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n412), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT49), .B(G64gat), .Z(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n730), .B2(new_n732), .ZN(G1333gat));
  AOI21_X1  g532(.A(new_n557), .B1(new_n726), .B2(new_n664), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n667), .A2(G71gat), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g536(.A1(new_n726), .A2(new_n407), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n600), .A2(new_n649), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n622), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT109), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n693), .A2(new_n694), .A3(new_n742), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n743), .A2(new_n727), .B1(new_n494), .B2(new_n496), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n682), .B(new_n740), .C1(new_n683), .C2(new_n684), .ZN(new_n745));
  NAND2_X1  g544(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n676), .A2(new_n740), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n622), .A3(new_n751), .ZN(new_n752));
  NOR4_X1   g551(.A1(new_n752), .A2(new_n385), .A3(new_n516), .A4(new_n515), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n744), .A2(new_n753), .ZN(G1336gat));
  NAND4_X1  g553(.A1(new_n693), .A2(new_n694), .A3(new_n412), .A4(new_n742), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G92gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n758), .A3(G92gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n700), .A2(G92gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n748), .A2(new_n751), .A3(new_n622), .A4(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n757), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n756), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n764), .B2(new_n756), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n762), .A2(new_n763), .B1(new_n766), .B2(new_n767), .ZN(G1337gat));
  OR2_X1    g567(.A1(new_n752), .A2(new_n667), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n665), .A2(new_n506), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n769), .A2(new_n506), .B1(new_n743), .B2(new_n770), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n751), .A3(new_n407), .A4(new_n622), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n507), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n408), .A2(new_n507), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n693), .A2(new_n694), .A3(new_n742), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n776), .A2(KEYINPUT114), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT114), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n743), .A2(new_n774), .B1(new_n772), .B2(new_n507), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(KEYINPUT53), .ZN(new_n782));
  AND4_X1   g581(.A1(new_n780), .A2(new_n773), .A3(KEYINPUT53), .A4(new_n775), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n778), .A2(new_n779), .B1(new_n782), .B2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n725), .A2(new_n785), .A3(new_n650), .A4(new_n623), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT115), .B1(new_n624), .B2(new_n649), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n611), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n609), .A2(new_n610), .A3(new_n605), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n792));
  AOI211_X1 g591(.A(KEYINPUT117), .B(new_n618), .C1(new_n611), .C2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n609), .A2(new_n610), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n604), .A3(new_n792), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n619), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n791), .B(KEYINPUT55), .C1(new_n793), .C2(new_n797), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n800), .A2(new_n649), .A3(new_n621), .A4(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n640), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n645), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n634), .A2(new_n635), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n644), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n622), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n603), .A3(new_n552), .ZN(new_n810));
  INV_X1    g609(.A(new_n792), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n605), .B(new_n811), .C1(new_n609), .C2(new_n610), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT117), .B1(new_n812), .B2(new_n618), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n794), .A3(new_n619), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n813), .A2(new_n814), .B1(new_n790), .B2(new_n789), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n621), .B1(new_n815), .B2(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(new_n801), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n804), .A2(new_n807), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n673), .B2(new_n674), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n810), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n786), .A2(new_n787), .B1(new_n821), .B2(new_n724), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n727), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n413), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n650), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n649), .A2(new_n281), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT118), .Z(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n826), .B2(new_n829), .ZN(G1340gat));
  NOR2_X1   g629(.A1(new_n826), .A2(new_n623), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(new_n282), .ZN(G1341gat));
  INV_X1    g631(.A(new_n826), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n600), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n682), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n836), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT56), .B1(new_n836), .B2(G134gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(G134gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(G1343gat));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n809), .A2(new_n841), .A3(new_n603), .A4(new_n552), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n724), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n810), .A2(KEYINPUT120), .A3(new_n820), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n843), .A2(new_n844), .B1(new_n786), .B2(new_n787), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n407), .A2(KEYINPUT57), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT121), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n724), .A3(new_n842), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n786), .A2(new_n787), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  INV_X1    g650(.A(new_n846), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n822), .B2(new_n408), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n847), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n385), .B(new_n412), .C1(new_n422), .C2(new_n424), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n649), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G141gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n700), .A2(new_n407), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n824), .A2(new_n664), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(G141gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n649), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT122), .Z(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n862), .B1(new_n858), .B2(KEYINPUT123), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n872), .A3(new_n649), .A4(new_n857), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT124), .B(new_n870), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n858), .A2(KEYINPUT123), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(G141gat), .A3(new_n873), .ZN(new_n877));
  INV_X1    g676(.A(new_n870), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n868), .B1(new_n874), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(new_n861), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n881), .A2(G148gat), .A3(new_n623), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n624), .A2(KEYINPUT125), .A3(new_n649), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n724), .B2(new_n821), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT125), .B1(new_n624), .B2(new_n649), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n408), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n823), .A2(new_n407), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n887), .A2(KEYINPUT57), .B1(new_n888), .B2(new_n854), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n622), .A3(new_n857), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n883), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n856), .A2(new_n622), .A3(new_n857), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(new_n883), .A3(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n882), .B1(new_n891), .B2(new_n893), .ZN(G1345gat));
  NAND3_X1  g693(.A1(new_n861), .A2(new_n322), .A3(new_n600), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n856), .A2(new_n600), .A3(new_n857), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n322), .ZN(G1346gat));
  OAI21_X1  g696(.A(new_n336), .B1(new_n881), .B2(new_n675), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n675), .A2(new_n336), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n856), .A2(new_n857), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n385), .A2(new_n412), .ZN(new_n902));
  NOR4_X1   g701(.A1(new_n822), .A2(new_n667), .A3(new_n407), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n649), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n622), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n600), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n222), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n235), .B2(new_n908), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n903), .A2(new_n682), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(G190gat), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT126), .B(new_n540), .C1(new_n903), .C2(new_n682), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n918));
  INV_X1    g717(.A(new_n221), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n913), .ZN(G1351gat));
  INV_X1    g719(.A(new_n888), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n664), .A2(new_n902), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n923), .A2(G197gat), .A3(new_n650), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n889), .A2(new_n649), .A3(new_n922), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G197gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(G1352gat));
  NOR3_X1   g729(.A1(new_n923), .A2(G204gat), .A3(new_n623), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT62), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n889), .A2(new_n622), .A3(new_n922), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G204gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  INV_X1    g734(.A(new_n923), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n254), .A3(new_n600), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n889), .A2(new_n600), .A3(new_n922), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n255), .A3(new_n682), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n889), .A2(new_n682), .A3(new_n922), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n255), .ZN(G1355gat));
endmodule


