//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT91), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G214), .A3(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT91), .B(G143), .ZN(new_n191));
  INV_X1    g005(.A(G214), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(G237), .A3(G953), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT18), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(KEYINPUT18), .A3(G131), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT64), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT64), .A2(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(new_n204), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n198), .A2(new_n199), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n210), .A2(new_n188), .B1(new_n189), .B2(G214), .ZN(new_n211));
  INV_X1    g025(.A(G237), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G214), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n209), .A2(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT92), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n194), .A2(KEYINPUT92), .A3(G131), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n219), .A2(new_n220), .B1(new_n195), .B2(new_n197), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n222));
  INV_X1    g036(.A(G125), .ZN(new_n223));
  OR3_X1    g037(.A1(new_n223), .A2(KEYINPUT16), .A3(G140), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(G146), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n204), .B(KEYINPUT19), .Z(new_n226));
  OR2_X1    g040(.A1(KEYINPUT64), .A2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n200), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n208), .B1(new_n221), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G113), .B(G122), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n231), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n225), .ZN(new_n240));
  AOI21_X1  g054(.A(G146), .B1(new_n222), .B2(new_n224), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT94), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n187), .A2(KEYINPUT91), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n214), .B1(new_n244), .B2(new_n215), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n218), .B(new_n197), .C1(new_n245), .C2(new_n190), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT92), .B1(new_n194), .B2(G131), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n243), .B1(new_n248), .B2(KEYINPUT17), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n219), .A2(new_n243), .A3(KEYINPUT17), .A4(new_n220), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT95), .B(new_n242), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT17), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n221), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n242), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n219), .A2(KEYINPUT17), .A3(new_n220), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT94), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n258), .B2(new_n250), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT95), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n235), .B(new_n208), .C1(new_n255), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT96), .ZN(new_n262));
  INV_X1    g076(.A(new_n208), .ZN(new_n263));
  INV_X1    g077(.A(new_n254), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n259), .B2(KEYINPUT95), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n242), .B1(new_n249), .B2(new_n251), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT95), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT96), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n235), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n239), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G475), .A2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n272), .A2(KEYINPUT20), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n272), .A2(KEYINPUT97), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT97), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n278), .B(new_n239), .C1(new_n262), .C2(new_n271), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n277), .A2(new_n279), .A3(new_n274), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT99), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT98), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n269), .A2(new_n235), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n262), .B2(new_n271), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(G902), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n269), .A2(new_n235), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n261), .A2(KEYINPUT96), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n270), .B1(new_n269), .B2(new_n235), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT98), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n293), .A3(G475), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n282), .A2(new_n283), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n292), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT12), .ZN(new_n298));
  INV_X1    g112(.A(G101), .ZN(new_n299));
  INV_X1    g113(.A(G107), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G104), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n234), .A2(G107), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n300), .A2(G104), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT84), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n234), .A2(G107), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n306), .A2(KEYINPUT84), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n304), .B1(new_n314), .B2(G101), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n302), .B1(new_n309), .B2(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n301), .B1(new_n307), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT85), .A3(new_n299), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n303), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n227), .A2(G143), .A3(new_n200), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n206), .A2(G143), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G128), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT1), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(new_n203), .B2(G143), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n187), .A2(G146), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n325), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT86), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n321), .A2(KEYINPUT86), .A3(new_n332), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n201), .A2(new_n202), .A3(new_n187), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n338));
  OAI21_X1  g152(.A(G128), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n330), .B1(new_n203), .B2(G143), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n339), .A2(new_n340), .B1(new_n328), .B2(new_n326), .ZN(new_n341));
  INV_X1    g155(.A(new_n303), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT85), .B1(new_n319), .B2(new_n299), .ZN(new_n343));
  NOR4_X1   g157(.A1(new_n316), .A2(new_n318), .A3(new_n304), .A4(G101), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n335), .A2(new_n336), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G137), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT11), .B1(new_n347), .B2(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(G134), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(KEYINPUT65), .A2(G137), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT65), .A2(G137), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT11), .A2(G134), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n350), .A2(new_n354), .A3(new_n197), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n197), .B1(new_n350), .B2(new_n354), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n298), .B1(new_n346), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n336), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT86), .B1(new_n321), .B2(new_n332), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n325), .B1(new_n322), .B2(KEYINPUT1), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n329), .B1(new_n228), .B2(new_n187), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n327), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI22_X1  g177(.A1(new_n359), .A2(new_n360), .B1(new_n363), .B2(new_n321), .ZN(new_n364));
  INV_X1    g178(.A(new_n357), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(KEYINPUT12), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT83), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n213), .A2(G227), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n359), .B2(new_n360), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n345), .A2(KEYINPUT87), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n321), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT10), .A4(new_n363), .ZN(new_n378));
  OAI221_X1 g192(.A(KEYINPUT4), .B1(new_n299), .B2(new_n319), .C1(new_n343), .C2(new_n344), .ZN(new_n379));
  AND2_X1   g193(.A1(KEYINPUT0), .A2(G128), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT0), .A2(G128), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G143), .B1(new_n227), .B2(new_n200), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(new_n329), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n322), .A2(new_n380), .A3(new_n324), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OR3_X1    g200(.A1(new_n319), .A2(KEYINPUT4), .A3(new_n299), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n357), .B(KEYINPUT88), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n374), .A2(new_n378), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n367), .A2(new_n372), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n378), .A2(new_n388), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT10), .B1(new_n335), .B2(new_n336), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n365), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n390), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n371), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n297), .B1(new_n397), .B2(new_n296), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n390), .A3(new_n372), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n367), .A2(new_n390), .ZN(new_n400));
  OAI211_X1 g214(.A(G469), .B(new_n399), .C1(new_n400), .C2(new_n372), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  OAI21_X1  g217(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G214), .B1(G237), .B2(G902), .ZN(new_n406));
  OAI21_X1  g220(.A(G210), .B1(G237), .B2(G902), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n341), .A2(new_n223), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n223), .B2(new_n386), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n213), .A2(G224), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g225(.A(G119), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G116), .ZN(new_n413));
  OAI21_X1  g227(.A(G113), .B1(new_n413), .B2(KEYINPUT5), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n415));
  INV_X1    g229(.A(G116), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G119), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n412), .A2(G116), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(G119), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n420), .A3(KEYINPUT67), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n414), .B1(new_n422), .B2(KEYINPUT5), .ZN(new_n423));
  XNOR2_X1  g237(.A(G116), .B(G119), .ZN(new_n424));
  OR2_X1    g238(.A1(KEYINPUT2), .A2(G113), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n426));
  AND3_X1   g240(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n375), .A2(new_n377), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n425), .B1(new_n427), .B2(new_n426), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(new_n432), .A3(new_n421), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n428), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n379), .A2(new_n434), .A3(new_n387), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G122), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n431), .A2(new_n435), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(KEYINPUT89), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n437), .A2(KEYINPUT6), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n411), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT90), .B(new_n411), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n436), .B(KEYINPUT8), .Z(new_n447));
  AND2_X1   g261(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n428), .B1(new_n448), .B2(new_n414), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n321), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n345), .A2(new_n430), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n410), .A2(KEYINPUT7), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n409), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n409), .A2(new_n453), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n456), .B2(new_n437), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n407), .B1(new_n446), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n407), .ZN(new_n459));
  INV_X1    g273(.A(new_n457), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n459), .B(new_n460), .C1(new_n444), .C2(new_n445), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n406), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n405), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n238), .B1(new_n289), .B2(new_n290), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n278), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n272), .A2(KEYINPUT97), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n273), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n275), .B1(new_n467), .B2(KEYINPUT20), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n287), .A2(new_n293), .A3(G475), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT99), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n187), .A2(G128), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT100), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(new_n325), .B2(G143), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n473), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G134), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n416), .A2(G122), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(G116), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n481), .A3(new_n300), .ZN(new_n482));
  OAI21_X1  g296(.A(G107), .B1(new_n477), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n472), .B1(G128), .B2(new_n187), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n476), .B(new_n484), .C1(G134), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(G134), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(KEYINPUT14), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT101), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n478), .B1(new_n481), .B2(KEYINPUT14), .ZN(new_n490));
  OAI21_X1  g304(.A(G107), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n482), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G217), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n403), .A2(new_n494), .A3(G953), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n493), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n292), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT102), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(G478), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n497), .B(new_n292), .C1(KEYINPUT15), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(G234), .A2(G237), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n505), .A2(G952), .A3(new_n213), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n505), .A2(G902), .A3(G953), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n295), .A2(new_n463), .A3(new_n470), .A4(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n512));
  INV_X1    g326(.A(G134), .ZN(new_n513));
  INV_X1    g327(.A(new_n352), .ZN(new_n514));
  NOR2_X1   g328(.A1(KEYINPUT65), .A2(G137), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n197), .B1(new_n516), .B2(new_n349), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n355), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n363), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n385), .B(new_n384), .C1(new_n355), .C2(new_n356), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n434), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n189), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT27), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT69), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n350), .A2(new_n354), .A3(new_n197), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n516), .A2(new_n349), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n197), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n521), .B1(new_n341), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n434), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n433), .A2(KEYINPUT68), .A3(new_n428), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n529), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n433), .A2(KEYINPUT68), .A3(new_n428), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT68), .B1(new_n433), .B2(new_n428), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n541), .A2(KEYINPUT69), .A3(new_n521), .A4(new_n519), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n524), .A2(new_n528), .A3(new_n538), .A4(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n538), .A2(new_n542), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n528), .A4(new_n524), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n533), .A2(new_n434), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n538), .A2(new_n542), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT28), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n533), .A2(new_n537), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n528), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n557), .A3(KEYINPUT70), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT32), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n560), .A2(new_n565), .A3(new_n561), .A4(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G472), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n551), .A2(new_n528), .A3(new_n554), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n524), .A2(new_n538), .A3(new_n542), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n556), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n569), .A2(KEYINPUT71), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n533), .A2(new_n537), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n533), .A2(new_n537), .A3(KEYINPUT72), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n538), .A3(new_n542), .A4(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n553), .B1(new_n578), .B2(KEYINPUT28), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n556), .A2(new_n572), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n569), .A2(new_n572), .A3(new_n571), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT71), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n568), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n512), .B1(new_n567), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(KEYINPUT73), .B(new_n586), .C1(new_n564), .C2(new_n566), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n325), .A2(G119), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n325), .A2(G119), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT23), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT77), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n596));
  OAI211_X1 g410(.A(G119), .B(new_n325), .C1(new_n596), .C2(KEYINPUT23), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G110), .ZN(new_n600));
  OAI22_X1  g414(.A1(new_n240), .A2(new_n241), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT24), .B(G110), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n603), .A2(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(KEYINPUT75), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n592), .A2(KEYINPUT74), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n592), .A2(KEYINPUT74), .ZN(new_n608));
  INV_X1    g422(.A(new_n593), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n607), .A2(new_n609), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n614), .A2(new_n604), .A3(new_n605), .A4(new_n608), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(KEYINPUT76), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n602), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n225), .A2(new_n205), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n606), .A2(new_n610), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n599), .A2(new_n600), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT78), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT22), .B(G137), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n617), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT79), .ZN(new_n629));
  INV_X1    g443(.A(new_n624), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(new_n625), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n625), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n626), .A2(KEYINPUT79), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n611), .A2(new_n612), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n615), .A2(KEYINPUT76), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n601), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n635), .B1(new_n638), .B2(new_n621), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n628), .A2(new_n639), .A3(new_n292), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT25), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n628), .A2(new_n639), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n494), .B1(G234), .B2(new_n292), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT80), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT80), .ZN(new_n647));
  INV_X1    g461(.A(new_n645), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n647), .B(new_n648), .C1(new_n642), .C2(new_n643), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n628), .A2(new_n639), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n292), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n591), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n654), .ZN(new_n656));
  NOR4_X1   g470(.A1(new_n646), .A2(new_n649), .A3(new_n656), .A4(KEYINPUT82), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n590), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n511), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n299), .ZN(G3));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n662));
  INV_X1    g476(.A(new_n497), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(KEYINPUT33), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT33), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n497), .A2(KEYINPUT103), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT104), .B1(new_n486), .B2(new_n492), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n665), .B1(new_n667), .B2(new_n496), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n496), .B2(new_n667), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n664), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(G478), .A3(new_n292), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n499), .A2(new_n502), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n295), .B2(new_n470), .ZN(new_n675));
  INV_X1    g489(.A(new_n404), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n398), .B2(new_n401), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n560), .A2(new_n292), .A3(new_n562), .ZN(new_n678));
  INV_X1    g492(.A(new_n562), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT70), .B1(new_n548), .B2(new_n557), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(G472), .A2(new_n678), .B1(new_n681), .B2(new_n561), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n677), .A2(new_n658), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n509), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n406), .B(new_n684), .C1(new_n458), .C2(new_n461), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n675), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT34), .B(G104), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G6));
  NOR2_X1   g503(.A1(new_n277), .A2(new_n279), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n281), .A3(new_n273), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n467), .A2(KEYINPUT20), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n469), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n685), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n504), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n683), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT35), .B(G107), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NOR2_X1   g512(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n617), .A2(new_n622), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n653), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n650), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n682), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n511), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT105), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G12));
  AND3_X1   g522(.A1(new_n590), .A2(new_n463), .A3(new_n703), .ZN(new_n709));
  INV_X1    g523(.A(G900), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n507), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n506), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n693), .A2(new_n504), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  NAND2_X1  g531(.A1(new_n295), .A2(new_n470), .ZN(new_n718));
  INV_X1    g532(.A(new_n703), .ZN(new_n719));
  INV_X1    g533(.A(new_n504), .ZN(new_n720));
  INV_X1    g534(.A(new_n406), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n723), .A2(KEYINPUT108), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(KEYINPUT108), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n713), .B(KEYINPUT39), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n677), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT40), .Z(new_n728));
  AOI21_X1  g542(.A(new_n460), .B1(new_n444), .B2(new_n445), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n407), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n578), .A2(KEYINPUT107), .A3(new_n556), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n543), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT107), .B1(new_n578), .B2(new_n556), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n292), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G472), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n567), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n724), .A2(new_n725), .A3(new_n728), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G143), .ZN(G45));
  AOI21_X1  g555(.A(new_n283), .B1(new_n282), .B2(new_n294), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n468), .A2(KEYINPUT99), .A3(new_n469), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n673), .B(new_n713), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n675), .A2(KEYINPUT109), .A3(new_n713), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n709), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n397), .A2(new_n296), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n397), .A2(new_n296), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n404), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n590), .A2(new_n658), .A3(new_n694), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n673), .B1(new_n742), .B2(new_n743), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n750), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n658), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n588), .A2(new_n589), .A3(new_n758), .A4(new_n753), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(KEYINPUT110), .A3(new_n675), .A4(new_n694), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT41), .B(G113), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G15));
  NAND2_X1  g577(.A1(new_n567), .A2(new_n587), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT73), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n567), .A2(new_n512), .A3(new_n587), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n658), .A4(new_n754), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n695), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n416), .ZN(G18));
  NOR2_X1   g583(.A1(new_n462), .A2(new_n753), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n765), .A2(new_n770), .A3(new_n766), .A4(new_n703), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n295), .A2(new_n470), .A3(new_n510), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n412), .ZN(G21));
  NAND2_X1  g588(.A1(new_n650), .A2(new_n654), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n548), .B1(new_n528), .B2(new_n579), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n561), .ZN(new_n778));
  INV_X1    g592(.A(new_n678), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT111), .B(G472), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n776), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n753), .A3(new_n509), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n718), .A2(new_n782), .A3(new_n730), .A4(new_n722), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT112), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G122), .ZN(G24));
  OAI211_X1 g599(.A(new_n703), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT113), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n746), .A2(new_n747), .A3(new_n770), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G125), .ZN(G27));
  NOR3_X1   g603(.A1(new_n405), .A2(new_n730), .A3(new_n721), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n590), .A2(new_n790), .A3(new_n658), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n746), .A2(new_n747), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n775), .B1(new_n567), .B2(new_n587), .ZN(new_n796));
  INV_X1    g610(.A(new_n790), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n746), .A2(new_n747), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  NAND2_X1  g615(.A1(new_n765), .A2(new_n766), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n758), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n715), .A3(KEYINPUT114), .A4(new_n790), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n791), .B2(new_n714), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n513), .ZN(G36));
  NOR2_X1   g622(.A1(new_n742), .A2(new_n743), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT43), .A3(new_n673), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n718), .B2(new_n674), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n682), .B(new_n719), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT44), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n730), .A2(new_n721), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n810), .A2(new_n812), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n682), .A2(new_n719), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT45), .B(new_n399), .C1(new_n400), .C2(new_n372), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n372), .B1(new_n367), .B2(new_n390), .ZN(new_n826));
  INV_X1    g640(.A(new_n399), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(G469), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n297), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(KEYINPUT46), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(KEYINPUT115), .A3(new_n752), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(KEYINPUT46), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n831), .B2(new_n752), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n404), .B(new_n726), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n814), .A2(KEYINPUT116), .A3(new_n815), .A4(new_n820), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n823), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G137), .ZN(G39));
  OAI21_X1  g654(.A(new_n404), .B1(new_n834), .B2(new_n835), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT47), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n746), .A2(new_n747), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n802), .A2(new_n758), .A3(new_n815), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(G140), .Z(G42));
  NAND2_X1  g660(.A1(new_n751), .A2(new_n752), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT117), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT49), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n776), .A2(new_n406), .A3(new_n404), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n732), .A2(new_n738), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n809), .A3(new_n673), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n718), .A2(new_n730), .A3(new_n722), .ZN(new_n854));
  INV_X1    g668(.A(new_n713), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n703), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT119), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n405), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n738), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n788), .A2(new_n748), .A3(new_n716), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT52), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n807), .B1(new_n795), .B2(new_n799), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n772), .A2(new_n771), .B1(new_n767), .B2(new_n695), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n295), .A2(new_n686), .A3(new_n470), .A4(new_n504), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n511), .B1(new_n659), .B2(new_n704), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n756), .A2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n675), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n686), .A3(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n761), .A2(new_n865), .A3(new_n867), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n746), .A2(new_n747), .A3(new_n787), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n504), .A2(new_n855), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n590), .A2(new_n693), .A3(new_n703), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n790), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n862), .A2(new_n872), .A3(new_n784), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n853), .B1(new_n861), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n748), .A2(new_n859), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n716), .A4(new_n788), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n860), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n866), .A2(new_n863), .A3(new_n864), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n784), .A3(new_n761), .A4(new_n871), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n797), .B1(new_n873), .B2(new_n875), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n884), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT54), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n712), .B1(new_n810), .B2(new_n812), .ZN(new_n892));
  NOR4_X1   g706(.A1(new_n732), .A2(new_n406), .A3(new_n753), .A4(new_n781), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT50), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n815), .A2(new_n754), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n712), .B(new_n896), .C1(new_n810), .C2(new_n812), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n787), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n896), .A2(new_n738), .A3(new_n758), .A4(new_n712), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n809), .A3(new_n674), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n781), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n842), .B1(new_n404), .B2(new_n848), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n815), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n895), .B(new_n901), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n892), .A2(new_n770), .A3(new_n902), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n899), .A2(new_n675), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT120), .B1(new_n213), .B2(G952), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(KEYINPUT120), .B2(new_n213), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n897), .A2(new_n796), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT48), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n917), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(KEYINPUT121), .B2(new_n916), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n909), .B(new_n914), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n891), .A2(new_n908), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(G952), .A2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n852), .B1(new_n922), .B2(new_n923), .ZN(G75));
  NOR2_X1   g738(.A1(new_n440), .A2(new_n441), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n411), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n292), .B1(new_n879), .B2(new_n889), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(KEYINPUT56), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n213), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n931), .A2(KEYINPUT56), .A3(new_n929), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G51));
  XNOR2_X1  g751(.A(new_n297), .B(KEYINPUT57), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n891), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n391), .A2(new_n396), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n930), .A2(G469), .A3(new_n824), .A4(new_n828), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(G54));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n944));
  AND2_X1   g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n930), .A2(new_n690), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n690), .B1(new_n930), .B2(new_n945), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n934), .B(new_n946), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n890), .A2(G902), .A3(new_n945), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n690), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n944), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT123), .B1(new_n950), .B2(new_n690), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n933), .B1(new_n950), .B2(new_n690), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n947), .A2(new_n948), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT124), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(G60));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT59), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n891), .A2(new_n670), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n670), .B1(new_n891), .B2(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n933), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT60), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n879), .B2(new_n889), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n701), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n934), .C1(new_n651), .C2(new_n965), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G66));
  INV_X1    g783(.A(G224), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n508), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n886), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n925), .B1(G898), .B2(new_n213), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT125), .Z(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  AND3_X1   g790(.A1(new_n788), .A2(new_n716), .A3(new_n748), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n740), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT62), .Z(new_n979));
  NAND2_X1  g793(.A1(new_n868), .A2(new_n870), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n718), .B2(new_n720), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n792), .A2(new_n726), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n845), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n839), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n213), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n522), .A2(new_n523), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(new_n226), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n837), .A2(new_n854), .A3(new_n796), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n845), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n991), .A2(new_n862), .A3(new_n977), .ZN(new_n992));
  AOI21_X1  g806(.A(G953), .B1(new_n992), .B2(new_n839), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n213), .A2(G900), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n987), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n993), .A2(new_n989), .A3(new_n994), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n988), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n213), .B1(G227), .B2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n988), .B(new_n1002), .C1(new_n997), .C2(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G72));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n984), .B2(new_n886), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n528), .A3(new_n570), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n992), .A2(new_n839), .A3(new_n972), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n1006), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n570), .A2(new_n528), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n933), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n571), .A2(new_n543), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n890), .A2(new_n1006), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(G57));
endmodule


