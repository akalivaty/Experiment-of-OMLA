//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(new_n203), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR3_X1   g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT66), .B(G238), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT67), .B(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n203), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n211), .A2(new_n216), .A3(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  AOI22_X1  g0045(.A1(new_n245), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n214), .A2(G33), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n255));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  OR3_X1    g0058(.A1(new_n258), .A2(KEYINPUT12), .A3(G68), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT12), .B1(new_n258), .B2(G68), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n256), .A2(new_n214), .A3(G1), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n252), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n214), .A2(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n203), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n259), .A2(new_n260), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n254), .A2(new_n255), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G226), .A2(G1698), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n229), .B2(G1698), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT72), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n274), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n270), .A2(new_n271), .B1(G33), .B2(G97), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT72), .B1(new_n280), .B2(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  INV_X1    g0083(.A(new_n215), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n276), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G238), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n277), .A2(new_n287), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n268), .B1(new_n282), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g0094(.A(KEYINPUT13), .B(new_n292), .C1(new_n279), .C2(new_n281), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n298));
  OAI211_X1 g0098(.A(G169), .B(new_n298), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n282), .A2(new_n293), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT13), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n282), .A2(new_n268), .A3(new_n293), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n298), .B1(new_n304), .B2(G169), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n267), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(G200), .B1(new_n294), .B2(new_n295), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n266), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT74), .ZN(new_n311));
  INV_X1    g0111(.A(new_n262), .ZN(new_n312));
  INV_X1    g0112(.A(new_n263), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G50), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n312), .A2(new_n314), .B1(G50), .B2(new_n258), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n204), .A2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(G150), .ZN(new_n317));
  INV_X1    g0117(.A(new_n245), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT8), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G58), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n316), .B1(new_n317), .B2(new_n318), .C1(new_n323), .C2(new_n248), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n315), .B1(new_n324), .B2(new_n252), .ZN(new_n325));
  INV_X1    g0125(.A(G226), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n289), .B1(new_n326), .B2(new_n291), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n271), .A2(G222), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n271), .A2(G1698), .ZN(new_n330));
  INV_X1    g0130(.A(G223), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n329), .B1(new_n218), .B2(new_n271), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n327), .B1(new_n332), .B2(new_n278), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G179), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n325), .B(new_n335), .C1(new_n336), .C2(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n324), .A2(new_n252), .ZN(new_n338));
  INV_X1    g0138(.A(new_n315), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n325), .A2(KEYINPUT71), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT71), .B1(new_n338), .B2(new_n339), .ZN(new_n346));
  AOI211_X1 g0146(.A(new_n341), .B(new_n315), .C1(new_n324), .C2(new_n252), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT9), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n333), .A2(G190), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n333), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT10), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n349), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n337), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n326), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n271), .B(new_n359), .C1(G223), .C2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n277), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n289), .B1(new_n229), .B2(new_n291), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n362), .A2(new_n363), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(G169), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT3), .A2(G33), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT3), .A2(G33), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT75), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n271), .B2(G20), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT7), .A4(new_n214), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT76), .B1(new_n202), .B2(new_n203), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(G58), .A3(G68), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n381), .A3(new_n212), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G20), .ZN(new_n383));
  INV_X1    g0183(.A(G159), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n318), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n203), .B1(new_n374), .B2(new_n371), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n252), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n322), .A2(new_n313), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n312), .B1(KEYINPUT77), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n261), .B2(new_n323), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n367), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n395), .ZN(new_n399));
  INV_X1    g0199(.A(new_n252), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n385), .B1(new_n377), .B2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n390), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT18), .B1(new_n403), .B2(new_n367), .ZN(new_n404));
  INV_X1    g0204(.A(G190), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n362), .A2(new_n363), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(G200), .B2(new_n366), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n391), .A2(new_n395), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n407), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n398), .A2(new_n404), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n214), .A2(new_n218), .B1(new_n414), .B2(new_n247), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n323), .A2(new_n318), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n252), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n263), .A2(new_n249), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n262), .A2(new_n418), .B1(new_n218), .B2(new_n261), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n289), .B1(new_n219), .B2(new_n291), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n271), .A2(G232), .A3(new_n328), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n423), .B2(new_n271), .C1(new_n330), .C2(new_n217), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n424), .B2(new_n278), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n420), .B1(new_n425), .B2(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT70), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT70), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n420), .C1(new_n425), .C2(G169), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n364), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(G190), .ZN(new_n432));
  INV_X1    g0232(.A(new_n420), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n351), .C2(new_n425), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n358), .A2(new_n413), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n311), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G264), .B(G1698), .C1(new_n368), .C2(new_n369), .ZN(new_n438));
  OAI211_X1 g0238(.A(G257), .B(new_n328), .C1(new_n368), .C2(new_n369), .ZN(new_n439));
  INV_X1    g0239(.A(G303), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n271), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n278), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n277), .A2(G274), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n443), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n286), .A2(G45), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(G41), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(new_n447), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n285), .A3(KEYINPUT79), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n278), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G270), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n442), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n261), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n286), .A2(G33), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n400), .A2(new_n258), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT78), .B(G97), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n214), .B(new_n468), .C1(new_n469), .C2(G33), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n251), .A2(new_n215), .B1(G20), .B2(new_n462), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT78), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G97), .ZN(new_n476));
  AOI21_X1  g0276(.A(G33), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n468), .A2(new_n214), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT20), .B(new_n471), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n467), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n461), .A2(new_n481), .A3(new_n482), .A4(G179), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n442), .A2(new_n458), .A3(G179), .A4(new_n460), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n400), .A2(new_n258), .A3(new_n465), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n463), .B1(new_n485), .B2(new_n462), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT20), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n477), .A2(new_n478), .ZN(new_n488));
  INV_X1    g0288(.A(new_n471), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n490), .B2(new_n479), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT82), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n442), .A2(new_n458), .A3(new_n460), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G169), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(G200), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n491), .C1(new_n405), .C2(new_n495), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n481), .A2(new_n495), .A3(KEYINPUT21), .A4(G169), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n493), .A2(new_n497), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n423), .A3(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n507));
  AND4_X1   g0307(.A1(new_n503), .A2(new_n504), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n214), .B(G87), .C1(new_n368), .C2(new_n369), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n271), .A2(new_n214), .A3(G87), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(KEYINPUT84), .B2(KEYINPUT24), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n508), .A2(new_n511), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n252), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT25), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n258), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n423), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n466), .A2(G107), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n271), .A2(G250), .A3(new_n328), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n278), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n459), .A2(G264), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n458), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G190), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n528), .A2(new_n278), .B1(G264), .B2(new_n459), .ZN(new_n533));
  AOI21_X1  g0333(.A(G200), .B1(new_n533), .B2(new_n458), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n520), .B(new_n524), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n336), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n364), .A3(new_n458), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n400), .B1(new_n516), .B2(new_n518), .ZN(new_n538));
  INV_X1    g0338(.A(new_n524), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n414), .A2(new_n261), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n469), .B2(new_n247), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G87), .A2(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n474), .A2(new_n476), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n214), .B1(new_n273), .B2(new_n542), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n271), .A2(new_n214), .A3(G68), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n541), .B1(new_n549), .B2(new_n252), .ZN(new_n550));
  XOR2_X1   g0350(.A(new_n414), .B(KEYINPUT80), .Z(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n466), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n277), .A2(G274), .A3(new_n446), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n277), .A2(G250), .A3(new_n452), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(G1698), .C1(new_n368), .C2(new_n369), .ZN(new_n556));
  OAI211_X1 g0356(.A(G238), .B(new_n328), .C1(new_n368), .C2(new_n369), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n278), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n550), .A2(new_n552), .B1(new_n560), .B2(new_n364), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n278), .ZN(new_n562));
  INV_X1    g0362(.A(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n336), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(G200), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(G190), .A3(new_n563), .ZN(new_n568));
  INV_X1    g0368(.A(G87), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT81), .B1(new_n485), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT81), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n262), .A2(new_n571), .A3(G87), .A4(new_n465), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(new_n550), .A3(new_n568), .A4(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n535), .A2(new_n540), .A3(new_n566), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n261), .A2(new_n473), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n485), .B2(new_n473), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  AND2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n423), .A2(KEYINPUT6), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n469), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(G20), .B1(G77), .B2(new_n245), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT7), .B1(new_n370), .B2(new_n214), .ZN(new_n585));
  NOR4_X1   g0385(.A1(new_n368), .A2(new_n369), .A3(new_n373), .A4(G20), .ZN(new_n586));
  OAI21_X1  g0386(.A(G107), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n577), .B1(new_n588), .B2(new_n252), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(new_n328), .C1(new_n368), .C2(new_n369), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n328), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n468), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n278), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n451), .A2(new_n457), .B1(new_n459), .B2(G257), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(G190), .ZN(new_n599));
  AOI21_X1  g0399(.A(G200), .B1(new_n596), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n589), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n589), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n336), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n596), .A2(new_n597), .A3(new_n364), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n575), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n437), .A2(new_n502), .A3(new_n607), .ZN(G372));
  NAND3_X1  g0408(.A1(new_n568), .A2(new_n550), .A3(new_n573), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT86), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n564), .B2(G200), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n564), .A2(new_n610), .A3(G200), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n564), .A2(new_n614), .A3(new_n336), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT85), .B1(new_n560), .B2(G169), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n612), .A2(new_n613), .B1(new_n561), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n605), .A3(new_n601), .A4(new_n535), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n493), .A2(new_n540), .A3(new_n497), .A4(new_n500), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n596), .A2(new_n597), .A3(new_n364), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n589), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(new_n603), .A3(new_n566), .A4(new_n574), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n617), .A2(new_n561), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n437), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n337), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n398), .A2(new_n404), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n306), .A2(new_n431), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n410), .A2(new_n411), .A3(new_n309), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n356), .B1(new_n349), .B2(new_n353), .ZN(new_n638));
  AOI211_X1 g0438(.A(KEYINPUT10), .B(new_n352), .C1(new_n345), .C2(new_n348), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n633), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n632), .A2(new_n642), .ZN(G369));
  AND2_X1   g0443(.A1(new_n497), .A2(new_n500), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n493), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n257), .A2(new_n214), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(G213), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n491), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT87), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n501), .B2(new_n653), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n535), .A2(new_n540), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n520), .B2(new_n524), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n540), .B2(new_n651), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n651), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n644), .B2(new_n493), .ZN(new_n662));
  INV_X1    g0462(.A(new_n657), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n540), .B2(new_n661), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n209), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n213), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n545), .A2(G116), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G1), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n619), .B2(new_n620), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n629), .B1(new_n627), .B2(KEYINPUT26), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n623), .B1(new_n618), .B2(new_n622), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n535), .A2(new_n601), .A3(new_n605), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n493), .A2(new_n540), .A3(new_n497), .A4(new_n500), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(KEYINPUT89), .A3(new_n683), .A4(new_n618), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT90), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n685), .A2(new_n686), .A3(new_n651), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n686), .B1(new_n685), .B2(new_n651), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT29), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n631), .A2(new_n651), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n607), .A2(new_n502), .A3(new_n651), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n495), .A2(new_n364), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n598), .A3(new_n531), .A4(new_n564), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n533), .A2(new_n560), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n696), .A2(new_n598), .A3(new_n484), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n695), .B1(KEYINPUT30), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(KEYINPUT30), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n661), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT31), .B(new_n661), .C1(new_n698), .C2(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n693), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n689), .A2(new_n692), .B1(G330), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n676), .B1(new_n705), .B2(G1), .ZN(G364));
  NOR2_X1   g0506(.A1(new_n256), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n286), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n669), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n209), .A2(G355), .A3(new_n271), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G116), .B2(new_n209), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n209), .A2(new_n370), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n445), .B2(new_n670), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n243), .A2(G45), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n215), .B1(G20), .B2(new_n336), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n710), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n405), .A2(G179), .A3(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n214), .ZN(new_n725));
  INV_X1    g0525(.A(G294), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n214), .A2(new_n364), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(KEYINPUT33), .A2(G317), .ZN(new_n732));
  NAND2_X1  g0532(.A1(KEYINPUT33), .A2(G317), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n729), .A2(new_n405), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n727), .B(new_n734), .C1(G326), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n728), .A2(G190), .A3(new_n351), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n271), .B1(new_n738), .B2(G322), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G190), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n214), .A2(G179), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n740), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G311), .A2(new_n742), .B1(new_n745), .B2(G329), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(new_n405), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT92), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n752), .A2(G283), .B1(G303), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n736), .A2(new_n739), .A3(new_n746), .A4(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n731), .A2(new_n203), .B1(new_n569), .B2(new_n753), .ZN(new_n757));
  INV_X1    g0557(.A(new_n735), .ZN(new_n758));
  INV_X1    g0558(.A(G50), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n745), .A2(G159), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(G107), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n271), .B1(new_n737), .B2(new_n202), .ZN(new_n764));
  INV_X1    g0564(.A(new_n218), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(new_n742), .ZN(new_n766));
  INV_X1    g0566(.A(new_n725), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n760), .A2(KEYINPUT32), .B1(new_n767), .B2(G97), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n762), .A2(new_n763), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n756), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n723), .B1(new_n770), .B2(new_n720), .ZN(new_n771));
  INV_X1    g0571(.A(new_n719), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n655), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n655), .A2(G330), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT91), .ZN(new_n775));
  INV_X1    g0575(.A(new_n656), .ZN(new_n776));
  INV_X1    g0576(.A(new_n710), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n773), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT94), .ZN(G396));
  NAND2_X1  g0580(.A1(new_n661), .A2(new_n420), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n431), .A2(new_n434), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n431), .B2(new_n781), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n690), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n651), .C1(new_n621), .C2(new_n630), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n704), .A2(G330), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT98), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n790), .B(new_n777), .C1(new_n788), .C2(new_n787), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n789), .A2(KEYINPUT98), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n784), .A2(new_n717), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n720), .A2(new_n717), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT95), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n710), .B1(G77), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n754), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n423), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G97), .A2(new_n767), .B1(new_n735), .B2(G303), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT96), .B(G283), .Z(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n731), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n271), .B1(new_n745), .B2(G311), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n803), .B1(new_n462), .B2(new_n741), .C1(new_n726), .C2(new_n737), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n751), .A2(new_n569), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n799), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n738), .A2(G143), .B1(new_n742), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n731), .B2(new_n317), .C1(new_n810), .C2(new_n758), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT34), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n271), .B1(new_n744), .B2(new_n813), .C1(new_n725), .C2(new_n202), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n752), .B2(G68), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n812), .B(new_n815), .C1(new_n759), .C2(new_n798), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n808), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n797), .B1(new_n818), .B2(new_n720), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G384));
  NOR3_X1   g0621(.A1(new_n215), .A2(new_n214), .A3(new_n462), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n583), .B(KEYINPUT99), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT35), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT36), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n670), .A2(new_n765), .A3(new_n381), .A4(new_n379), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n201), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n286), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT38), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n408), .B1(new_n403), .B2(new_n367), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n649), .B1(new_n391), .B2(new_n395), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n834), .A2(KEYINPUT37), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n378), .A2(new_n386), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n388), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n399), .B1(new_n838), .B2(new_n402), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT102), .B1(new_n839), .B2(new_n649), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n387), .A2(new_n252), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n395), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT102), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n650), .ZN(new_n845));
  INV_X1    g0645(.A(new_n367), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n840), .A2(new_n845), .A3(new_n408), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n836), .B1(KEYINPUT37), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n840), .A2(new_n845), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n412), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n833), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n408), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n396), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n391), .A2(new_n395), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n650), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n857), .A3(new_n858), .A4(new_n408), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n412), .A2(new_n850), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n296), .C2(new_n336), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n297), .A3(new_n299), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n307), .A2(new_n308), .A3(new_n266), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n267), .B(new_n661), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n267), .A2(new_n661), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n306), .A2(new_n309), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n431), .A2(new_n661), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT100), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT101), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n786), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n786), .B2(new_n872), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n863), .B(new_n870), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n634), .A2(new_n649), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(KEYINPUT103), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  AOI221_X4 g0680(.A(new_n833), .B1(new_n412), .B2(new_n850), .C1(new_n854), .C2(new_n859), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n859), .A2(KEYINPUT104), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n391), .A2(new_n395), .A3(new_n407), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n396), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(new_n858), .A4(new_n857), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n834), .B2(new_n835), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n412), .A2(new_n835), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n880), .B1(new_n881), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n865), .A2(new_n267), .A3(new_n651), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n852), .A2(new_n862), .A3(KEYINPUT39), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n879), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n870), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n786), .A2(new_n872), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT101), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n874), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n900), .A2(new_n863), .B1(new_n634), .B2(new_n649), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n689), .A2(new_n437), .A3(new_n692), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n689), .A2(new_n437), .A3(new_n906), .A4(new_n692), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n641), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n903), .B(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n881), .A2(new_n890), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n702), .A2(new_n703), .ZN(new_n911));
  NOR4_X1   g0711(.A1(new_n575), .A2(new_n501), .A3(new_n606), .A4(new_n661), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT106), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n784), .B1(new_n867), .B2(new_n869), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n693), .A2(new_n915), .A3(new_n702), .A4(new_n703), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT40), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n863), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n437), .A2(new_n913), .A3(new_n916), .ZN(new_n923));
  OAI21_X1  g0723(.A(G330), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n909), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n286), .B2(new_n707), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n909), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n832), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NOR2_X1   g0732(.A1(new_n713), .A2(new_n235), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n721), .B1(new_n209), .B2(new_n414), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n710), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(G107), .A2(new_n767), .B1(new_n735), .B2(G311), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n726), .B2(new_n731), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n271), .B1(new_n745), .B2(G317), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n440), .B2(new_n737), .C1(new_n741), .C2(new_n801), .ZN(new_n939));
  INV_X1    g0739(.A(new_n753), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT46), .B1(new_n940), .B2(G116), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n754), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n469), .C2(new_n751), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n725), .A2(new_n203), .B1(new_n737), .B2(new_n317), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT110), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n731), .A2(new_n384), .B1(new_n202), .B2(new_n753), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G143), .B2(new_n735), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n271), .B1(new_n744), .B2(new_n810), .C1(new_n201), .C2(new_n741), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(new_n218), .C2(new_n751), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n944), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n935), .B1(new_n953), .B2(new_n720), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n550), .A2(new_n573), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n661), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n618), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n629), .B2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n954), .B1(new_n772), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n601), .B(new_n605), .C1(new_n589), .C2(new_n651), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(new_n605), .C2(new_n651), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n665), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n666), .A2(new_n963), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n660), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n664), .A2(KEYINPUT109), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT109), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n659), .B2(new_n662), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n972), .B1(new_n974), .B2(new_n664), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n776), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n705), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n705), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n669), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n709), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n961), .A2(new_n962), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n605), .B1(new_n982), .B2(new_n540), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n963), .A2(new_n663), .A3(new_n662), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n651), .A2(new_n983), .B1(new_n984), .B2(KEYINPUT42), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(KEYINPUT42), .B2(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n986), .A2(KEYINPUT43), .A3(new_n958), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n660), .A2(new_n964), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n959), .B1(new_n981), .B2(new_n994), .ZN(G387));
  OR2_X1    g0795(.A1(new_n659), .A2(new_n772), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n232), .A2(new_n445), .A3(new_n271), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT50), .B1(new_n323), .B2(G50), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n445), .C1(new_n203), .C2(new_n249), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n323), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n370), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n672), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n668), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n721), .B1(new_n209), .B2(new_n423), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n710), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n753), .A2(new_n218), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n731), .A2(new_n323), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G159), .C2(new_n735), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n752), .A2(G97), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n551), .A2(new_n767), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n737), .A2(new_n759), .B1(new_n741), .B2(new_n203), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n370), .B(new_n1011), .C1(G150), .C2(new_n745), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n271), .B1(new_n745), .B2(G326), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n725), .A2(new_n801), .B1(new_n753), .B2(new_n726), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n738), .A2(G317), .B1(new_n742), .B2(G303), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n730), .A2(G311), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n735), .A2(G322), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT48), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1014), .B1(new_n462), .B2(new_n751), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1013), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1005), .B1(new_n1027), .B2(new_n720), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n976), .A2(new_n709), .B1(new_n996), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n977), .A2(new_n669), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n705), .A2(new_n976), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT112), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(G393));
  NOR2_X1   g0834(.A1(new_n971), .A2(new_n977), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n669), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n971), .A2(new_n977), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n971), .A2(new_n708), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n240), .A2(new_n713), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n721), .B1(new_n209), .B2(new_n469), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n710), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G150), .A2(new_n735), .B1(new_n738), .B2(G159), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT51), .ZN(new_n1045));
  INV_X1    g0845(.A(G143), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n271), .B1(new_n744), .B2(new_n1046), .C1(new_n323), .C2(new_n741), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n767), .A2(G77), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n203), .B2(new_n753), .C1(new_n731), .C2(new_n201), .ZN(new_n1049));
  NOR4_X1   g0849(.A1(new_n1045), .A2(new_n805), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G317), .A2(new_n735), .B1(new_n738), .B2(G311), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT52), .Z(new_n1054));
  OAI22_X1  g0854(.A1(new_n725), .A2(new_n462), .B1(new_n801), .B2(new_n753), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G303), .B2(new_n730), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n370), .B1(new_n741), .B2(new_n726), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G322), .B2(new_n745), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n763), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1052), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1043), .B1(new_n1061), .B2(new_n720), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n963), .B2(new_n772), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1039), .A2(new_n1040), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  INV_X1    g0865(.A(KEYINPUT115), .ZN(new_n1066));
  INV_X1    g0866(.A(G330), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n784), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n913), .A2(new_n916), .A3(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(new_n897), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n685), .A2(new_n651), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT90), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n685), .A2(new_n686), .A3(new_n651), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n784), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n871), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n783), .B1(new_n687), .B2(new_n688), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(KEYINPUT114), .A3(new_n871), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n870), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n910), .A2(new_n893), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1083), .A2(new_n892), .B1(new_n891), .B2(new_n894), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1070), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1068), .A2(new_n704), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n897), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1084), .B(new_n1088), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1066), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1088), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1082), .A2(new_n1085), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1084), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(KEYINPUT115), .C1(new_n1093), .C2(new_n1070), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n923), .A2(G330), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1087), .A2(new_n897), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1070), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n899), .A2(new_n874), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1069), .A2(new_n897), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1091), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n908), .B(new_n1095), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n905), .A2(new_n907), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n642), .A3(new_n1095), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1102), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT116), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1108), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1090), .A2(new_n1094), .A3(new_n1105), .A4(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1036), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n891), .A2(new_n894), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n717), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n710), .B1(new_n322), .B2(new_n796), .ZN(new_n1122));
  INV_X1    g0922(.A(G283), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1048), .B1(new_n731), .B2(new_n423), .C1(new_n1123), .C2(new_n758), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n370), .B1(new_n744), .B2(new_n726), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n737), .A2(new_n462), .B1(new_n741), .B2(new_n469), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n203), .B2(new_n751), .C1(new_n569), .C2(new_n798), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1130), .A2(new_n742), .B1(G137), .B2(new_n730), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT118), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n271), .B1(new_n737), .B2(new_n813), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n735), .A2(G128), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n384), .B2(new_n725), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(G125), .C2(new_n745), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n753), .A2(new_n317), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(new_n201), .C2(new_n751), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1128), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1122), .B1(new_n1140), .B2(new_n720), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1116), .A2(new_n709), .B1(new_n1121), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1119), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT119), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT119), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1119), .A2(new_n1145), .A3(new_n1142), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(G378));
  OAI21_X1  g0948(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n342), .A2(new_n344), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n650), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n633), .B(new_n1151), .C1(new_n638), .C2(new_n639), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n922), .B2(G330), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1067), .B(new_n1158), .C1(new_n918), .C2(new_n921), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1160), .A2(new_n1161), .B1(new_n902), .B2(new_n896), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n888), .A2(new_n889), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n862), .B1(new_n1163), .B2(KEYINPUT38), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n920), .B1(new_n1164), .B2(new_n919), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n913), .A2(new_n914), .A3(new_n920), .A4(new_n916), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n862), .B2(new_n852), .ZN(new_n1167));
  OAI21_X1  g0967(.A(G330), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1158), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n901), .B2(KEYINPUT103), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n877), .A2(new_n878), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT103), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n922), .A2(G330), .A3(new_n1159), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1169), .A2(new_n1171), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1162), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1070), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n1117), .A3(new_n1092), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1177), .B1(new_n1181), .B2(new_n1108), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT121), .B1(new_n1182), .B2(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1036), .B1(new_n1182), .B2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1162), .A2(new_n1176), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1086), .A2(new_n1104), .A3(new_n1089), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n1107), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT57), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1183), .A2(new_n1184), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n201), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n710), .B1(new_n1192), .B2(new_n796), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n271), .A2(G41), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n759), .B1(G33), .B2(G41), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1194), .B1(new_n1123), .B2(new_n744), .C1(new_n423), .C2(new_n737), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n551), .B2(new_n742), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n752), .A2(G58), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1006), .B1(G68), .B2(new_n767), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G97), .A2(new_n730), .B1(new_n735), .B2(G116), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G150), .A2(new_n767), .B1(new_n735), .B2(G125), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1130), .A2(new_n940), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n730), .A2(G132), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n738), .A2(G128), .B1(new_n742), .B2(G137), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n745), .C2(G124), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n384), .C2(new_n751), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1204), .B1(new_n1203), .B2(new_n1202), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1193), .B1(new_n1214), .B2(new_n720), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1159), .B2(new_n718), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT120), .Z(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1185), .B2(new_n709), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1191), .A2(new_n1218), .ZN(G375));
  NAND2_X1  g1019(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1114), .A2(new_n1105), .A3(new_n980), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n897), .A2(new_n717), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n710), .B1(G68), .B2(new_n796), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n370), .B1(new_n745), .B2(G128), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n810), .B2(new_n737), .C1(new_n317), .C2(new_n741), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n758), .A2(new_n813), .B1(new_n759), .B2(new_n725), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1130), .A2(new_n730), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n754), .A2(G159), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1227), .A2(new_n1199), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n754), .A2(G97), .B1(G303), .B2(new_n745), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n752), .A2(G77), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n370), .B1(new_n737), .B2(new_n1123), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G107), .B2(new_n742), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G116), .A2(new_n730), .B1(new_n735), .B2(G294), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1010), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1223), .B1(new_n1238), .B2(new_n720), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1112), .A2(new_n709), .B1(new_n1222), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1221), .A2(new_n1240), .ZN(G381));
  XNOR2_X1  g1041(.A(G375), .B(KEYINPUT124), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT123), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1143), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1119), .A2(KEYINPUT123), .A3(new_n1142), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(G390), .A2(G387), .A3(G384), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  AND4_X1   g1048(.A1(new_n1240), .A2(new_n1247), .A3(new_n1221), .A4(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1242), .A2(new_n1246), .A3(new_n1249), .ZN(G407));
  INV_X1    g1050(.A(G343), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1242), .A2(new_n1246), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G407), .A2(new_n1254), .A3(G213), .ZN(G409));
  NAND4_X1  g1055(.A1(new_n1191), .A2(new_n1144), .A3(new_n1146), .A4(new_n1218), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n980), .B(new_n1185), .C1(new_n1186), .C2(new_n1107), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1182), .A2(new_n1259), .A3(new_n980), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1260), .A3(new_n1218), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1244), .A2(new_n1261), .A3(new_n1245), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1256), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1252), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1265), .A2(new_n1220), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n669), .B1(new_n1265), .B2(new_n1220), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1240), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1268), .A2(new_n820), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n820), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G2897), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1252), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1269), .B(new_n1270), .C1(new_n1272), .C2(new_n1252), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1264), .B2(new_n1271), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1064), .A2(G387), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1064), .A2(G387), .ZN(new_n1282));
  AND2_X1   g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1281), .A2(new_n1282), .B1(new_n1248), .B2(new_n1283), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1064), .A2(G387), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1283), .A2(new_n1248), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1064), .A2(G387), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1253), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1271), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1278), .A2(new_n1280), .A3(new_n1290), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1291), .A2(new_n1295), .A3(new_n1292), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1291), .B2(new_n1276), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1296), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1294), .B1(new_n1300), .B2(new_n1290), .ZN(G405));
  NAND2_X1  g1101(.A1(new_n1246), .A2(G375), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1256), .B1(new_n1302), .B2(KEYINPUT127), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1289), .B(new_n1271), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1305), .B(new_n1306), .ZN(G402));
endmodule


