//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(G58), .A2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n208), .B1(new_n212), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n217), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n238), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT70), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT14), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1698), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G226), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n255), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n251), .B1(new_n261), .B2(KEYINPUT69), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(KEYINPUT69), .B2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT13), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G41), .A2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n265), .A2(G1), .A3(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(KEYINPUT64), .A2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT64), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n265), .ZN(new_n271));
  INV_X1    g0071(.A(new_n251), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n267), .B1(new_n273), .B2(G238), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n263), .A2(new_n264), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n264), .B1(new_n263), .B2(new_n274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G169), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n248), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI221_X1 g0080(.A(G169), .B1(new_n246), .B2(new_n247), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(G179), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n268), .A2(G13), .A3(G20), .A4(new_n269), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n240), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT12), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n209), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT64), .B(G1), .Z(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n287), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n217), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n210), .A2(G33), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n299), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n289), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(new_n301), .B(KEYINPUT11), .Z(new_n302));
  NOR2_X1   g0102(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n283), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n278), .B2(G190), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n278), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n296), .A2(G150), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n310), .B1(new_n201), .B2(new_n210), .C1(new_n311), .C2(new_n299), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(new_n289), .B1(new_n217), .B2(new_n285), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n293), .A2(G50), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n291), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT9), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n254), .B2(new_n255), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n320), .A2(G223), .B1(new_n323), .B2(G77), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n256), .A2(G222), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n272), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n267), .B1(new_n273), .B2(G226), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n318), .B1(new_n329), .B2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n316), .B(new_n330), .C1(new_n331), .C2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(new_n279), .ZN(new_n335));
  AND2_X1   g0135(.A1(KEYINPUT65), .A2(G179), .ZN(new_n336));
  NOR2_X1   g0136(.A1(KEYINPUT65), .A2(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n335), .B(new_n315), .C1(new_n339), .C2(new_n329), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n273), .A2(G244), .ZN(new_n342));
  INV_X1    g0142(.A(new_n267), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n320), .A2(G238), .B1(new_n323), .B2(G107), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n258), .A2(G232), .A3(new_n319), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n251), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n338), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n279), .B1(new_n344), .B2(new_n347), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n270), .A2(new_n210), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n291), .A2(new_n351), .A3(new_n202), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G20), .A2(G77), .ZN(new_n353));
  INV_X1    g0153(.A(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT15), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G87), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n353), .B1(new_n311), .B2(new_n297), .C1(new_n359), .C2(new_n299), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n352), .B1(new_n289), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n285), .A2(new_n202), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT67), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n349), .A2(new_n350), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n348), .A2(G190), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n363), .A3(new_n361), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n348), .A2(new_n307), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n334), .A2(new_n341), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n240), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n373), .B2(new_n213), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n296), .A2(G159), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n254), .A2(new_n210), .A3(new_n255), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n255), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(KEYINPUT71), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n383), .A2(KEYINPUT72), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT72), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n384), .A2(G68), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n377), .C1(new_n386), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n240), .B1(new_n380), .B2(new_n382), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n376), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT73), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(KEYINPUT73), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n391), .A2(new_n289), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n311), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n293), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n291), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n293), .A2(KEYINPUT74), .A3(new_n398), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n401), .A2(new_n402), .B1(new_n285), .B2(new_n311), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n218), .A2(G1698), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(G223), .B2(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n272), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n251), .B(G232), .C1(new_n270), .C2(new_n265), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n343), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n338), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G169), .B2(new_n411), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n404), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n404), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n409), .A2(new_n331), .A3(new_n343), .A4(new_n410), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n410), .A2(new_n343), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n251), .B1(new_n406), .B2(new_n407), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n307), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT75), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT75), .B1(new_n419), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n397), .A2(new_n403), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n425), .A4(new_n403), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n416), .A2(new_n418), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n309), .A2(new_n371), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n268), .A2(G45), .A3(new_n269), .ZN(new_n432));
  AND2_X1   g0232(.A1(KEYINPUT5), .A2(G41), .ZN(new_n433));
  NOR2_X1   g0233(.A1(KEYINPUT5), .A2(G41), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(G257), .B(new_n251), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n266), .B1(new_n249), .B2(new_n250), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT5), .B(G41), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n292), .A2(new_n437), .A3(G45), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(G244), .B(new_n319), .C1(new_n321), .C2(new_n322), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n442), .A2(KEYINPUT77), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n442), .B2(KEYINPUT77), .ZN(new_n445));
  OAI211_X1 g0245(.A(G250), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n441), .B1(new_n449), .B2(new_n251), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n284), .A2(G97), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n291), .B1(G33), .B2(new_n292), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n296), .A2(G77), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT76), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT6), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n456), .A2(new_n457), .A3(G107), .ZN(new_n458));
  XNOR2_X1  g0258(.A(G97), .B(G107), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n455), .B1(new_n210), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G107), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n380), .B2(new_n382), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n289), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n450), .A2(new_n279), .B1(new_n453), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT78), .B1(new_n449), .B2(new_n251), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  INV_X1    g0267(.A(new_n448), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n442), .A2(KEYINPUT77), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n443), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n272), .C1(new_n470), .C2(new_n444), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n440), .A2(KEYINPUT79), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n436), .A2(new_n439), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n466), .A2(new_n471), .A3(new_n338), .A4(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n466), .A2(new_n471), .A3(new_n475), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT80), .A4(new_n475), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(G200), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n464), .A2(new_n453), .ZN(new_n483));
  INV_X1    g0283(.A(new_n450), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G190), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n477), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n284), .A2(G107), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT25), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n452), .A2(G107), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n210), .B(G87), .C1(new_n321), .C2(new_n322), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n258), .A2(new_n494), .A3(new_n210), .A4(G87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G116), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(G20), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n499), .A2(new_n498), .A3(G20), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n496), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n496), .B2(new_n504), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n289), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n491), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(G264), .B(new_n251), .C1(new_n432), .C2(new_n435), .ZN(new_n510));
  OAI211_X1 g0310(.A(G250), .B(new_n319), .C1(new_n321), .C2(new_n322), .ZN(new_n511));
  INV_X1    g0311(.A(G294), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n253), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n320), .A2(new_n514), .A3(G257), .ZN(new_n515));
  OAI211_X1 g0315(.A(G257), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT84), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n510), .B(new_n439), .C1(new_n518), .C2(new_n251), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n279), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n509), .B(new_n520), .C1(G179), .C2(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(G200), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n320), .B2(G257), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n516), .A2(KEYINPUT84), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n272), .B1(new_n525), .B2(new_n513), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(G190), .A3(new_n439), .A4(new_n510), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n522), .A2(new_n527), .A3(new_n491), .A4(new_n508), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n521), .A2(KEYINPUT85), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n320), .A2(G264), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n258), .A2(G257), .A3(new_n319), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n323), .A2(G303), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n272), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n251), .B1(new_n432), .B2(new_n435), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n539), .A2(new_n220), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n540), .A3(new_n439), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n285), .A2(new_n219), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n268), .A2(G33), .A3(new_n269), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n284), .A2(new_n290), .A3(new_n545), .A4(G116), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n288), .A2(new_n209), .B1(G20), .B2(new_n219), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n447), .B(new_n210), .C1(G33), .C2(new_n457), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n547), .A2(KEYINPUT20), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n547), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n544), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n541), .B2(new_n331), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n543), .A2(new_n553), .A3(KEYINPUT82), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n537), .A2(new_n272), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n439), .B1(new_n539), .B2(new_n220), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n551), .B1(new_n558), .B2(G190), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n559), .B2(new_n542), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n292), .A2(new_n437), .A3(G45), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n432), .A2(G250), .A3(new_n251), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G244), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n565));
  OAI211_X1 g0365(.A(G238), .B(new_n319), .C1(new_n321), .C2(new_n322), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n499), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n272), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G200), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n284), .A2(new_n358), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n210), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n354), .A2(new_n457), .A3(new_n462), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n210), .B(G68), .C1(new_n321), .C2(new_n322), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n299), .B2(new_n457), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n571), .B1(new_n579), .B2(new_n289), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n284), .A2(new_n290), .A3(new_n545), .A4(G87), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n564), .A2(G190), .A3(new_n568), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n570), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n564), .A2(new_n338), .A3(new_n568), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n284), .A2(new_n290), .A3(new_n545), .A4(new_n358), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n562), .A2(new_n563), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n272), .B2(new_n567), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n585), .B(new_n587), .C1(new_n589), .C2(G169), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n584), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n541), .A2(G169), .A3(new_n551), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  INV_X1    g0397(.A(G179), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n556), .A2(new_n598), .A3(new_n557), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n596), .A2(new_n597), .B1(new_n599), .B2(new_n551), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n541), .A2(KEYINPUT21), .A3(G169), .A4(new_n551), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n561), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n431), .A2(new_n486), .A3(new_n533), .A4(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n341), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n416), .A2(new_n418), .ZN(new_n606));
  INV_X1    g0406(.A(new_n365), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n283), .B2(new_n304), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n428), .A2(new_n429), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n308), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT87), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n334), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n605), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n465), .A2(new_n476), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT86), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n579), .A2(new_n289), .ZN(new_n619));
  INV_X1    g0419(.A(new_n571), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n581), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n580), .B2(new_n581), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n583), .B1(new_n589), .B2(new_n307), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n590), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n617), .A2(new_n625), .A3(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n477), .A2(new_n594), .A3(new_n592), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(KEYINPUT26), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n482), .A2(new_n485), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n520), .B1(G179), .B2(new_n519), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n491), .A2(new_n508), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n600), .B(new_n601), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n570), .B(new_n583), .C1(new_n621), .C2(new_n622), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n528), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n629), .A2(new_n617), .A3(new_n632), .A4(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n628), .A2(new_n636), .A3(new_n590), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n431), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n616), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n292), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n552), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n561), .A2(new_n602), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n602), .B2(new_n649), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT88), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n509), .A2(new_n647), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT89), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n533), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n521), .A2(new_n648), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n596), .A2(new_n597), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n599), .A2(new_n551), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n661), .A2(new_n601), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n647), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n533), .A2(new_n655), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n521), .B2(new_n647), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n660), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n206), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n574), .A2(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n215), .B2(new_n670), .ZN(new_n673));
  XOR2_X1   g0473(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n674));
  XNOR2_X1  g0474(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n590), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n634), .B1(new_n663), .B2(new_n521), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n486), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT26), .B1(new_n617), .B2(new_n625), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(KEYINPUT29), .A3(new_n648), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n647), .B1(new_n678), .B2(new_n628), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(KEYINPUT29), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n533), .A2(new_n603), .A3(new_n486), .A4(new_n648), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n526), .A2(new_n510), .ZN(new_n686));
  NOR2_X1   g0486(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n569), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n484), .A2(new_n686), .A3(new_n599), .A4(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n688), .A2(new_n526), .A3(new_n510), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n484), .A3(new_n599), .A4(new_n692), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n558), .A2(new_n339), .A3(new_n589), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n478), .A3(new_n519), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n647), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n685), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n684), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n675), .B1(new_n707), .B2(G1), .ZN(G364));
  XNOR2_X1  g0508(.A(new_n641), .B(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G45), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G1), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n669), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n652), .B2(G330), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G330), .B2(new_n652), .ZN(new_n714));
  INV_X1    g0514(.A(new_n712), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n209), .B1(G20), .B2(new_n279), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n210), .A2(new_n331), .A3(new_n307), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n339), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G190), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n720), .A2(G326), .B1(G294), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  NOR2_X1   g0525(.A1(new_n210), .A2(new_n331), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n307), .A2(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n210), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n721), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(G303), .A2(new_n729), .B1(new_n732), .B2(G329), .ZN(new_n733));
  INV_X1    g0533(.A(G283), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n727), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n323), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n730), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n338), .A2(new_n737), .A3(new_n307), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT33), .B(G317), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n339), .A2(new_n307), .A3(new_n726), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n338), .A2(new_n737), .A3(G200), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n742), .A2(G322), .B1(G311), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n725), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n731), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT32), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n719), .A2(new_n217), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n728), .A2(new_n354), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n258), .B1(new_n735), .B2(new_n462), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n723), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n457), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n738), .A2(G68), .B1(new_n747), .B2(new_n748), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n742), .A2(G58), .B1(G77), .B2(new_n743), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n752), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n717), .B1(new_n745), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n668), .A2(new_n323), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G355), .B1(new_n219), .B2(new_n668), .ZN(new_n761));
  INV_X1    g0561(.A(G45), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n244), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n668), .A2(new_n258), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G45), .B2(new_n215), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n761), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT93), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n771), .B(new_n716), .C1(new_n766), .C2(new_n767), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n715), .B(new_n759), .C1(new_n768), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n771), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n652), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n714), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  NAND2_X1  g0577(.A1(new_n364), .A2(new_n647), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n607), .B1(new_n370), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n365), .A2(new_n647), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n637), .A2(new_n648), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(KEYINPUT97), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT97), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n683), .A2(new_n784), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n683), .B2(new_n781), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(new_n705), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT98), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n712), .B1(new_n787), .B2(new_n705), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n716), .A2(new_n769), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n712), .B1(G77), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT95), .Z(new_n797));
  AOI22_X1  g0597(.A1(G107), .A2(new_n729), .B1(new_n732), .B2(G311), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n798), .B(new_n323), .C1(new_n354), .C2(new_n735), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n754), .B(new_n799), .C1(G303), .C2(new_n720), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n742), .A2(G294), .B1(G116), .B2(new_n743), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n738), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n803), .A2(KEYINPUT96), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(KEYINPUT96), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n802), .B1(G283), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n720), .A2(G137), .B1(new_n738), .B2(G150), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n742), .A2(G143), .ZN(new_n810));
  INV_X1    g0610(.A(new_n743), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n810), .C1(new_n746), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n258), .B1(new_n728), .B2(new_n217), .ZN(new_n814));
  INV_X1    g0614(.A(new_n735), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G68), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n731), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n814), .B(new_n818), .C1(G58), .C2(new_n723), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n808), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n797), .B1(new_n820), .B2(new_n717), .C1(new_n781), .C2(new_n770), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n793), .A2(new_n821), .ZN(G384));
  NOR2_X1   g0622(.A1(new_n709), .A2(new_n292), .ZN(new_n823));
  INV_X1    g0623(.A(G330), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  INV_X1    g0626(.A(new_n403), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT72), .B1(new_n383), .B2(new_n385), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n388), .A2(new_n387), .A3(new_n389), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n376), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n290), .B1(new_n830), .B2(KEYINPUT16), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n377), .B1(new_n386), .B2(new_n390), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n392), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n827), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n426), .B(KEYINPUT99), .C1(new_n834), .C2(new_n413), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n391), .A2(new_n289), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n830), .A2(KEYINPUT16), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n403), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n645), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n838), .A2(new_n414), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT99), .B1(new_n842), .B2(new_n426), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n826), .B(KEYINPUT37), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n840), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n430), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n404), .A2(new_n839), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n415), .A2(new_n848), .A3(new_n849), .A4(new_n426), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT100), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n426), .B1(new_n834), .B2(new_n413), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n835), .A3(new_n840), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n855), .B2(KEYINPUT37), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n825), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n841), .B2(new_n843), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n850), .A2(KEYINPUT100), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n844), .A4(new_n846), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n702), .A2(KEYINPUT102), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n700), .A2(new_n864), .A3(new_n701), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n685), .A2(new_n863), .A3(new_n703), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n303), .A2(new_n648), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n305), .A2(new_n308), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n283), .A2(new_n867), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n866), .A2(new_n871), .A3(new_n781), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n848), .B1(new_n606), .B2(new_n609), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n415), .A2(new_n848), .A3(new_n426), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(new_n849), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n825), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n861), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n873), .A2(new_n881), .A3(KEYINPUT40), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n431), .A2(new_n866), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n824), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n606), .A2(new_n839), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n780), .B1(new_n783), .B2(new_n785), .ZN(new_n889));
  INV_X1    g0689(.A(new_n871), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n891), .B2(new_n862), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n305), .A2(new_n647), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n431), .B(new_n682), .C1(KEYINPUT29), .C2(new_n683), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n616), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n898), .B(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n823), .B1(new_n887), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n902), .B2(new_n887), .ZN(new_n904));
  INV_X1    g0704(.A(new_n460), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n219), .B(new_n212), .C1(new_n905), .C2(KEYINPUT35), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(KEYINPUT35), .B2(new_n905), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  OAI21_X1  g0708(.A(G77), .B1(new_n372), .B2(new_n240), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n239), .B1(new_n215), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n640), .A3(new_n270), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n908), .A3(new_n911), .ZN(G367));
  NOR2_X1   g0712(.A1(new_n771), .A2(new_n716), .ZN(new_n913));
  INV_X1    g0713(.A(new_n764), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n913), .B1(new_n206), .B2(new_n359), .C1(new_n234), .C2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n712), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n623), .A2(new_n647), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n590), .A3(new_n633), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n590), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n753), .A2(new_n240), .ZN(new_n920));
  AOI22_X1  g0720(.A1(G77), .A2(new_n815), .B1(new_n732), .B2(G137), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n258), .C1(new_n372), .C2(new_n728), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n920), .B(new_n922), .C1(G143), .C2(new_n720), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n742), .A2(G150), .B1(G50), .B2(new_n743), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n746), .C2(new_n806), .ZN(new_n925));
  INV_X1    g0725(.A(G311), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n728), .A2(new_n219), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n719), .A2(new_n926), .B1(new_n927), .B2(KEYINPUT46), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(KEYINPUT46), .B2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(G317), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n323), .B1(new_n731), .B2(new_n930), .C1(new_n457), .C2(new_n735), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n742), .B2(G303), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n929), .B(new_n932), .C1(new_n806), .C2(new_n512), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n743), .A2(G283), .B1(G107), .B2(new_n723), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT108), .Z(new_n935));
  OAI21_X1  g0735(.A(new_n925), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT47), .Z(new_n937));
  OAI221_X1 g0737(.A(new_n916), .B1(new_n774), .B2(new_n919), .C1(new_n937), .C2(new_n717), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT104), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n483), .A2(new_n647), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n486), .A2(new_n941), .B1(new_n477), .B2(new_n647), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n665), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n521), .B1(new_n482), .B2(new_n485), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n648), .B1(new_n945), .B2(new_n477), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT43), .B1(new_n919), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n919), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n660), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n942), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(new_n955), .C2(new_n953), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n711), .B(KEYINPUT107), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n660), .A2(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n666), .A2(new_n942), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT44), .Z(new_n964));
  NOR2_X1   g0764(.A1(new_n666), .A2(new_n942), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n653), .B(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n706), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n962), .A2(new_n967), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n707), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n669), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n961), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n938), .B1(new_n959), .B2(new_n977), .ZN(G387));
  NOR2_X1   g0778(.A1(new_n970), .A2(new_n960), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT109), .Z(new_n980));
  OAI22_X1  g0780(.A1(new_n803), .A2(new_n311), .B1(new_n359), .B2(new_n753), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G159), .B2(new_n720), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n258), .B1(new_n735), .B2(new_n457), .ZN(new_n983));
  INV_X1    g0783(.A(G150), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n728), .A2(new_n202), .B1(new_n731), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(G68), .C2(new_n743), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n982), .B(new_n986), .C1(new_n217), .C2(new_n741), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n729), .A2(G294), .B1(new_n723), .B2(G283), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n807), .A2(G311), .B1(G322), .B2(new_n720), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n743), .A2(G303), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n930), .B2(new_n741), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT111), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT48), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n988), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT112), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n996), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n258), .B1(new_n732), .B2(G326), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n219), .C2(new_n735), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT49), .B1(new_n998), .B2(new_n999), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n987), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n716), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n231), .A2(new_n762), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n398), .A2(new_n217), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n671), .B(new_n762), .C1(new_n240), .C2(new_n202), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n764), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1006), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n760), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(G107), .B2(new_n206), .C1(new_n671), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n715), .B1(new_n1015), .B2(new_n913), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1005), .B(new_n1016), .C1(new_n658), .C2(new_n774), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n980), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n971), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n970), .A2(new_n706), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n669), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1021), .ZN(G393));
  XNOR2_X1  g0822(.A(new_n967), .B(new_n954), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n973), .B(new_n669), .C1(new_n971), .C2(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n238), .A2(new_n764), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n913), .B1(new_n457), .B2(new_n206), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n741), .A2(new_n926), .B1(new_n719), .B2(new_n930), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT52), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n728), .A2(new_n734), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n323), .B1(new_n735), .B2(new_n462), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G322), .C2(new_n732), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n219), .B2(new_n753), .C1(new_n512), .C2(new_n811), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n807), .B2(G303), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n728), .A2(new_n240), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n258), .B1(new_n735), .B2(new_n354), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G143), .C2(new_n732), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n202), .B2(new_n753), .C1(new_n311), .C2(new_n811), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n807), .B2(G50), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n741), .A2(new_n746), .B1(new_n719), .B2(new_n984), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1028), .A2(new_n1033), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n712), .B1(new_n1025), .B2(new_n1026), .C1(new_n1041), .C2(new_n717), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n942), .B2(new_n771), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1023), .B2(new_n961), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1024), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(KEYINPUT113), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1024), .A2(KEYINPUT113), .A3(new_n1044), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G390));
  INV_X1    g0849(.A(KEYINPUT116), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n895), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n889), .B2(new_n890), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT39), .B1(new_n861), .B2(new_n880), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n780), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n681), .A2(new_n648), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n779), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT114), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT114), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n1056), .C1(new_n1057), .C2(new_n779), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n871), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n895), .B1(new_n861), .B2(new_n880), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1055), .A2(KEYINPUT115), .A3(new_n1064), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n779), .A2(new_n824), .A3(new_n780), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n866), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n871), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT115), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1050), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1055), .A2(new_n1064), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(KEYINPUT116), .A3(new_n1065), .A4(new_n1069), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n704), .A2(new_n1066), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n890), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1072), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n885), .A2(new_n824), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT117), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n901), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n889), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n871), .B1(new_n704), .B2(new_n1066), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n1069), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1078), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n871), .C2(new_n1067), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1083), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1080), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1072), .A2(new_n1076), .A3(new_n1079), .A4(new_n1091), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n669), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1072), .A2(new_n1076), .A3(new_n961), .A4(new_n1079), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n712), .B1(new_n398), .B2(new_n795), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n753), .A2(new_n746), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n729), .A2(G150), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G128), .C2(new_n720), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n742), .A2(G132), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n258), .B1(new_n731), .B2(new_n1103), .C1(new_n217), .C2(new_n735), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n743), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n807), .A2(G137), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1101), .A2(new_n1102), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n806), .A2(new_n462), .B1(new_n457), .B2(new_n811), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n719), .A2(new_n734), .B1(new_n753), .B2(new_n202), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n750), .A2(new_n258), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n816), .C1(new_n512), .C2(new_n731), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G116), .C2(new_n742), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1109), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1097), .B1(new_n1118), .B2(new_n716), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n894), .A2(new_n896), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1121), .B2(new_n770), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1096), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1095), .A2(new_n1124), .ZN(G378));
  NAND2_X1  g0925(.A1(new_n334), .A2(new_n340), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n315), .A2(new_n839), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n769), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n803), .A2(new_n457), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n920), .B(new_n1134), .C1(G116), .C2(new_n720), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n735), .A2(new_n372), .B1(new_n731), .B2(new_n734), .ZN(new_n1136));
  INV_X1    g0936(.A(G41), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n323), .C1(new_n728), .C2(new_n202), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(new_n742), .C2(G107), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1135), .B(new_n1139), .C1(new_n359), .C2(new_n811), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT58), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n720), .A2(G125), .B1(G150), .B2(new_n723), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n743), .A2(G137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n742), .A2(G128), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n729), .A2(KEYINPUT119), .A3(new_n1106), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT119), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n728), .B2(new_n1105), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(new_n803), .C2(new_n817), .ZN(new_n1150));
  OR3_X1    g0950(.A1(new_n1146), .A2(KEYINPUT59), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT59), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n815), .A2(G159), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G33), .B(G41), .C1(new_n732), .C2(G124), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n217), .B1(new_n321), .B2(G41), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1142), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n716), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n794), .A2(new_n217), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1133), .A2(new_n712), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n872), .B1(new_n861), .B2(new_n857), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n875), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n882), .B(G330), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1132), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1132), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n876), .A2(new_n1167), .A3(G330), .A4(new_n882), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1166), .A2(new_n898), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n898), .B1(new_n1168), .B2(new_n1166), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1162), .B1(new_n1173), .B2(new_n961), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1083), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1094), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n669), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1173), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1174), .B1(new_n1180), .B2(new_n1181), .ZN(G375));
  INV_X1    g0982(.A(new_n1090), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1175), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n976), .A3(new_n1092), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT120), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n960), .B(KEYINPUT121), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n715), .B1(new_n240), .B2(new_n794), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n811), .A2(new_n984), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n720), .A2(G132), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G137), .C2(new_n742), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G159), .A2(new_n729), .B1(new_n732), .B2(G128), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n323), .B1(new_n815), .B2(G58), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n217), .C2(new_n753), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n807), .B2(new_n1106), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n807), .A2(G116), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G97), .A2(new_n729), .B1(new_n732), .B2(G303), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n323), .C1(new_n202), .C2(new_n735), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n811), .A2(new_n462), .B1(new_n734), .B2(new_n741), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n719), .A2(new_n512), .B1(new_n753), .B2(new_n359), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1194), .A2(new_n1198), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1190), .B1(new_n717), .B2(new_n1205), .C1(new_n871), .C2(new_n770), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1189), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1187), .A2(new_n1208), .ZN(G381));
  OR2_X1    g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  INV_X1    g1010(.A(G384), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1048), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OR4_X1    g1013(.A1(G387), .A2(new_n1210), .A3(G381), .A4(new_n1213), .ZN(G407));
  OAI211_X1 g1014(.A(G407), .B(G213), .C1(G343), .C2(new_n1210), .ZN(G409));
  NAND2_X1  g1015(.A1(new_n1048), .A2(G387), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n959), .A2(new_n977), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n938), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT124), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1048), .B2(G387), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n776), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1212), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1219), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1216), .A2(new_n1218), .A3(new_n1220), .A4(new_n1223), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n646), .A2(G213), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G378), .B(new_n1174), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n670), .B1(new_n1080), .B2(new_n1092), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1123), .B1(new_n1231), .B2(new_n1094), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1162), .B1(new_n1173), .B2(new_n1188), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n976), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1094), .B2(new_n1175), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT123), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g1037(.A(KEYINPUT123), .B(new_n1234), .C1(new_n1175), .C2(new_n1094), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1232), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1229), .B1(new_n1230), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1184), .B1(KEYINPUT60), .B2(new_n1092), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1083), .A2(new_n1090), .A3(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n669), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1208), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1211), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G384), .B(new_n1208), .C1(new_n1241), .C2(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT62), .B1(new_n1240), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1230), .A2(new_n1239), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1228), .ZN(new_n1252));
  AOI211_X1 g1052(.A(KEYINPUT125), .B(new_n1229), .C1(new_n1230), .C2(new_n1239), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1248), .A2(KEYINPUT62), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1249), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1229), .A2(G2897), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1247), .B(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1227), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1254), .A2(KEYINPUT63), .A3(new_n1248), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT63), .B1(new_n1258), .B2(new_n1240), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1240), .A2(new_n1248), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1227), .A2(KEYINPUT61), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1264), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1263), .A2(new_n1269), .ZN(G405));
  NAND3_X1  g1070(.A1(G375), .A2(new_n1248), .A3(new_n1232), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G375), .A2(new_n1232), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1247), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1227), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1271), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1226), .A3(new_n1225), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1230), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1274), .A2(new_n1279), .A3(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


