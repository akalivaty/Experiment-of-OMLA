//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT65), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n211), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G223), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G222), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n202), .B2(new_n249), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n258), .A2(new_n262), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G226), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G169), .ZN(new_n268));
  INV_X1    g0068(.A(G179), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n267), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G150), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n214), .A2(G33), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n272), .B1(new_n206), .B2(new_n201), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n255), .B1(new_n207), .B2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(G50), .B1(new_n206), .B2(G1), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n282), .A2(new_n283), .B1(G50), .B2(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n284), .A2(new_n285), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n270), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n267), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n267), .A2(G200), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT9), .B(new_n278), .C1(new_n287), .C2(new_n288), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n294), .A2(new_n300), .A3(new_n296), .A4(new_n297), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n290), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n249), .A2(G232), .A3(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  INV_X1    g0104(.A(G226), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n304), .C1(new_n253), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n258), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n264), .B1(new_n265), .B2(G238), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(G169), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(G169), .C1(new_n310), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n307), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(G179), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n280), .A2(G20), .A3(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(new_n322), .B(KEYINPUT12), .Z(new_n323));
  INV_X1    g0123(.A(new_n282), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n321), .B1(new_n205), .B2(G20), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n321), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n273), .B2(new_n202), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n277), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n277), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n310), .B2(new_n311), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n317), .A2(new_n337), .A3(new_n318), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n333), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n273), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n271), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n202), .A2(new_n214), .B1(new_n274), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n277), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n202), .B1(new_n205), .B2(G20), .ZN(new_n348));
  INV_X1    g0148(.A(new_n281), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n202), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT72), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n281), .B2(G77), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n324), .A2(new_n348), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT70), .B(G107), .ZN(new_n356));
  INV_X1    g0156(.A(G232), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n355), .B1(new_n249), .B2(new_n356), .C1(new_n253), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n258), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n264), .B1(new_n265), .B2(G244), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n337), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n335), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n354), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n269), .B2(new_n362), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n354), .B2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n302), .A2(new_n334), .A3(new_n340), .A4(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n274), .B1(new_n205), .B2(G20), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n324), .A2(new_n369), .B1(new_n349), .B2(new_n274), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n321), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n271), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT64), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n378), .B1(new_n382), .B2(new_n249), .ZN(new_n383));
  AND2_X1   g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n377), .B1(new_n388), .B2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n276), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n214), .A3(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n247), .A2(new_n206), .A3(new_n248), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n378), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n321), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(new_n377), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n371), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n257), .A2(G232), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n263), .ZN(new_n400));
  OAI211_X1 g0200(.A(G223), .B(new_n252), .C1(new_n384), .C2(new_n385), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n258), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n269), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G169), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n407), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n386), .B2(new_n214), .ZN(new_n410));
  NOR4_X1   g0210(.A1(new_n384), .A2(new_n385), .A3(new_n378), .A4(G20), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n377), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n396), .A2(new_n414), .A3(new_n277), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n370), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n409), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n404), .A2(new_n258), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n399), .A2(new_n263), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n337), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G200), .B2(new_n405), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n423), .A3(new_n370), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n415), .A2(new_n423), .A3(KEYINPUT17), .A4(new_n370), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT74), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT74), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n419), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n368), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n205), .B(G45), .C1(new_n260), .C2(KEYINPUT5), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT78), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n257), .A2(G274), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n436), .ZN(new_n439));
  OAI211_X1 g0239(.A(G257), .B(new_n257), .C1(new_n439), .C2(new_n434), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT79), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n249), .A2(G244), .A3(new_n252), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(KEYINPUT4), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n445), .A2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n258), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n434), .B(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n437), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(new_n440), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n442), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G200), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n349), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n205), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n276), .A2(new_n281), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n392), .A2(new_n394), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n271), .A2(G77), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT75), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n459), .A2(new_n465), .A3(KEYINPUT6), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(KEYINPUT6), .B2(new_n459), .ZN(new_n474));
  XOR2_X1   g0274(.A(KEYINPUT76), .B(G107), .Z(new_n475));
  XNOR2_X1  g0275(.A(new_n474), .B(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n470), .B(new_n472), .C1(new_n476), .C2(new_n214), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n463), .B1(new_n477), .B2(new_n277), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n442), .A2(G190), .A3(new_n450), .A4(new_n456), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n458), .B(new_n478), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n341), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n281), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT19), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n214), .B1(new_n486), .B2(new_n304), .ZN(new_n487));
  INV_X1    g0287(.A(G87), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n356), .A2(new_n488), .A3(new_n459), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n249), .A2(new_n214), .A3(G68), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n486), .B1(new_n273), .B2(new_n459), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT81), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n485), .B1(new_n496), .B2(new_n277), .ZN(new_n497));
  INV_X1    g0297(.A(new_n462), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(G250), .B1(new_n261), .B2(G1), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(new_n257), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n249), .A2(G244), .A3(G1698), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(G238), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n507), .C1(new_n253), .C2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n509), .B2(new_n258), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G200), .ZN(new_n511));
  AOI211_X1 g0311(.A(G190), .B(new_n505), .C1(new_n509), .C2(new_n258), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n497), .B1(new_n341), .B2(new_n462), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(G179), .ZN(new_n516));
  INV_X1    g0316(.A(G169), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n501), .A2(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n349), .A2(new_n465), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT25), .ZN(new_n521));
  OR3_X1    g0321(.A1(new_n520), .A2(KEYINPUT83), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT83), .B1(new_n520), .B2(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n498), .A2(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  XOR2_X1   g0328(.A(KEYINPUT84), .B(G294), .Z(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G33), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n249), .A2(G257), .A3(G1698), .ZN(new_n531));
  INV_X1    g0331(.A(G250), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(new_n253), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n258), .ZN(new_n534));
  OAI211_X1 g0334(.A(G264), .B(new_n257), .C1(new_n439), .C2(new_n434), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n454), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n335), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G190), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT23), .B1(new_n469), .B2(new_n206), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n507), .A2(G20), .ZN(new_n540));
  NOR2_X1   g0340(.A1(KEYINPUT23), .A2(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n382), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n543), .A2(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n249), .A2(new_n214), .A3(G87), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n277), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n549), .B1(new_n544), .B2(new_n545), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(KEYINPUT24), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n528), .B(new_n538), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n457), .A2(G169), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n442), .A2(G179), .A3(new_n450), .A4(new_n456), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n478), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n483), .A2(new_n519), .A3(new_n556), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n249), .A2(G264), .A3(G1698), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n249), .A2(G257), .A3(new_n252), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n249), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n565), .A2(new_n258), .ZN(new_n566));
  OAI211_X1 g0366(.A(G270), .B(new_n257), .C1(new_n439), .C2(new_n434), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n454), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(KEYINPUT21), .B(G169), .C1(new_n566), .C2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n454), .A2(new_n567), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n565), .A2(new_n258), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n269), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n498), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n349), .A2(G116), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n206), .A2(G116), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n276), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n214), .B(new_n443), .C1(G33), .C2(new_n459), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n575), .A2(new_n576), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n572), .A2(new_n582), .A3(G169), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n573), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n582), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n572), .A2(G190), .ZN(new_n587));
  AOI21_X1  g0387(.A(G200), .B1(new_n570), .B2(new_n571), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n551), .A2(new_n552), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n276), .B1(new_n554), .B2(KEYINPUT24), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n527), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n536), .A2(new_n269), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(G169), .B2(new_n536), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n585), .B(new_n589), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n433), .A2(new_n561), .A3(new_n595), .ZN(G372));
  NAND2_X1  g0396(.A1(new_n408), .A2(new_n418), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n366), .A2(new_n354), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n334), .B1(new_n339), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n426), .A2(new_n427), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT74), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n428), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n597), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n604), .A2(KEYINPUT86), .B1(new_n299), .B2(new_n301), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n290), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n585), .B1(new_n592), .B2(new_n594), .ZN(new_n608));
  INV_X1    g0408(.A(new_n518), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n462), .A2(new_n341), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n485), .B(new_n610), .C1(new_n496), .C2(new_n277), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n609), .A2(new_n611), .B1(new_n500), .B2(new_n513), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n559), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n613), .A3(new_n556), .A4(new_n483), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n559), .A2(KEYINPUT85), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n617), .B(new_n478), .C1(new_n557), .C2(new_n558), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n615), .B(new_n519), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n515), .A2(new_n518), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n559), .B(new_n620), .C1(new_n500), .C2(new_n513), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(KEYINPUT26), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n432), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n607), .A2(new_n625), .ZN(G369));
  INV_X1    g0426(.A(new_n585), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n214), .A2(new_n280), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT27), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n214), .A2(new_n632), .A3(new_n280), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(G213), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n633), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n628), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n635), .A2(KEYINPUT88), .A3(G343), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n582), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n627), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n585), .A2(new_n589), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n592), .A2(new_n594), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n642), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n556), .B1(new_n651), .B2(new_n592), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n650), .A2(new_n642), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n585), .A2(new_n642), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n209), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G41), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n213), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n205), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n489), .A2(G116), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n624), .A2(new_n651), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n519), .A2(new_n615), .A3(new_n559), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n620), .B(KEYINPUT90), .Z(new_n673));
  NAND3_X1  g0473(.A1(new_n614), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n616), .A2(new_n618), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n615), .B1(new_n675), .B2(new_n519), .ZN(new_n676));
  OAI211_X1 g0476(.A(KEYINPUT29), .B(new_n651), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n442), .A2(new_n450), .A3(new_n456), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n566), .A2(new_n568), .A3(new_n269), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n510), .A2(new_n535), .A3(new_n534), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT89), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n510), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(G179), .B1(new_n570), .B2(new_n571), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n687), .A2(new_n536), .A3(new_n457), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n681), .A4(new_n682), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n642), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n642), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n561), .A2(new_n595), .A3(new_n642), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n679), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n678), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n668), .B1(new_n703), .B2(G1), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT91), .Z(G364));
  NOR2_X1   g0505(.A1(new_n382), .A2(new_n279), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G45), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n664), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n215), .B1(G20), .B2(new_n517), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n661), .A2(new_n386), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G355), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G116), .B2(new_n209), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n240), .A2(G45), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G45), .B2(new_n213), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n661), .A2(new_n249), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n214), .A2(G190), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT93), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n335), .A2(G179), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(KEYINPUT93), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G107), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(G20), .A3(G190), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n249), .C1(new_n488), .C2(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  NAND3_X1  g0533(.A1(new_n724), .A2(G179), .A3(G200), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n724), .A2(G179), .A3(new_n335), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n321), .A2(new_n734), .B1(new_n735), .B2(new_n202), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n214), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G97), .ZN(new_n740));
  NOR4_X1   g0540(.A1(new_n214), .A2(new_n269), .A3(new_n337), .A4(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G50), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n214), .A2(new_n269), .A3(new_n337), .A4(new_n335), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n740), .B1(new_n742), .B2(new_n372), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n725), .A2(new_n727), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT32), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT94), .B(G159), .Z(new_n750));
  OR3_X1    g0550(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n736), .B(new_n746), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n748), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G283), .A2(new_n729), .B1(new_n754), .B2(G329), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT96), .Z(new_n756));
  NAND2_X1  g0556(.A1(new_n741), .A2(G322), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n739), .A2(new_n529), .ZN(new_n758));
  INV_X1    g0558(.A(new_n731), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n249), .B1(new_n759), .B2(G303), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n735), .B1(new_n734), .B2(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n761), .B(new_n764), .C1(G326), .C2(new_n744), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n733), .A2(new_n753), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n714), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n710), .B1(new_n716), .B2(new_n723), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  INV_X1    g0569(.A(new_n713), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n646), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n648), .A2(new_n710), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n646), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  AOI22_X1  g0575(.A1(new_n640), .A2(new_n641), .B1(new_n347), .B2(new_n353), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n598), .B1(new_n364), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n651), .A2(new_n354), .A3(new_n366), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n669), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n779), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n624), .A2(new_n651), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n701), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n700), .A2(new_n780), .A3(new_n782), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(new_n709), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n714), .A2(new_n711), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n709), .B1(new_n202), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n729), .A2(G87), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n762), .B2(new_n748), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n741), .A2(G294), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n744), .A2(G303), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n249), .B1(new_n759), .B2(G107), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n791), .A2(new_n792), .A3(new_n740), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n574), .A2(new_n735), .B1(new_n734), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n790), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n729), .A2(G68), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n249), .B1(new_n731), .B2(new_n743), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G58), .B2(new_n739), .ZN(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n798), .B(new_n800), .C1(new_n801), .C2(new_n748), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT34), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G137), .A2(new_n744), .B1(new_n741), .B2(G143), .ZN(new_n804));
  INV_X1    g0604(.A(G150), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n805), .B2(new_n734), .C1(new_n750), .C2(new_n735), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n803), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n797), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n788), .B1(new_n809), .B2(new_n767), .C1(new_n781), .C2(new_n712), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n786), .A2(new_n810), .ZN(G384));
  XNOR2_X1  g0611(.A(new_n476), .B(KEYINPUT98), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT35), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT35), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n813), .A2(G116), .A3(new_n216), .A4(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n816));
  XNOR2_X1  g0616(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n213), .B(G77), .C1(new_n372), .C2(new_n321), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n743), .A2(G68), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n205), .B(G13), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n333), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n640), .B2(new_n641), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n339), .B(new_n823), .C1(new_n320), .C2(new_n333), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n642), .B(new_n333), .C1(new_n320), .C2(new_n339), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n781), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n697), .B2(new_n699), .ZN(new_n828));
  INV_X1    g0628(.A(new_n391), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n414), .B(new_n277), .C1(new_n389), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n370), .ZN(new_n831));
  INV_X1    g0631(.A(new_n638), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n424), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n407), .B1(new_n370), .B2(new_n830), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n409), .A2(new_n416), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n416), .A2(new_n832), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n424), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n597), .B1(new_n602), .B2(new_n428), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n833), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(KEYINPUT38), .B(new_n841), .C1(new_n842), .C2(new_n833), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT40), .B1(new_n828), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n823), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n334), .A2(new_n340), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n779), .B1(new_n851), .B2(new_n825), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n852), .B(KEYINPUT40), .C1(new_n696), .C2(new_n698), .ZN(new_n853));
  INV_X1    g0653(.A(new_n833), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n431), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n855), .A2(KEYINPUT101), .A3(KEYINPUT38), .A4(new_n841), .ZN(new_n856));
  XOR2_X1   g0656(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n416), .B(new_n832), .C1(new_n597), .C2(new_n600), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n837), .A2(new_n838), .A3(new_n424), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n840), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n846), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n853), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n849), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT104), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n697), .A2(new_n699), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n432), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(G330), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n334), .A2(new_n642), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n846), .A2(new_n863), .ZN(new_n876));
  INV_X1    g0676(.A(new_n862), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n856), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n845), .A2(KEYINPUT39), .A3(new_n846), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(KEYINPUT102), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT102), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT39), .B1(new_n864), .B2(new_n856), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n845), .A2(KEYINPUT39), .A3(new_n846), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n875), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n824), .A2(new_n826), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n782), .B2(new_n778), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n847), .B1(new_n597), .B2(new_n638), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT103), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n678), .B2(new_n433), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n671), .A2(new_n432), .A3(KEYINPUT103), .A4(new_n677), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n894), .A2(new_n607), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n892), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n873), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n205), .B2(new_n706), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n873), .A2(new_n897), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n821), .B1(new_n899), .B2(new_n900), .ZN(G367));
  OAI22_X1  g0701(.A1(new_n743), .A2(new_n735), .B1(new_n734), .B2(new_n750), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n739), .A2(G68), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n386), .B1(new_n759), .B2(G58), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n903), .B(new_n904), .C1(new_n742), .C2(new_n805), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n902), .B(new_n905), .C1(G143), .C2(new_n744), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n729), .A2(G77), .ZN(new_n907));
  INV_X1    g0707(.A(G137), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n748), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT109), .ZN(new_n910));
  AOI22_X1  g0710(.A1(G97), .A2(new_n729), .B1(new_n754), .B2(G317), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n759), .A2(G116), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT46), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n912), .A2(new_n913), .B1(new_n356), .B2(new_n738), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n249), .B(new_n914), .C1(new_n913), .C2(new_n912), .ZN(new_n915));
  AOI22_X1  g0715(.A1(G303), .A2(new_n741), .B1(new_n744), .B2(G311), .ZN(new_n916));
  INV_X1    g0716(.A(new_n735), .ZN(new_n917));
  INV_X1    g0717(.A(new_n734), .ZN(new_n918));
  AOI22_X1  g0718(.A1(G283), .A2(new_n917), .B1(new_n918), .B2(new_n529), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n911), .A2(new_n915), .A3(new_n916), .A4(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n910), .A2(KEYINPUT47), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT47), .B1(new_n910), .B2(new_n920), .ZN(new_n922));
  OR3_X1    g0722(.A1(new_n921), .A2(new_n922), .A3(new_n767), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n235), .A2(new_n722), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n716), .B1(new_n661), .B2(new_n484), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n709), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n651), .A2(new_n501), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n519), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n620), .B2(new_n927), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n923), .B(new_n926), .C1(new_n770), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n708), .A2(G1), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n656), .A2(new_n658), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(KEYINPUT106), .B1(new_n648), .B2(KEYINPUT107), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT106), .B1(new_n656), .B2(new_n658), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n656), .B2(new_n658), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n648), .A2(KEYINPUT107), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n483), .B(new_n560), .C1(new_n651), .C2(new_n478), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n559), .A2(new_n642), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n659), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT45), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT44), .B1(new_n659), .B2(new_n944), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n659), .A2(KEYINPUT44), .A3(new_n944), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n657), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n941), .A2(new_n703), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n947), .A2(new_n657), .A3(new_n948), .A4(new_n949), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT108), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n702), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n662), .B(KEYINPUT41), .Z(new_n957));
  OAI21_X1  g0757(.A(new_n933), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n560), .B1(new_n942), .B2(new_n650), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT105), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n642), .B1(new_n960), .B2(KEYINPUT105), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n656), .A2(new_n658), .A3(new_n944), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n961), .A2(new_n962), .B1(KEYINPUT42), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n929), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n968), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n951), .A2(new_n944), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n931), .B1(new_n958), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(G387));
  INV_X1    g0776(.A(new_n662), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n941), .B2(new_n703), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n703), .B2(new_n941), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n386), .B1(new_n728), .B2(new_n574), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G317), .A2(new_n741), .B1(new_n744), .B2(G322), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n564), .B2(new_n735), .C1(new_n762), .C2(new_n734), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT110), .Z(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT48), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT48), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n739), .A2(G283), .B1(new_n529), .B2(new_n759), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n980), .B(new_n989), .C1(G326), .C2(new_n754), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n738), .A2(new_n341), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n386), .B(new_n991), .C1(G77), .C2(new_n759), .ZN(new_n992));
  INV_X1    g0792(.A(G159), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n743), .B2(new_n742), .C1(new_n993), .C2(new_n745), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n321), .A2(new_n735), .B1(new_n734), .B2(new_n274), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n459), .A2(new_n728), .B1(new_n748), .B2(new_n805), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n714), .B1(new_n990), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n656), .A2(new_n770), .ZN(new_n999));
  INV_X1    g0799(.A(new_n722), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n231), .B2(G45), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n666), .B2(new_n717), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n274), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n743), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n261), .B1(new_n321), .B2(new_n202), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1005), .A2(new_n666), .A3(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1002), .A2(new_n1007), .B1(G107), .B2(new_n209), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n709), .B(new_n999), .C1(new_n715), .C2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n941), .A2(new_n932), .B1(new_n998), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n979), .A2(new_n1010), .ZN(G393));
  INV_X1    g0811(.A(KEYINPUT112), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n952), .B(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n955), .A3(new_n932), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n715), .B1(new_n459), .B2(new_n209), .C1(new_n1000), .C2(new_n243), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n710), .A2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n754), .A2(G143), .B1(G68), .B2(new_n759), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT114), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n249), .B1(new_n202), .B2(new_n738), .C1(new_n735), .C2(new_n274), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G50), .B2(new_n918), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n805), .A2(new_n745), .B1(new_n742), .B2(new_n993), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT51), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1023), .A3(new_n789), .A4(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n386), .B1(new_n795), .B2(new_n731), .C1(new_n738), .C2(new_n574), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G294), .B2(new_n917), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n564), .B2(new_n734), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G311), .A2(new_n741), .B1(new_n744), .B2(G317), .ZN(new_n1029));
  XOR2_X1   g0829(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n754), .A2(G322), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n730), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1018), .A2(new_n1025), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1016), .B1(new_n1034), .B2(new_n714), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT116), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n944), .A2(new_n770), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT113), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT113), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n953), .A2(new_n955), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n662), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1013), .A2(new_n955), .B1(new_n703), .B2(new_n941), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1014), .B(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(G390));
  NAND2_X1  g0844(.A1(new_n782), .A2(new_n778), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n888), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n875), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n882), .A2(new_n886), .A3(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n651), .B(new_n777), .C1(new_n674), .C2(new_n676), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n778), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n1046), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n878), .A3(new_n875), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n852), .B(G330), .C1(new_n696), .C2(new_n698), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1055), .B(KEYINPUT117), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1049), .A2(new_n1053), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(G330), .B(new_n781), .C1(new_n696), .C2(new_n698), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1051), .B1(new_n888), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n888), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n1055), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1062), .A2(new_n1058), .B1(new_n1064), .B2(new_n1045), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n432), .A2(G330), .A3(new_n869), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n894), .A2(new_n607), .A3(new_n895), .A4(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n977), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1057), .A2(new_n1059), .A3(new_n1068), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n882), .A2(new_n886), .A3(new_n711), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n787), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n710), .B1(new_n1003), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n754), .A2(G294), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n744), .A2(G283), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n386), .B1(new_n731), .B2(new_n488), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n738), .A2(new_n202), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G116), .C2(new_n741), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n798), .A2(new_n1076), .A3(new_n1077), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n459), .A2(new_n735), .B1(new_n734), .B2(new_n356), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT118), .Z(new_n1083));
  OAI21_X1  g0883(.A(new_n249), .B1(new_n738), .B2(new_n993), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G132), .B2(new_n741), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT54), .B(G143), .Z(new_n1086));
  NAND2_X1  g0886(.A1(new_n917), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n918), .A2(G137), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n759), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n731), .B2(new_n805), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1089), .A2(new_n1091), .B1(new_n744), .B2(G128), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(G125), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n743), .A2(new_n728), .B1(new_n748), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1081), .A2(new_n1083), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1075), .B1(new_n1096), .B2(new_n714), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1073), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1060), .B2(new_n933), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1072), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G378));
  INV_X1    g0901(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n289), .A2(new_n832), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n302), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n302), .A2(new_n1103), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1106));
  OR3_X1    g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n849), .A2(new_n866), .A3(G330), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT102), .B1(new_n880), .B2(new_n881), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n884), .A2(new_n885), .A3(new_n883), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n874), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1115), .B2(new_n890), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n848), .A2(new_n865), .A3(new_n679), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n887), .A2(new_n891), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n890), .A3(new_n1112), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1117), .B1(new_n887), .B2(new_n891), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1111), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1067), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1119), .A2(new_n1123), .B1(new_n1071), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1102), .B1(new_n1125), .B2(KEYINPUT57), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n977), .B1(new_n1125), .B2(KEYINPUT57), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT57), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1049), .A2(new_n1053), .A3(new_n1058), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1055), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1067), .B1(new_n1134), .B2(new_n1068), .ZN(new_n1135));
  OAI211_X1 g0935(.A(KEYINPUT122), .B(new_n1128), .C1(new_n1131), .C2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1126), .A2(new_n1127), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n729), .A2(G58), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n795), .B2(new_n748), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n386), .A2(new_n260), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n759), .B2(G77), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n903), .A2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n465), .B2(new_n742), .C1(new_n574), .C2(new_n745), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n459), .A2(new_n734), .B1(new_n735), .B2(new_n341), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(G50), .B1(new_n246), .B2(new_n260), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1145), .A2(KEYINPUT58), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n759), .A2(new_n1086), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n805), .B2(new_n738), .C1(new_n745), .C2(new_n1094), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n801), .A2(new_n734), .B1(new_n735), .B2(new_n908), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G128), .C2(new_n741), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n246), .B(new_n260), .C1(new_n728), .C2(new_n750), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G124), .B2(new_n754), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT59), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n1151), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1147), .B1(KEYINPUT58), .B2(new_n1145), .C1(new_n1153), .C2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n714), .B1(new_n1158), .B2(KEYINPUT119), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(KEYINPUT119), .B2(new_n1158), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT120), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n709), .B(new_n1161), .C1(new_n743), .C2(new_n787), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1109), .A2(new_n711), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1131), .B2(new_n933), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1137), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(KEYINPUT123), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(KEYINPUT123), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(G375));
  INV_X1    g0970(.A(new_n1065), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(new_n1124), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1172), .A2(new_n957), .A3(new_n1068), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n710), .B1(G68), .B2(new_n1074), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT124), .Z(new_n1175));
  OAI221_X1 g0975(.A(new_n249), .B1(new_n993), .B2(new_n731), .C1(new_n738), .C2(new_n743), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n742), .A2(new_n908), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G132), .C2(new_n744), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G150), .A2(new_n917), .B1(new_n918), .B2(new_n1086), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n754), .A2(G128), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1178), .A2(new_n1138), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n742), .A2(new_n795), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n744), .A2(G294), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n386), .B1(new_n731), .B2(new_n459), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n991), .A4(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G116), .A2(new_n918), .B1(new_n917), .B2(new_n469), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n754), .A2(G303), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n907), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1181), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1175), .B1(new_n767), .B2(new_n1189), .C1(new_n1046), .C2(new_n712), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1065), .B2(new_n933), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1173), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(G381));
  OAI21_X1  g0993(.A(new_n1100), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n979), .A2(new_n774), .A3(new_n1010), .ZN(new_n1195));
  OR4_X1    g0995(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1195), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1194), .A2(G387), .A3(new_n1196), .ZN(G407));
  OAI211_X1 g0997(.A(G407), .B(G213), .C1(G343), .C2(new_n1194), .ZN(G409));
  INV_X1    g0998(.A(G390), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(G393), .A2(G396), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(G387), .A2(new_n1199), .A3(new_n1195), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G387), .A2(new_n1199), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT126), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(new_n1195), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n975), .B2(G390), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1201), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(G387), .A2(new_n1204), .A3(new_n1199), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT61), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n639), .A2(G213), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1137), .A2(G378), .A3(new_n1166), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1131), .A2(new_n1135), .A3(new_n957), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1100), .B1(new_n1165), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(G384), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1069), .A2(new_n662), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT60), .B1(new_n1171), .B2(new_n1124), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT60), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1172), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1217), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1216), .B1(new_n1221), .B2(new_n1191), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1218), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1068), .A2(new_n977), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1191), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(G384), .A3(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1210), .A2(KEYINPUT125), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1222), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1211), .A2(G2897), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1229), .B(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT63), .B1(new_n1215), .B2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1215), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT63), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1209), .B(new_n1235), .C1(new_n1236), .C2(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1210), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1231), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1215), .A2(new_n1243), .A3(new_n1233), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(KEYINPUT127), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1208), .ZN(new_n1246));
  AND4_X1   g1046(.A1(new_n1243), .A2(new_n1238), .A3(new_n1210), .A4(new_n1233), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1215), .B2(new_n1231), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT127), .B1(new_n1250), .B2(new_n1242), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1237), .B1(new_n1246), .B2(new_n1251), .ZN(G405));
  OR2_X1    g1052(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1207), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n1233), .A3(new_n1254), .A4(new_n1201), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1233), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1194), .B1(new_n1100), .B2(new_n1167), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1258), .B(new_n1259), .ZN(G402));
endmodule


