

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n715), .A2(n714), .ZN(n755) );
  NOR2_X1 U552 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U553 ( .A(n525), .B(KEYINPUT0), .ZN(n630) );
  NOR2_X1 U554 ( .A1(n630), .A2(n531), .ZN(n519) );
  XOR2_X1 U555 ( .A(n752), .B(KEYINPUT31), .Z(n520) );
  OR2_X1 U556 ( .A1(n745), .A2(G301), .ZN(n521) );
  AND2_X1 U557 ( .A1(n720), .A2(n719), .ZN(n724) );
  INV_X1 U558 ( .A(n755), .ZN(n741) );
  NAND2_X1 U559 ( .A1(n764), .A2(G286), .ZN(n754) );
  NOR2_X1 U560 ( .A1(n798), .A2(n797), .ZN(n800) );
  INV_X1 U561 ( .A(G543), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n570), .A2(n569), .ZN(n925) );
  XOR2_X1 U563 ( .A(KEYINPUT4), .B(KEYINPUT77), .Z(n523) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U565 ( .A1(G89), .A2(n639), .ZN(n522) );
  XNOR2_X1 U566 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U567 ( .A(KEYINPUT76), .B(n524), .ZN(n527) );
  INV_X1 U568 ( .A(G651), .ZN(n531) );
  NAND2_X1 U569 ( .A1(n519), .A2(G76), .ZN(n526) );
  NAND2_X1 U570 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U571 ( .A(n528), .B(KEYINPUT5), .ZN(n537) );
  NOR2_X1 U572 ( .A1(G651), .A2(n630), .ZN(n529) );
  XNOR2_X1 U573 ( .A(KEYINPUT64), .B(n529), .ZN(n643) );
  NAND2_X1 U574 ( .A1(G51), .A2(n643), .ZN(n530) );
  XNOR2_X1 U575 ( .A(n530), .B(KEYINPUT78), .ZN(n534) );
  NOR2_X1 U576 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X2 U577 ( .A(KEYINPUT1), .B(n532), .Z(n642) );
  NAND2_X1 U578 ( .A1(G63), .A2(n642), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n535), .Z(n536) );
  NAND2_X1 U581 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U582 ( .A(n538), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .ZN(n539) );
  XNOR2_X1 U584 ( .A(n539), .B(KEYINPUT79), .ZN(G286) );
  XNOR2_X1 U585 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n541) );
  NOR2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  XNOR2_X2 U587 ( .A(n541), .B(n540), .ZN(n867) );
  NAND2_X1 U588 ( .A1(n867), .A2(G137), .ZN(n544) );
  INV_X1 U589 ( .A(G2105), .ZN(n545) );
  AND2_X4 U590 ( .A1(n545), .A2(G2104), .ZN(n869) );
  NAND2_X1 U591 ( .A1(G101), .A2(n869), .ZN(n542) );
  XOR2_X1 U592 ( .A(n542), .B(KEYINPUT23), .Z(n543) );
  NAND2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n549) );
  NOR2_X1 U594 ( .A1(G2104), .A2(n545), .ZN(n873) );
  NAND2_X1 U595 ( .A1(G125), .A2(n873), .ZN(n547) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U597 ( .A1(G113), .A2(n874), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U599 ( .A1(n549), .A2(n548), .ZN(G160) );
  NAND2_X1 U600 ( .A1(n642), .A2(G64), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G52), .A2(n643), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n557) );
  NAND2_X1 U603 ( .A1(G90), .A2(n639), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G77), .A2(n519), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U606 ( .A(KEYINPUT67), .B(n554), .ZN(n555) );
  XNOR2_X1 U607 ( .A(KEYINPUT9), .B(n555), .ZN(n556) );
  NOR2_X1 U608 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U609 ( .A(KEYINPUT68), .B(n558), .ZN(G171) );
  INV_X1 U610 ( .A(G171), .ZN(G301) );
  AND2_X1 U611 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U616 ( .A(G223), .ZN(n817) );
  NAND2_X1 U617 ( .A1(n817), .A2(G567), .ZN(n560) );
  XOR2_X1 U618 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U619 ( .A1(G68), .A2(n519), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n639), .A2(G81), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT12), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT13), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G43), .A2(n643), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U626 ( .A1(G56), .A2(n642), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n567), .B(KEYINPUT71), .ZN(n568) );
  XNOR2_X1 U628 ( .A(n568), .B(KEYINPUT14), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n925), .A2(G860), .ZN(G153) );
  INV_X1 U630 ( .A(G868), .ZN(n596) );
  NOR2_X1 U631 ( .A1(n596), .A2(G171), .ZN(n571) );
  XOR2_X1 U632 ( .A(n571), .B(KEYINPUT72), .Z(n583) );
  NAND2_X1 U633 ( .A1(G79), .A2(n519), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n572), .B(KEYINPUT74), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G92), .A2(n639), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G54), .A2(n643), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G66), .A2(n642), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT73), .B(n575), .ZN(n576) );
  NOR2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n580) );
  XNOR2_X2 U643 ( .A(n581), .B(n580), .ZN(n916) );
  INV_X1 U644 ( .A(n916), .ZN(n725) );
  NAND2_X1 U645 ( .A1(n596), .A2(n725), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U647 ( .A1(G91), .A2(n639), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G78), .A2(n519), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G65), .A2(n642), .ZN(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT69), .B(n586), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G53), .A2(n643), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(G299) );
  NOR2_X1 U655 ( .A1(G286), .A2(n596), .ZN(n592) );
  NOR2_X1 U656 ( .A1(G868), .A2(G299), .ZN(n591) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U658 ( .A(G860), .ZN(n612) );
  NAND2_X1 U659 ( .A1(n612), .A2(G559), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n593), .A2(n916), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U662 ( .A1(G559), .A2(n596), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n916), .A2(n595), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n925), .A2(n596), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U666 ( .A(KEYINPUT80), .B(n599), .Z(G282) );
  NAND2_X1 U667 ( .A1(G123), .A2(n873), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT18), .B(n600), .Z(n601) );
  XNOR2_X1 U669 ( .A(n601), .B(KEYINPUT81), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G111), .A2(n874), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G135), .A2(n867), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G99), .A2(n869), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n965) );
  XNOR2_X1 U676 ( .A(n965), .B(G2096), .ZN(n608) );
  XNOR2_X1 U677 ( .A(n608), .B(KEYINPUT82), .ZN(n610) );
  INV_X1 U678 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G559), .A2(n916), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n611), .B(n925), .ZN(n657) );
  NAND2_X1 U682 ( .A1(n612), .A2(n657), .ZN(n619) );
  NAND2_X1 U683 ( .A1(n642), .A2(G67), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G55), .A2(n643), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U686 ( .A1(G93), .A2(n639), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G80), .A2(n519), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n659) );
  XOR2_X1 U690 ( .A(n619), .B(n659), .Z(G145) );
  NAND2_X1 U691 ( .A1(G86), .A2(n639), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G48), .A2(n643), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n519), .A2(G73), .ZN(n622) );
  XOR2_X1 U695 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n642), .A2(G61), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U699 ( .A1(G651), .A2(G74), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G49), .A2(n643), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n642), .A2(n629), .ZN(n632) );
  NAND2_X1 U703 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G88), .A2(n639), .ZN(n634) );
  NAND2_X1 U706 ( .A1(G75), .A2(n519), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n642), .A2(G62), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G50), .A2(n643), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G85), .A2(n639), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G72), .A2(n519), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n642), .A2(G60), .ZN(n645) );
  NAND2_X1 U716 ( .A1(G47), .A2(n643), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(n648), .Z(G290) );
  XNOR2_X1 U720 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n650) );
  XNOR2_X1 U721 ( .A(G288), .B(KEYINPUT85), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U723 ( .A(n651), .B(KEYINPUT83), .Z(n653) );
  XNOR2_X1 U724 ( .A(G166), .B(n659), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U726 ( .A(G305), .B(n654), .ZN(n656) );
  INV_X1 U727 ( .A(G299), .ZN(n909) );
  XNOR2_X1 U728 ( .A(G290), .B(n909), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n656), .B(n655), .ZN(n885) );
  XNOR2_X1 U730 ( .A(n657), .B(n885), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n658), .A2(G868), .ZN(n661) );
  OR2_X1 U732 ( .A1(G868), .A2(n659), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U740 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  NOR2_X1 U741 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U742 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U743 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U744 ( .A1(G96), .A2(n668), .ZN(n822) );
  AND2_X1 U745 ( .A1(G2106), .A2(n822), .ZN(n673) );
  NAND2_X1 U746 ( .A1(G108), .A2(G120), .ZN(n669) );
  NOR2_X1 U747 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U748 ( .A1(G69), .A2(n670), .ZN(n821) );
  NAND2_X1 U749 ( .A1(G567), .A2(n821), .ZN(n671) );
  XOR2_X1 U750 ( .A(KEYINPUT86), .B(n671), .Z(n672) );
  NOR2_X1 U751 ( .A1(n673), .A2(n672), .ZN(G319) );
  INV_X1 U752 ( .A(G319), .ZN(n675) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n674) );
  NOR2_X1 U754 ( .A1(n675), .A2(n674), .ZN(n820) );
  NAND2_X1 U755 ( .A1(n820), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G138), .A2(n867), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G102), .A2(n869), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U759 ( .A1(G126), .A2(n873), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G114), .A2(n874), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U762 ( .A1(n681), .A2(n680), .ZN(G164) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n714) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n812) );
  XNOR2_X1 U767 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NAND2_X1 U768 ( .A1(G140), .A2(n867), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G104), .A2(n869), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U771 ( .A(KEYINPUT34), .B(n684), .ZN(n689) );
  NAND2_X1 U772 ( .A1(G128), .A2(n873), .ZN(n686) );
  NAND2_X1 U773 ( .A1(G116), .A2(n874), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U775 ( .A(KEYINPUT35), .B(n687), .Z(n688) );
  NOR2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U777 ( .A(KEYINPUT36), .B(n690), .ZN(n882) );
  NOR2_X1 U778 ( .A1(n810), .A2(n882), .ZN(n967) );
  NAND2_X1 U779 ( .A1(n812), .A2(n967), .ZN(n691) );
  XOR2_X1 U780 ( .A(KEYINPUT87), .B(n691), .Z(n808) );
  NAND2_X1 U781 ( .A1(G105), .A2(n869), .ZN(n692) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n692), .Z(n697) );
  NAND2_X1 U783 ( .A1(G129), .A2(n873), .ZN(n694) );
  NAND2_X1 U784 ( .A1(G117), .A2(n874), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U786 ( .A(KEYINPUT89), .B(n695), .Z(n696) );
  NOR2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n867), .A2(G141), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n864) );
  NAND2_X1 U790 ( .A1(G1996), .A2(n864), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n700), .B(KEYINPUT90), .ZN(n709) );
  NAND2_X1 U792 ( .A1(G95), .A2(n869), .ZN(n702) );
  NAND2_X1 U793 ( .A1(G107), .A2(n874), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n867), .A2(G131), .ZN(n703) );
  XOR2_X1 U796 ( .A(KEYINPUT88), .B(n703), .Z(n704) );
  NOR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n873), .A2(G119), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n858) );
  NAND2_X1 U800 ( .A1(G1991), .A2(n858), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U802 ( .A(KEYINPUT91), .B(n710), .ZN(n977) );
  INV_X1 U803 ( .A(n977), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n711), .A2(n812), .ZN(n801) );
  NAND2_X1 U805 ( .A1(n808), .A2(n801), .ZN(n712) );
  XNOR2_X1 U806 ( .A(n712), .B(KEYINPUT92), .ZN(n798) );
  XNOR2_X1 U807 ( .A(G1981), .B(G305), .ZN(n929) );
  XNOR2_X1 U808 ( .A(n713), .B(KEYINPUT93), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n741), .A2(G1348), .ZN(n717) );
  NOR2_X1 U810 ( .A1(G2067), .A2(n755), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n726) );
  NAND2_X1 U812 ( .A1(n725), .A2(n726), .ZN(n720) );
  NAND2_X1 U813 ( .A1(G1996), .A2(n741), .ZN(n718) );
  XNOR2_X1 U814 ( .A(KEYINPUT26), .B(n718), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n755), .A2(G1341), .ZN(n721) );
  XNOR2_X1 U816 ( .A(n721), .B(KEYINPUT94), .ZN(n722) );
  AND2_X1 U817 ( .A1(n722), .A2(n925), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n728) );
  OR2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U821 ( .A(KEYINPUT95), .B(n729), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n741), .A2(G2072), .ZN(n730) );
  XNOR2_X1 U823 ( .A(n730), .B(KEYINPUT27), .ZN(n732) );
  AND2_X1 U824 ( .A1(G1956), .A2(n755), .ZN(n731) );
  NOR2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n735), .A2(n909), .ZN(n733) );
  NAND2_X1 U827 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n735), .A2(n909), .ZN(n736) );
  XOR2_X1 U829 ( .A(n736), .B(KEYINPUT28), .Z(n737) );
  NAND2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U831 ( .A(n739), .B(KEYINPUT29), .ZN(n740) );
  INV_X1 U832 ( .A(n740), .ZN(n744) );
  NAND2_X1 U833 ( .A1(G1961), .A2(n755), .ZN(n743) );
  XOR2_X1 U834 ( .A(KEYINPUT25), .B(G2078), .Z(n942) );
  NAND2_X1 U835 ( .A1(n741), .A2(n942), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n744), .A2(n521), .ZN(n753) );
  NAND2_X1 U838 ( .A1(G301), .A2(n745), .ZN(n746) );
  XOR2_X1 U839 ( .A(KEYINPUT96), .B(n746), .Z(n751) );
  NAND2_X1 U840 ( .A1(G8), .A2(n755), .ZN(n792) );
  NOR2_X1 U841 ( .A1(G1966), .A2(n792), .ZN(n766) );
  NOR2_X1 U842 ( .A1(G2084), .A2(n755), .ZN(n767) );
  NOR2_X1 U843 ( .A1(n766), .A2(n767), .ZN(n747) );
  NAND2_X1 U844 ( .A1(G8), .A2(n747), .ZN(n748) );
  XNOR2_X1 U845 ( .A(KEYINPUT30), .B(n748), .ZN(n749) );
  NOR2_X1 U846 ( .A1(G168), .A2(n749), .ZN(n750) );
  NOR2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U848 ( .A1(n753), .A2(n520), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n754), .B(KEYINPUT98), .ZN(n761) );
  NOR2_X1 U850 ( .A1(G1971), .A2(n792), .ZN(n757) );
  NOR2_X1 U851 ( .A1(G2090), .A2(n755), .ZN(n756) );
  NOR2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U853 ( .A1(n758), .A2(G303), .ZN(n759) );
  XOR2_X1 U854 ( .A(KEYINPUT99), .B(n759), .Z(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n762), .A2(G8), .ZN(n763) );
  XNOR2_X1 U857 ( .A(n763), .B(KEYINPUT32), .ZN(n772) );
  INV_X1 U858 ( .A(n764), .ZN(n765) );
  NOR2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U860 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U862 ( .A(KEYINPUT97), .B(n770), .Z(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n790) );
  NOR2_X1 U864 ( .A1(G288), .A2(G1976), .ZN(n773) );
  XNOR2_X1 U865 ( .A(n773), .B(KEYINPUT100), .ZN(n781) );
  NOR2_X1 U866 ( .A1(G1971), .A2(G303), .ZN(n774) );
  NOR2_X1 U867 ( .A1(n781), .A2(n774), .ZN(n913) );
  NAND2_X1 U868 ( .A1(n790), .A2(n913), .ZN(n775) );
  XNOR2_X1 U869 ( .A(n775), .B(KEYINPUT101), .ZN(n778) );
  NAND2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n912) );
  INV_X1 U871 ( .A(n792), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n912), .A2(n776), .ZN(n777) );
  NOR2_X1 U873 ( .A1(KEYINPUT33), .A2(n779), .ZN(n780) );
  NOR2_X1 U874 ( .A1(n929), .A2(n780), .ZN(n785) );
  INV_X1 U875 ( .A(n781), .ZN(n782) );
  NOR2_X1 U876 ( .A1(n792), .A2(n782), .ZN(n783) );
  NAND2_X1 U877 ( .A1(KEYINPUT33), .A2(n783), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n796) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XOR2_X1 U880 ( .A(n786), .B(KEYINPUT24), .Z(n787) );
  OR2_X1 U881 ( .A1(n792), .A2(n787), .ZN(n794) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G8), .A2(n788), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  AND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n795) );
  AND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U888 ( .A(G1986), .B(G290), .ZN(n918) );
  NAND2_X1 U889 ( .A1(n918), .A2(n812), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n815) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n864), .ZN(n960) );
  INV_X1 U892 ( .A(n801), .ZN(n805) );
  NOR2_X1 U893 ( .A1(n858), .A2(G1991), .ZN(n802) );
  XNOR2_X1 U894 ( .A(n802), .B(KEYINPUT102), .ZN(n966) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n966), .A2(n803), .ZN(n804) );
  NOR2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U898 ( .A1(n960), .A2(n806), .ZN(n807) );
  XNOR2_X1 U899 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n810), .A2(n882), .ZN(n962) );
  NAND2_X1 U902 ( .A1(n811), .A2(n962), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U905 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U908 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(G188) );
  INV_X1 U912 ( .A(G120), .ZN(G236) );
  INV_X1 U913 ( .A(G108), .ZN(G238) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  XOR2_X1 U918 ( .A(G2100), .B(G2096), .Z(n824) );
  XNOR2_X1 U919 ( .A(KEYINPUT42), .B(G2678), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT43), .B(G2090), .Z(n826) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2072), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U924 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U925 ( .A(G2078), .B(G2084), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(G227) );
  XNOR2_X1 U927 ( .A(G1996), .B(KEYINPUT106), .ZN(n840) );
  XOR2_X1 U928 ( .A(G1981), .B(G1961), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1991), .B(G1966), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U931 ( .A(G1976), .B(G1971), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1986), .B(G1956), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2474), .B(KEYINPUT41), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(G229) );
  NAND2_X1 U938 ( .A1(G100), .A2(n869), .ZN(n842) );
  NAND2_X1 U939 ( .A1(G112), .A2(n874), .ZN(n841) );
  NAND2_X1 U940 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n843), .B(KEYINPUT107), .ZN(n845) );
  NAND2_X1 U942 ( .A1(G136), .A2(n867), .ZN(n844) );
  NAND2_X1 U943 ( .A1(n845), .A2(n844), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n873), .A2(G124), .ZN(n846) );
  XOR2_X1 U945 ( .A(KEYINPUT44), .B(n846), .Z(n847) );
  NOR2_X1 U946 ( .A1(n848), .A2(n847), .ZN(G162) );
  NAND2_X1 U947 ( .A1(G130), .A2(n873), .ZN(n850) );
  NAND2_X1 U948 ( .A1(G118), .A2(n874), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT108), .B(n851), .ZN(n857) );
  NAND2_X1 U951 ( .A1(n869), .A2(G106), .ZN(n852) );
  XOR2_X1 U952 ( .A(KEYINPUT109), .B(n852), .Z(n854) );
  NAND2_X1 U953 ( .A1(n867), .A2(G142), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(n855), .B(KEYINPUT45), .Z(n856) );
  NOR2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U958 ( .A(n860), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U959 ( .A(G164), .B(KEYINPUT46), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U961 ( .A(G162), .B(n965), .Z(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(n881) );
  NAND2_X1 U964 ( .A1(n867), .A2(G139), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT110), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G103), .A2(n869), .ZN(n870) );
  NAND2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT111), .B(n872), .Z(n879) );
  NAND2_X1 U969 ( .A1(G127), .A2(n873), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G115), .A2(n874), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U973 ( .A1(n879), .A2(n878), .ZN(n970) );
  XNOR2_X1 U974 ( .A(G160), .B(n970), .ZN(n880) );
  XNOR2_X1 U975 ( .A(n881), .B(n880), .ZN(n883) );
  XOR2_X1 U976 ( .A(n883), .B(n882), .Z(n884) );
  NOR2_X1 U977 ( .A1(G37), .A2(n884), .ZN(G395) );
  XOR2_X1 U978 ( .A(KEYINPUT112), .B(n885), .Z(n887) );
  XNOR2_X1 U979 ( .A(n925), .B(G286), .ZN(n886) );
  XNOR2_X1 U980 ( .A(n887), .B(n886), .ZN(n889) );
  XOR2_X1 U981 ( .A(n916), .B(G301), .Z(n888) );
  XNOR2_X1 U982 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U983 ( .A1(G37), .A2(n890), .ZN(G397) );
  XOR2_X1 U984 ( .A(G2451), .B(KEYINPUT104), .Z(n892) );
  XNOR2_X1 U985 ( .A(G2443), .B(G2446), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U987 ( .A(n893), .B(KEYINPUT105), .Z(n895) );
  XNOR2_X1 U988 ( .A(G1348), .B(G1341), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U990 ( .A(G2435), .B(G2438), .Z(n897) );
  XNOR2_X1 U991 ( .A(G2454), .B(G2430), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U994 ( .A(G2427), .B(KEYINPUT103), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U996 ( .A1(n902), .A2(G14), .ZN(n908) );
  NAND2_X1 U997 ( .A1(G319), .A2(n908), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(n908), .ZN(G401) );
  XNOR2_X1 U1005 ( .A(n909), .B(G1956), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G1971), .A2(G303), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n920) );
  XOR2_X1 U1010 ( .A(G1348), .B(n916), .Z(n917) );
  NOR2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1012 ( .A1(n920), .A2(n919), .ZN(n923) );
  XOR2_X1 U1013 ( .A(G1961), .B(G301), .Z(n921) );
  XNOR2_X1 U1014 ( .A(KEYINPUT119), .B(n921), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(KEYINPUT120), .B(n924), .ZN(n927) );
  XNOR2_X1 U1017 ( .A(n925), .B(G1341), .ZN(n926) );
  NAND2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n934) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n928) );
  XNOR2_X1 U1020 ( .A(n928), .B(KEYINPUT117), .ZN(n930) );
  NOR2_X1 U1021 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1022 ( .A(KEYINPUT118), .B(n931), .ZN(n932) );
  XNOR2_X1 U1023 ( .A(KEYINPUT57), .B(n932), .ZN(n933) );
  NOR2_X1 U1024 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(KEYINPUT121), .B(n935), .ZN(n938) );
  XNOR2_X1 U1026 ( .A(G16), .B(KEYINPUT116), .ZN(n936) );
  XNOR2_X1 U1027 ( .A(n936), .B(KEYINPUT56), .ZN(n937) );
  NAND2_X1 U1028 ( .A1(n938), .A2(n937), .ZN(n988) );
  XOR2_X1 U1029 ( .A(G1991), .B(G25), .Z(n939) );
  NAND2_X1 U1030 ( .A1(n939), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(G1996), .B(G32), .ZN(n944) );
  XNOR2_X1 U1035 ( .A(G27), .B(n942), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1039 ( .A(KEYINPUT53), .B(n949), .Z(n952) );
  XOR2_X1 U1040 ( .A(KEYINPUT54), .B(G34), .Z(n950) );
  XNOR2_X1 U1041 ( .A(G2084), .B(n950), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n953) );
  NOR2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(KEYINPUT55), .B(KEYINPUT113), .ZN(n981) );
  XOR2_X1 U1046 ( .A(n955), .B(n981), .Z(n957) );
  XNOR2_X1 U1047 ( .A(G29), .B(KEYINPUT115), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n958), .ZN(n986) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n961), .Z(n963) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n979) );
  XOR2_X1 U1054 ( .A(G2084), .B(G160), .Z(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n969) );
  NOR2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1057 ( .A1(n969), .A2(n968), .ZN(n975) );
  XOR2_X1 U1058 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1059 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n973), .Z(n974) );
  NOR2_X1 U1062 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1063 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1064 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1065 ( .A(KEYINPUT52), .B(n980), .ZN(n982) );
  NAND2_X1 U1066 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1067 ( .A1(n983), .A2(G29), .ZN(n984) );
  XOR2_X1 U1068 ( .A(KEYINPUT114), .B(n984), .Z(n985) );
  NOR2_X1 U1069 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1070 ( .A1(n988), .A2(n987), .ZN(n1015) );
  XOR2_X1 U1071 ( .A(G1976), .B(G23), .Z(n990) );
  XOR2_X1 U1072 ( .A(G1971), .B(G22), .Z(n989) );
  NAND2_X1 U1073 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1074 ( .A(G24), .B(G1986), .ZN(n991) );
  NOR2_X1 U1075 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1076 ( .A(KEYINPUT58), .B(n993), .Z(n1011) );
  XOR2_X1 U1077 ( .A(G1961), .B(G5), .Z(n1006) );
  XOR2_X1 U1078 ( .A(G1348), .B(KEYINPUT59), .Z(n994) );
  XNOR2_X1 U1079 ( .A(G4), .B(n994), .ZN(n1003) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n995), .B(KEYINPUT122), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G6), .B(G1981), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(KEYINPUT123), .B(n998), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(KEYINPUT124), .B(n1001), .Z(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(KEYINPUT60), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G21), .B(G1966), .ZN(n1007) );
  NOR2_X1 U1092 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1094 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1012), .Z(n1013) );
  NOR2_X1 U1096 ( .A1(G16), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1097 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(n1016), .B(KEYINPUT62), .ZN(G311) );
  XOR2_X1 U1099 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

