//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT18), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT83), .B(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G29gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(KEYINPUT15), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n219), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n220), .A2(KEYINPUT82), .B1(new_n225), .B2(KEYINPUT14), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n226), .A2(new_n228), .B1(G29gat), .B2(new_n212), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT84), .B1(new_n229), .B2(new_n216), .ZN(new_n230));
  NOR3_X1   g029(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n221), .B1(new_n231), .B2(new_n227), .ZN(new_n232));
  INV_X1    g031(.A(new_n228), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n213), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235));
  INV_X1    g034(.A(new_n216), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n224), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT16), .ZN(new_n240));
  INV_X1    g039(.A(G22gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G15gat), .ZN(new_n242));
  INV_X1    g041(.A(G15gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G22gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(G1gat), .B1(new_n242), .B2(new_n244), .ZN(new_n247));
  OAI21_X1  g046(.A(G8gat), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT85), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(G8gat), .C1(new_n246), .C2(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(KEYINPUT86), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n247), .A2(G8gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n249), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n211), .B1(new_n238), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n215), .A2(new_n223), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n220), .A2(KEYINPUT82), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n221), .A3(new_n228), .ZN(new_n261));
  AOI211_X1 g060(.A(KEYINPUT84), .B(new_n216), .C1(new_n261), .C2(new_n213), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT17), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT17), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n266), .B(new_n259), .C1(new_n262), .C2(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n258), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n256), .A3(new_n251), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n211), .B(new_n270), .C1(new_n265), .C2(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n210), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n264), .B(new_n257), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n207), .B(KEYINPUT13), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n230), .A2(new_n237), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n266), .B1(new_n279), .B2(new_n259), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT17), .B(new_n224), .C1(new_n230), .C2(new_n237), .ZN(new_n281));
  OAI211_X1 g080(.A(KEYINPUT87), .B(new_n257), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n270), .B1(new_n265), .B2(new_n267), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n258), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT18), .B1(new_n284), .B2(new_n207), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n206), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n273), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n206), .B1(new_n287), .B2(new_n274), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n257), .B1(new_n280), .B2(new_n281), .ZN(new_n289));
  INV_X1    g088(.A(new_n258), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n208), .B1(new_n291), .B2(new_n282), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n272), .B(new_n288), .C1(new_n292), .C2(KEYINPUT18), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n296));
  XOR2_X1   g095(.A(G1gat), .B(G29gat), .Z(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  INV_X1    g106(.A(G162gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G141gat), .B(G148gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n306), .B(new_n309), .C1(new_n310), .C2(KEYINPUT2), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .A4(G141gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n306), .B1(new_n309), .B2(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT71), .B1(new_n312), .B2(G141gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT70), .B(G148gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(G141gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n311), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(KEYINPUT1), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(new_n324), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n323), .B(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n311), .C1(new_n319), .C2(new_n322), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n331), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n313), .A2(new_n315), .A3(G141gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n320), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n317), .A3(new_n318), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n337), .B1(new_n343), .B2(new_n311), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT72), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n323), .A2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n331), .A4(new_n338), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n334), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n327), .A2(new_n330), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n343), .A4(new_n311), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n323), .A2(new_n331), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT4), .B1(new_n323), .B2(new_n331), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n336), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n352), .A2(new_n357), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n349), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n304), .B(new_n305), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n349), .A2(new_n358), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT5), .A3(new_n335), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n360), .A3(new_n361), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n365), .A2(new_n366), .A3(new_n303), .A4(new_n302), .ZN(new_n367));
  AND2_X1   g166(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G169gat), .ZN(new_n378));
  INV_X1    g177(.A(G176gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT23), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n377), .B(new_n380), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n368), .A2(new_n370), .B1(G169gat), .B2(G176gat), .ZN(new_n382));
  OR2_X1    g181(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(G190gat), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT64), .A4(new_n373), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n373), .A4(new_n380), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT27), .B(G183gat), .ZN(new_n390));
  OR2_X1    g189(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n391));
  NAND2_X1  g190(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n390), .A2(new_n370), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G183gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT27), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G183gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n397), .A3(new_n370), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n392), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n393), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT66), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n403), .A2(KEYINPUT26), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(KEYINPUT26), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n375), .A3(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n381), .A2(new_n389), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G226gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  OAI22_X1  g208(.A1(new_n407), .A2(KEYINPUT29), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G211gat), .A2(G218gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(G211gat), .A2(G218gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(G197gat), .A2(G204gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(G197gat), .A2(G204gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G211gat), .B(G218gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G197gat), .B(G204gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n418), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n423), .A3(KEYINPUT69), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n414), .B(new_n425), .C1(new_n417), .C2(new_n418), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n406), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n387), .B1(new_n388), .B2(new_n386), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n408), .A2(new_n409), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n410), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n410), .B2(new_n433), .ZN(new_n435));
  XNOR2_X1  g234(.A(G8gat), .B(G36gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(KEYINPUT37), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT38), .ZN(new_n440));
  OR3_X1    g239(.A1(new_n434), .A2(new_n435), .A3(new_n440), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n434), .A2(new_n435), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n363), .A2(new_n367), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  INV_X1    g243(.A(G228gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n409), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n419), .A2(new_n423), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT29), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n450), .A2(new_n337), .B1(new_n343), .B2(new_n311), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n338), .A2(new_n449), .B1(new_n426), .B2(new_n424), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT77), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n338), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n427), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n419), .B2(new_n423), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n323), .B1(new_n458), .B2(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT77), .A3(new_n447), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n424), .A2(new_n449), .A3(new_n426), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n449), .A4(new_n426), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n337), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n323), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n447), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n462), .A2(new_n241), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n241), .B1(new_n462), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n444), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT77), .B1(new_n460), .B2(new_n447), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n454), .B(new_n446), .C1(new_n457), .C2(new_n459), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G22gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n241), .A3(new_n470), .ZN(new_n479));
  INV_X1    g278(.A(new_n444), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n473), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n474), .B1(new_n473), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n443), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n345), .A2(new_n348), .B1(new_n352), .B2(new_n357), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n485), .A2(KEYINPUT39), .A3(new_n333), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT79), .B1(new_n486), .B2(new_n302), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n345), .A2(new_n348), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n361), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n334), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n301), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n485), .A2(new_n333), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT39), .B1(new_n332), .B2(new_n334), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT40), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT40), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n500), .B(new_n497), .C1(new_n487), .C2(new_n493), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n502));
  INV_X1    g301(.A(new_n427), .ZN(new_n503));
  INV_X1    g302(.A(new_n433), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n432), .B1(new_n431), .B2(new_n449), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n438), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n410), .A2(new_n433), .A3(new_n427), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT30), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n511), .B(new_n438), .C1(new_n434), .C2(new_n435), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n302), .B1(new_n359), .B2(new_n362), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n499), .A2(new_n501), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n296), .B1(new_n484), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n431), .A2(new_n331), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n407), .A2(new_n350), .ZN(new_n518));
  NAND2_X1  g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n381), .A2(new_n389), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n525), .A2(new_n350), .A3(new_n428), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n350), .B1(new_n525), .B2(new_n428), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT32), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT33), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT67), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G15gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n532), .B(KEYINPUT67), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n243), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n534), .A2(new_n536), .A3(G43gat), .ZN(new_n537));
  AOI21_X1  g336(.A(G43gat), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n529), .A2(new_n531), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n528), .B(KEYINPUT32), .C1(new_n541), .C2(new_n530), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT34), .B1(new_n520), .B2(new_n521), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n540), .B2(new_n542), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n523), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n519), .B1(new_n517), .B2(new_n518), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n539), .B1(new_n548), .B2(KEYINPUT33), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n542), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n543), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n540), .A2(new_n544), .A3(new_n542), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n522), .A3(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n547), .A2(new_n556), .A3(KEYINPUT36), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT36), .B1(new_n547), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n494), .A2(new_n498), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n500), .ZN(new_n561));
  INV_X1    g360(.A(new_n514), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n494), .A2(KEYINPUT40), .A3(new_n498), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n474), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n471), .A2(new_n472), .A3(new_n444), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n480), .B1(new_n478), .B2(new_n479), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n473), .A2(new_n474), .A3(new_n481), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n570), .A3(KEYINPUT80), .A4(new_n443), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n510), .A2(new_n512), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n363), .A2(new_n367), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT76), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT76), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n575), .A2(new_n569), .A3(new_n568), .A4(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n516), .A2(new_n559), .A3(new_n571), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n547), .A2(new_n556), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT76), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(new_n574), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT35), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n572), .ZN(new_n584));
  INV_X1    g383(.A(new_n573), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT35), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n570), .A3(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT81), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n578), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n295), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT88), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(KEYINPUT88), .A3(new_n595), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT90), .ZN(new_n603));
  NAND2_X1  g402(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n603), .B(G57gat), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n600), .B1(new_n594), .B2(new_n595), .ZN(new_n608));
  INV_X1    g407(.A(G57gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(G64gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT90), .B1(new_n612), .B2(G57gat), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n607), .B(new_n608), .C1(new_n611), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n602), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n257), .B1(new_n616), .B2(new_n615), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT91), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n621), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT92), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G85gat), .A2(G92gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT7), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(G85gat), .ZN(new_n640));
  INV_X1    g439(.A(G92gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G99gat), .B(G106gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n638), .A3(new_n642), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n645), .A2(KEYINPUT93), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT93), .B1(new_n645), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n268), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G190gat), .B(G218gat), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n650), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n654), .A2(new_n264), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n651), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n636), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n635), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n629), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n615), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n648), .B2(new_n649), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n645), .A2(new_n647), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n615), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n645), .A2(new_n602), .A3(new_n614), .A4(new_n647), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n665), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n665), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(new_n678));
  OR2_X1    g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n668), .A2(new_n672), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n664), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n674), .A2(new_n665), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n663), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n593), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n573), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n239), .ZN(G1324gat));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  NAND4_X1  g488(.A1(new_n593), .A2(new_n584), .A3(new_n685), .A4(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT95), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT94), .ZN(new_n696));
  OAI21_X1  g495(.A(G8gat), .B1(new_n686), .B2(new_n572), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(G1325gat));
  INV_X1    g497(.A(KEYINPUT96), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n557), .B2(new_n558), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT36), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n579), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n547), .A2(new_n556), .A3(KEYINPUT36), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(KEYINPUT96), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G15gat), .B1(new_n686), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n579), .A2(new_n243), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n686), .B2(new_n707), .ZN(G1326gat));
  INV_X1    g507(.A(new_n570), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n593), .A2(new_n709), .A3(new_n685), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT97), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n711), .B(new_n712), .Z(G1327gat));
  INV_X1    g512(.A(new_n662), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT44), .B1(new_n589), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n590), .A2(new_n592), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n662), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n684), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n628), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n295), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n585), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G29gat), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n721), .A2(new_n662), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n716), .A2(new_n294), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n573), .A2(G29gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n725), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n727), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n728), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n724), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT98), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n724), .A2(new_n735), .A3(new_n730), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1328gat));
  INV_X1    g536(.A(KEYINPUT99), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n212), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(new_n584), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n719), .A2(new_n584), .A3(new_n722), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n212), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1329gat));
  INV_X1    g544(.A(KEYINPUT100), .ZN(new_n746));
  INV_X1    g545(.A(new_n559), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n719), .A2(new_n746), .A3(new_n747), .A4(new_n722), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n578), .A2(new_n588), .A3(new_n591), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n591), .B1(new_n578), .B2(new_n588), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n718), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n589), .A2(new_n714), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n717), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n751), .A2(new_n747), .A3(new_n753), .A4(new_n722), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(new_n755), .A3(G43gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n579), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n593), .A2(new_n726), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n705), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n751), .A2(new_n763), .A3(new_n753), .A4(new_n722), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G43gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n759), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n762), .A2(KEYINPUT101), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT101), .ZN(new_n770));
  INV_X1    g569(.A(G43gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n754), .B2(KEYINPUT100), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n760), .B1(new_n772), .B2(new_n748), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT47), .B1(new_n765), .B2(new_n759), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n769), .A2(new_n775), .ZN(G1330gat));
  NAND3_X1  g575(.A1(new_n719), .A2(new_n709), .A3(new_n722), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G50gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n570), .A2(G50gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n731), .A2(new_n779), .B1(KEYINPUT102), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n780), .A2(KEYINPUT102), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1331gat));
  NOR3_X1   g583(.A1(new_n663), .A2(new_n294), .A3(new_n720), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n589), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n585), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G57gat), .ZN(G1332gat));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n584), .B1(new_n789), .B2(new_n612), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT103), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n612), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1333gat));
  NAND2_X1  g595(.A1(new_n786), .A2(new_n763), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n757), .A2(G71gat), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n797), .A2(G71gat), .B1(new_n786), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1334gat));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n709), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g602(.A1(new_n294), .A2(new_n629), .A3(new_n720), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n719), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G85gat), .B1(new_n805), .B2(new_n573), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n589), .A2(new_n295), .A3(new_n628), .A4(new_n714), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT51), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n585), .A2(new_n640), .A3(new_n684), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT51), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n720), .A2(G92gat), .A3(new_n572), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n719), .A2(new_n584), .A3(new_n804), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n813), .A2(new_n814), .B1(new_n815), .B2(G92gat), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n815), .A2(G92gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(KEYINPUT108), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n817), .A2(KEYINPUT108), .ZN(new_n820));
  INV_X1    g619(.A(new_n814), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n819), .B(new_n820), .C1(new_n808), .C2(new_n821), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n816), .A2(new_n817), .B1(new_n818), .B2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n805), .B2(new_n705), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n757), .A2(G99gat), .A3(new_n720), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n808), .B2(new_n825), .ZN(G1338gat));
  NOR3_X1   g625(.A1(new_n570), .A2(G106gat), .A3(new_n720), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n719), .A2(new_n709), .A3(new_n804), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n813), .A2(new_n827), .B1(new_n828), .B2(G106gat), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n828), .A2(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n827), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n808), .B2(new_n832), .ZN(new_n833));
  OAI22_X1  g632(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n833), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n668), .A2(new_n672), .A3(new_n665), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n681), .A2(new_n836), .A3(KEYINPUT54), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n678), .B1(new_n673), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(KEYINPUT55), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n683), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(new_n837), .B2(new_n839), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n282), .B(new_n208), .C1(new_n283), .C2(new_n258), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n273), .A2(new_n275), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n205), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n293), .A2(new_n684), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n294), .A2(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n293), .A2(new_n684), .A3(new_n847), .A4(KEYINPUT109), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n714), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n843), .A2(new_n661), .A3(new_n659), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n293), .A2(new_n847), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n835), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n848), .A2(new_n849), .ZN(new_n857));
  INV_X1    g656(.A(new_n206), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n207), .B1(new_n269), .B2(new_n271), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n209), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n276), .B1(new_n284), .B2(new_n210), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n272), .A2(new_n288), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n285), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n843), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n865), .A3(new_n851), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n855), .B1(new_n866), .B2(new_n662), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT110), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n856), .A2(new_n628), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n685), .A2(new_n295), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n580), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n573), .A3(new_n584), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n295), .A2(G113gat), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT112), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n294), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(KEYINPUT111), .A3(G113gat), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT111), .B1(new_n877), .B2(G113gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(G1340gat));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G120gat), .ZN(new_n882));
  XOR2_X1   g681(.A(KEYINPUT113), .B(G120gat), .Z(new_n883));
  NAND2_X1  g682(.A1(new_n873), .A2(new_n684), .ZN(new_n884));
  MUX2_X1   g683(.A(new_n882), .B(new_n883), .S(new_n884), .Z(G1341gat));
  NAND2_X1  g684(.A1(new_n873), .A2(new_n629), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g686(.A1(new_n873), .A2(new_n714), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n888), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(G134gat), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT56), .B1(new_n888), .B2(G134gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G1343gat));
  AOI21_X1  g691(.A(new_n570), .B1(new_n869), .B2(new_n870), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n559), .A2(new_n585), .A3(new_n572), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n714), .B1(new_n865), .B2(new_n848), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n628), .B1(new_n897), .B2(new_n855), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n870), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n709), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G141gat), .B1(new_n902), .B2(new_n295), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n573), .B1(new_n869), .B2(new_n870), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT114), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(KEYINPUT114), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n570), .B1(new_n700), .B2(new_n704), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n572), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n295), .A2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT58), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n903), .B(new_n914), .C1(new_n909), .C2(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1344gat));
  INV_X1    g715(.A(new_n909), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n321), .A3(new_n684), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n628), .B1(new_n867), .B2(KEYINPUT110), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n835), .B(new_n855), .C1(new_n866), .C2(new_n662), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n870), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n894), .B1(new_n922), .B2(new_n709), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n870), .B(new_n924), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT57), .B(new_n570), .C1(new_n925), .C2(new_n898), .ZN(new_n926));
  NOR4_X1   g725(.A1(new_n923), .A2(new_n926), .A3(new_n720), .A4(new_n896), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n312), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n919), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n902), .A2(new_n720), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(KEYINPUT59), .A3(new_n321), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n918), .B1(new_n931), .B2(new_n933), .ZN(G1345gat));
  OAI21_X1  g733(.A(G155gat), .B1(new_n902), .B2(new_n628), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n629), .A2(new_n307), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n909), .B2(new_n936), .ZN(G1346gat));
  OAI21_X1  g736(.A(G162gat), .B1(new_n902), .B2(new_n662), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n714), .A2(new_n308), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n909), .B2(new_n939), .ZN(G1347gat));
  INV_X1    g739(.A(new_n580), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n585), .A2(new_n572), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n378), .A3(new_n294), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(KEYINPUT117), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n922), .A2(new_n947), .A3(new_n941), .A4(new_n942), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n295), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n378), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n949), .A2(KEYINPUT118), .A3(new_n378), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n379), .A3(new_n684), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n720), .B1(new_n946), .B2(new_n948), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n379), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n944), .A2(new_n390), .A3(new_n629), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n628), .B1(new_n946), .B2(new_n948), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n394), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n947), .B1(new_n871), .B2(new_n942), .ZN(new_n964));
  INV_X1    g763(.A(new_n948), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n714), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n963), .B1(new_n966), .B2(G190gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n662), .B1(new_n946), .B2(new_n948), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(KEYINPUT120), .A3(new_n370), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n963), .A3(G190gat), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT120), .B1(new_n968), .B2(new_n370), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n944), .A2(new_n370), .A3(new_n714), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT119), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(G1351gat));
  NAND2_X1  g775(.A1(new_n907), .A2(new_n584), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n573), .B1(new_n977), .B2(KEYINPUT121), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT121), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n979), .B1(new_n907), .B2(new_n584), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n981), .A2(new_n922), .ZN(new_n982));
  INV_X1    g781(.A(G197gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n983), .A3(new_n294), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n705), .A2(new_n942), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT123), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT122), .B1(new_n923), .B2(new_n926), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n925), .A2(new_n898), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n894), .A3(new_n709), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n988), .B(new_n990), .C1(new_n893), .C2(new_n894), .ZN(new_n991));
  AOI211_X1 g790(.A(new_n295), .B(new_n986), .C1(new_n987), .C2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n993));
  OAI21_X1  g792(.A(G197gat), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n986), .B1(new_n987), .B2(new_n991), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(new_n993), .A3(new_n294), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n984), .B1(new_n994), .B2(new_n996), .ZN(G1352gat));
  AND2_X1   g796(.A1(new_n907), .A2(new_n584), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n585), .B1(new_n998), .B2(new_n979), .ZN(new_n999));
  INV_X1    g798(.A(new_n980), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n720), .A2(G204gat), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n999), .A2(new_n922), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n981), .A2(KEYINPUT125), .A3(new_n922), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(KEYINPUT126), .B1(new_n1006), .B2(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n1004), .A2(new_n1008), .A3(new_n1005), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n684), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(G204gat), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(G1353gat));
  INV_X1    g814(.A(G211gat), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n982), .A2(new_n1016), .A3(new_n629), .ZN(new_n1017));
  OR4_X1    g816(.A1(new_n628), .A2(new_n923), .A3(new_n926), .A4(new_n985), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(G1354gat));
  NAND2_X1  g820(.A1(new_n982), .A2(new_n714), .ZN(new_n1022));
  INV_X1    g821(.A(G218gat), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1024), .A2(KEYINPUT127), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1022), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1027));
  NOR2_X1   g826(.A1(new_n662), .A2(new_n1023), .ZN(new_n1028));
  AOI22_X1  g827(.A1(new_n1025), .A2(new_n1027), .B1(new_n995), .B2(new_n1028), .ZN(G1355gat));
endmodule


