

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818;

  OR2_X1 U369 ( .A1(n702), .A2(G902), .ZN(n481) );
  INV_X1 U370 ( .A(G113), .ZN(n710) );
  INV_X1 U371 ( .A(G122), .ZN(n730) );
  INV_X1 U372 ( .A(G953), .ZN(n623) );
  XNOR2_X1 U373 ( .A(n353), .B(n492), .ZN(n697) );
  BUF_X1 U374 ( .A(n618), .Z(n671) );
  AND2_X1 U375 ( .A1(n352), .A2(n376), .ZN(n347) );
  OR2_X1 U376 ( .A1(n440), .A2(KEYINPUT47), .ZN(n348) );
  INV_X1 U377 ( .A(n629), .ZN(n759) );
  XNOR2_X2 U378 ( .A(n535), .B(KEYINPUT33), .ZN(n776) );
  OR2_X2 U379 ( .A1(n354), .A2(G902), .ZN(n532) );
  NOR2_X1 U380 ( .A1(n708), .A2(n656), .ZN(n667) );
  XNOR2_X1 U381 ( .A(n475), .B(n474), .ZN(n723) );
  NOR2_X1 U382 ( .A1(n756), .A2(n412), .ZN(n485) );
  AND2_X1 U383 ( .A1(n686), .A2(n685), .ZN(n756) );
  XNOR2_X1 U384 ( .A(n359), .B(KEYINPUT45), .ZN(n684) );
  NOR2_X2 U385 ( .A1(n602), .A2(n469), .ZN(n363) );
  XNOR2_X1 U386 ( .A(n358), .B(n357), .ZN(n356) );
  NOR2_X1 U387 ( .A1(n645), .A2(n778), .ZN(n471) );
  INV_X1 U388 ( .A(n751), .ZN(n349) );
  OR2_X1 U389 ( .A1(n607), .A2(n563), .ZN(n377) );
  XNOR2_X1 U390 ( .A(n562), .B(n561), .ZN(n607) );
  NOR2_X1 U391 ( .A1(n366), .A2(G953), .ZN(n509) );
  INV_X1 U392 ( .A(G234), .ZN(n366) );
  INV_X1 U393 ( .A(G902), .ZN(n369) );
  NAND2_X1 U394 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U395 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U396 ( .A1(n391), .A2(n382), .ZN(n380) );
  AND2_X1 U397 ( .A1(n394), .A2(n392), .ZN(n389) );
  NAND2_X1 U398 ( .A1(n391), .A2(n390), .ZN(n388) );
  AND2_X1 U399 ( .A1(n385), .A2(n383), .ZN(n381) );
  XNOR2_X1 U400 ( .A(n361), .B(n615), .ZN(n360) );
  AND2_X1 U401 ( .A1(n462), .A2(n460), .ZN(n459) );
  NAND2_X1 U402 ( .A1(n776), .A2(n378), .ZN(n352) );
  OR2_X1 U403 ( .A1(n771), .A2(n612), .ZN(n609) );
  NAND2_X1 U404 ( .A1(n349), .A2(n781), .ZN(n440) );
  XNOR2_X1 U405 ( .A(n355), .B(n659), .ZN(n817) );
  NAND2_X1 U406 ( .A1(n356), .A2(n595), .ZN(n355) );
  AND2_X1 U407 ( .A1(n377), .A2(n589), .ZN(n376) );
  OR2_X2 U408 ( .A1(n371), .A2(n367), .ZN(n479) );
  NAND2_X1 U409 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U410 ( .A1(n393), .A2(n735), .ZN(n392) );
  AND2_X1 U411 ( .A1(n384), .A2(n735), .ZN(n383) );
  XNOR2_X1 U412 ( .A(n364), .B(G478), .ZN(n614) );
  OR2_X1 U413 ( .A1(n691), .A2(G210), .ZN(n384) );
  INV_X1 U414 ( .A(n691), .ZN(n382) );
  INV_X1 U415 ( .A(n732), .ZN(n390) );
  OR2_X1 U416 ( .A1(n732), .A2(G472), .ZN(n393) );
  NAND2_X1 U417 ( .A1(n738), .A2(n369), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n570), .ZN(n738) );
  XNOR2_X1 U419 ( .A(n723), .B(n547), .ZN(n690) );
  NOR2_X1 U420 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U421 ( .A1(n370), .A2(n369), .ZN(n368) );
  INV_X1 U422 ( .A(n374), .ZN(n370) );
  NAND2_X1 U423 ( .A1(n374), .A2(G902), .ZN(n372) );
  INV_X1 U424 ( .A(n563), .ZN(n375) );
  INV_X1 U425 ( .A(n441), .ZN(n374) );
  INV_X1 U426 ( .A(n658), .ZN(n357) );
  INV_X1 U427 ( .A(G110), .ZN(n398) );
  XNOR2_X1 U428 ( .A(G110), .B(G128), .ZN(n421) );
  XNOR2_X1 U429 ( .A(G140), .B(G137), .ZN(n510) );
  XNOR2_X1 U430 ( .A(G119), .B(KEYINPUT23), .ZN(n420) );
  INV_X1 U431 ( .A(G101), .ZN(n397) );
  NAND2_X1 U432 ( .A1(n347), .A2(n350), .ZN(n590) );
  NAND2_X1 U433 ( .A1(n351), .A2(n375), .ZN(n350) );
  INV_X1 U434 ( .A(n776), .ZN(n351) );
  XNOR2_X1 U435 ( .A(n529), .B(n353), .ZN(n354) );
  XNOR2_X2 U436 ( .A(n804), .B(G146), .ZN(n353) );
  XNOR2_X1 U437 ( .A(n354), .B(n731), .ZN(n732) );
  NAND2_X1 U438 ( .A1(n667), .A2(n480), .ZN(n358) );
  NAND2_X1 U439 ( .A1(n362), .A2(n360), .ZN(n359) );
  NAND2_X1 U440 ( .A1(n456), .A2(n729), .ZN(n361) );
  XNOR2_X1 U441 ( .A(n363), .B(KEYINPUT44), .ZN(n362) );
  XNOR2_X1 U442 ( .A(n571), .B(n573), .ZN(n365) );
  XNOR2_X2 U443 ( .A(n479), .B(KEYINPUT1), .ZN(n594) );
  NOR2_X1 U444 ( .A1(n697), .A2(n368), .ZN(n367) );
  NAND2_X1 U445 ( .A1(n697), .A2(n374), .ZN(n373) );
  AND2_X1 U446 ( .A1(n607), .A2(n563), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n693), .ZN(G51) );
  NAND2_X1 U448 ( .A1(n413), .A2(n386), .ZN(n385) );
  AND2_X1 U449 ( .A1(n691), .A2(G210), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U451 ( .A(n401), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n401), .A2(n395), .ZN(n394) );
  AND2_X1 U453 ( .A1(n732), .A2(G472), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n569), .B(n495), .ZN(n570) );
  BUF_X1 U455 ( .A(n423), .Z(n396) );
  NAND2_X1 U456 ( .A1(G101), .A2(n398), .ZN(n399) );
  NAND2_X1 U457 ( .A1(n397), .A2(G110), .ZN(n400) );
  NAND2_X1 U458 ( .A1(n399), .A2(n400), .ZN(n499) );
  XNOR2_X1 U459 ( .A(n687), .B(n443), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n687), .B(n443), .ZN(n413) );
  NAND2_X1 U461 ( .A1(n452), .A2(n465), .ZN(n456) );
  NOR2_X1 U462 ( .A1(n467), .A2(n466), .ZN(n465) );
  INV_X1 U463 ( .A(KEYINPUT78), .ZN(n477) );
  XNOR2_X1 U464 ( .A(n588), .B(n587), .ZN(n702) );
  INV_X1 U465 ( .A(KEYINPUT100), .ZN(n468) );
  XNOR2_X1 U466 ( .A(G104), .B(G107), .ZN(n501) );
  NOR2_X1 U467 ( .A1(n407), .A2(n418), .ZN(n417) );
  NOR2_X1 U468 ( .A1(n668), .A2(KEYINPUT19), .ZN(n418) );
  NAND2_X1 U469 ( .A1(n415), .A2(n556), .ZN(n414) );
  NOR2_X2 U470 ( .A1(G953), .A2(G237), .ZN(n578) );
  XNOR2_X1 U471 ( .A(KEYINPUT4), .B(G131), .ZN(n498) );
  XNOR2_X1 U472 ( .A(n471), .B(n470), .ZN(n666) );
  INV_X1 U473 ( .A(KEYINPUT39), .ZN(n470) );
  NOR2_X1 U474 ( .A1(n764), .A2(KEYINPUT79), .ZN(n461) );
  NOR2_X1 U475 ( .A1(n595), .A2(n603), .ZN(n463) );
  NOR2_X1 U476 ( .A1(n444), .A2(n438), .ZN(n437) );
  INV_X1 U477 ( .A(n744), .ZN(n464) );
  NOR2_X1 U478 ( .A1(n744), .A2(n409), .ZN(n467) );
  NOR2_X1 U479 ( .A1(n781), .A2(n468), .ZN(n466) );
  INV_X1 U480 ( .A(n680), .ZN(n490) );
  XNOR2_X1 U481 ( .A(G902), .B(KEYINPUT15), .ZN(n678) );
  XNOR2_X1 U482 ( .A(G131), .B(KEYINPUT93), .ZN(n576) );
  XNOR2_X1 U483 ( .A(G143), .B(G140), .ZN(n583) );
  XOR2_X1 U484 ( .A(KEYINPUT94), .B(G122), .Z(n584) );
  INV_X1 U485 ( .A(n800), .ZN(n493) );
  XNOR2_X1 U486 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n541) );
  XNOR2_X1 U487 ( .A(KEYINPUT83), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U488 ( .A1(G234), .A2(G237), .ZN(n557) );
  INV_X1 U489 ( .A(G237), .ZN(n548) );
  NAND2_X1 U490 ( .A1(n416), .A2(n414), .ZN(n562) );
  AND2_X1 U491 ( .A1(n419), .A2(n417), .ZN(n416) );
  XNOR2_X1 U492 ( .A(n421), .B(n420), .ZN(n507) );
  XNOR2_X1 U493 ( .A(G116), .B(KEYINPUT99), .ZN(n567) );
  NAND2_X1 U494 ( .A1(n436), .A2(n735), .ZN(n435) );
  NAND2_X1 U495 ( .A1(n698), .A2(n441), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n621), .B(n620), .ZN(n792) );
  INV_X1 U497 ( .A(n657), .ZN(n480) );
  NAND2_X1 U498 ( .A1(n473), .A2(n472), .ZN(n645) );
  XNOR2_X1 U499 ( .A(n634), .B(n410), .ZN(n472) );
  AND2_X1 U500 ( .A1(n636), .A2(n635), .ZN(n473) );
  XNOR2_X1 U501 ( .A(G113), .B(G137), .ZN(n526) );
  XNOR2_X1 U502 ( .A(n537), .B(n574), .ZN(n474) );
  XNOR2_X1 U503 ( .A(n538), .B(n539), .ZN(n475) );
  XNOR2_X1 U504 ( .A(n639), .B(n638), .ZN(n727) );
  NAND2_X1 U505 ( .A1(n476), .A2(n596), .ZN(n597) );
  NAND2_X1 U506 ( .A1(n459), .A2(n457), .ZN(n729) );
  NAND2_X1 U507 ( .A1(n458), .A2(n603), .ZN(n457) );
  NOR2_X1 U508 ( .A1(n461), .A2(n629), .ZN(n460) );
  XNOR2_X1 U509 ( .A(n439), .B(n703), .ZN(n704) );
  NAND2_X1 U510 ( .A1(n427), .A2(n403), .ZN(n425) );
  INV_X1 U511 ( .A(n437), .ZN(n427) );
  AND2_X1 U512 ( .A1(n676), .A2(KEYINPUT65), .ZN(n402) );
  AND2_X1 U513 ( .A1(n434), .A2(n426), .ZN(n403) );
  XOR2_X1 U514 ( .A(KEYINPUT13), .B(G475), .Z(n404) );
  AND2_X1 U515 ( .A1(n668), .A2(KEYINPUT19), .ZN(n405) );
  XOR2_X1 U516 ( .A(n657), .B(KEYINPUT19), .Z(n406) );
  AND2_X1 U517 ( .A1(n627), .A2(n560), .ZN(n407) );
  OR2_X1 U518 ( .A1(n468), .A2(n464), .ZN(n408) );
  NAND2_X1 U519 ( .A1(n781), .A2(n468), .ZN(n409) );
  XOR2_X1 U520 ( .A(KEYINPUT106), .B(KEYINPUT30), .Z(n410) );
  AND2_X1 U521 ( .A1(n680), .A2(n681), .ZN(n411) );
  AND2_X1 U522 ( .A1(n490), .A2(KEYINPUT65), .ZN(n412) );
  INV_X1 U523 ( .A(G469), .ZN(n441) );
  INV_X1 U524 ( .A(KEYINPUT64), .ZN(n443) );
  INV_X1 U525 ( .A(KEYINPUT65), .ZN(n681) );
  NAND2_X1 U526 ( .A1(n618), .A2(n668), .ZN(n657) );
  INV_X1 U527 ( .A(n618), .ZN(n415) );
  NAND2_X1 U528 ( .A1(n618), .A2(n405), .ZN(n419) );
  XNOR2_X2 U529 ( .A(n552), .B(n551), .ZN(n618) );
  OR2_X2 U530 ( .A1(n423), .A2(G902), .ZN(n517) );
  XNOR2_X1 U531 ( .A(n396), .B(n422), .ZN(n733) );
  INV_X1 U532 ( .A(KEYINPUT123), .ZN(n422) );
  XNOR2_X1 U533 ( .A(n513), .B(n512), .ZN(n423) );
  XNOR2_X2 U534 ( .A(n424), .B(G143), .ZN(n565) );
  XNOR2_X2 U535 ( .A(G128), .B(G134), .ZN(n424) );
  NAND2_X1 U536 ( .A1(n428), .A2(n425), .ZN(G54) );
  NOR2_X1 U537 ( .A1(n435), .A2(n699), .ZN(n426) );
  INV_X1 U538 ( .A(n429), .ZN(n428) );
  NAND2_X1 U539 ( .A1(n433), .A2(n430), .ZN(n429) );
  NAND2_X1 U540 ( .A1(n431), .A2(n699), .ZN(n430) );
  NAND2_X1 U541 ( .A1(n434), .A2(n432), .ZN(n431) );
  INV_X1 U542 ( .A(n435), .ZN(n432) );
  NAND2_X1 U543 ( .A1(n437), .A2(n699), .ZN(n433) );
  NAND2_X1 U544 ( .A1(n444), .A2(n698), .ZN(n434) );
  OR2_X1 U545 ( .A1(n698), .A2(n441), .ZN(n438) );
  NAND2_X1 U546 ( .A1(n448), .A2(G475), .ZN(n439) );
  XNOR2_X1 U547 ( .A(n442), .B(n443), .ZN(n448) );
  NAND2_X1 U548 ( .A1(n440), .A2(KEYINPUT47), .ZN(n649) );
  NOR2_X2 U549 ( .A1(n778), .A2(n777), .ZN(n494) );
  NAND2_X2 U550 ( .A1(n484), .A2(n483), .ZN(n687) );
  XNOR2_X2 U551 ( .A(n478), .B(n477), .ZN(n486) );
  NAND2_X2 U552 ( .A1(n598), .A2(n655), .ZN(n478) );
  NAND2_X2 U553 ( .A1(n594), .A2(n762), .ZN(n523) );
  XNOR2_X2 U554 ( .A(KEYINPUT74), .B(KEYINPUT88), .ZN(n504) );
  NAND2_X1 U555 ( .A1(n484), .A2(n483), .ZN(n442) );
  XNOR2_X1 U556 ( .A(n687), .B(KEYINPUT64), .ZN(n444) );
  BUF_X1 U557 ( .A(n469), .Z(n445) );
  BUF_X2 U558 ( .A(n684), .Z(n685) );
  XNOR2_X1 U559 ( .A(n590), .B(KEYINPUT35), .ZN(n469) );
  OR2_X2 U560 ( .A1(n614), .A2(n642), .ZN(n591) );
  XNOR2_X2 U561 ( .A(n597), .B(KEYINPUT32), .ZN(n716) );
  BUF_X1 U562 ( .A(n697), .Z(n446) );
  XNOR2_X1 U563 ( .A(n503), .B(n493), .ZN(n492) );
  XNOR2_X1 U564 ( .A(n508), .B(n801), .ZN(n513) );
  XNOR2_X2 U565 ( .A(n633), .B(n632), .ZN(n818) );
  OR2_X2 U566 ( .A1(n792), .A2(n641), .ZN(n633) );
  XNOR2_X2 U567 ( .A(n671), .B(KEYINPUT38), .ZN(n778) );
  XNOR2_X1 U568 ( .A(G143), .B(G128), .ZN(n447) );
  NAND2_X1 U569 ( .A1(n685), .A2(n616), .ZN(n449) );
  NAND2_X1 U570 ( .A1(n684), .A2(n616), .ZN(n617) );
  XNOR2_X1 U571 ( .A(n449), .B(KEYINPUT75), .ZN(n450) );
  BUF_X1 U572 ( .A(n804), .Z(n451) );
  XNOR2_X1 U573 ( .A(n617), .B(KEYINPUT75), .ZN(n677) );
  NOR2_X2 U574 ( .A1(n727), .A2(n818), .ZN(n640) );
  NAND2_X1 U575 ( .A1(n454), .A2(n453), .ZN(n452) );
  NAND2_X1 U576 ( .A1(n408), .A2(n713), .ZN(n453) );
  NAND2_X1 U577 ( .A1(n455), .A2(n409), .ZN(n454) );
  INV_X1 U578 ( .A(n713), .ZN(n455) );
  INV_X1 U579 ( .A(n486), .ZN(n458) );
  NAND2_X1 U580 ( .A1(n486), .A2(n463), .ZN(n462) );
  XNOR2_X1 U581 ( .A(n445), .B(n730), .ZN(G24) );
  OR2_X2 U582 ( .A1(n690), .A2(n616), .ZN(n552) );
  INV_X1 U583 ( .A(n478), .ZN(n476) );
  AND2_X1 U584 ( .A1(n479), .A2(n762), .ZN(n636) );
  NAND2_X1 U585 ( .A1(n497), .A2(n479), .ZN(n631) );
  AND2_X2 U586 ( .A1(n759), .A2(n758), .ZN(n762) );
  INV_X1 U587 ( .A(n642), .ZN(n613) );
  NAND2_X1 U588 ( .A1(n482), .A2(n642), .ZN(n652) );
  XNOR2_X2 U589 ( .A(n481), .B(n404), .ZN(n642) );
  INV_X1 U590 ( .A(n614), .ZN(n482) );
  NAND2_X1 U591 ( .A1(n402), .A2(n450), .ZN(n483) );
  AND2_X2 U592 ( .A1(n489), .A2(n485), .ZN(n484) );
  NAND2_X1 U593 ( .A1(n677), .A2(n676), .ZN(n491) );
  XNOR2_X2 U594 ( .A(n488), .B(n487), .ZN(n538) );
  XNOR2_X2 U595 ( .A(KEYINPUT3), .B(G119), .ZN(n487) );
  XNOR2_X2 U596 ( .A(G116), .B(G101), .ZN(n488) );
  NAND2_X1 U597 ( .A1(n491), .A2(n411), .ZN(n489) );
  XNOR2_X2 U598 ( .A(n517), .B(n516), .ZN(n629) );
  XNOR2_X1 U599 ( .A(n586), .B(n585), .ZN(n587) );
  BUF_X1 U600 ( .A(n776), .Z(n791) );
  XNOR2_X1 U601 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X2 U602 ( .A(n609), .B(n608), .ZN(n713) );
  XOR2_X1 U603 ( .A(n568), .B(n567), .Z(n495) );
  AND2_X1 U604 ( .A1(n779), .A2(n758), .ZN(n496) );
  XOR2_X1 U605 ( .A(n630), .B(KEYINPUT28), .Z(n497) );
  INV_X1 U606 ( .A(KEYINPUT71), .ZN(n675) );
  XNOR2_X1 U607 ( .A(n754), .B(n675), .ZN(n676) );
  BUF_X1 U608 ( .A(n754), .Z(n805) );
  INV_X1 U609 ( .A(KEYINPUT22), .ZN(n592) );
  INV_X1 U610 ( .A(KEYINPUT60), .ZN(n705) );
  XNOR2_X2 U611 ( .A(n565), .B(n498), .ZN(n804) );
  XNOR2_X1 U612 ( .A(n510), .B(KEYINPUT87), .ZN(n800) );
  NAND2_X1 U613 ( .A1(G227), .A2(n623), .ZN(n500) );
  XNOR2_X1 U614 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U615 ( .A(KEYINPUT24), .B(KEYINPUT72), .ZN(n505) );
  XNOR2_X1 U616 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U617 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U618 ( .A(G146), .B(G125), .ZN(n543) );
  XNOR2_X1 U619 ( .A(n543), .B(KEYINPUT10), .ZN(n801) );
  XNOR2_X1 U620 ( .A(n509), .B(KEYINPUT8), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n566), .A2(G221), .ZN(n511) );
  XNOR2_X1 U622 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U623 ( .A1(n678), .A2(G234), .ZN(n514) );
  XNOR2_X1 U624 ( .A(n514), .B(KEYINPUT20), .ZN(n518) );
  NAND2_X1 U625 ( .A1(n518), .A2(G217), .ZN(n515) );
  XNOR2_X1 U626 ( .A(n515), .B(KEYINPUT25), .ZN(n516) );
  INV_X1 U627 ( .A(n518), .ZN(n520) );
  INV_X1 U628 ( .A(G221), .ZN(n519) );
  OR2_X1 U629 ( .A1(n520), .A2(n519), .ZN(n522) );
  INV_X1 U630 ( .A(KEYINPUT21), .ZN(n521) );
  XNOR2_X1 U631 ( .A(n522), .B(n521), .ZN(n758) );
  XNOR2_X2 U632 ( .A(n523), .B(KEYINPUT70), .ZN(n604) );
  INV_X1 U633 ( .A(KEYINPUT104), .ZN(n524) );
  XNOR2_X1 U634 ( .A(n604), .B(n524), .ZN(n534) );
  NAND2_X1 U635 ( .A1(n578), .A2(G210), .ZN(n525) );
  XNOR2_X1 U636 ( .A(n525), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U637 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n538), .B(n528), .ZN(n529) );
  INV_X1 U639 ( .A(KEYINPUT89), .ZN(n530) );
  XNOR2_X1 U640 ( .A(n530), .B(G472), .ZN(n531) );
  XNOR2_X2 U641 ( .A(n532), .B(n531), .ZN(n769) );
  XNOR2_X1 U642 ( .A(n769), .B(KEYINPUT6), .ZN(n655) );
  INV_X1 U643 ( .A(n655), .ZN(n533) );
  NAND2_X1 U644 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U645 ( .A(KEYINPUT68), .B(KEYINPUT16), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n536), .B(G110), .ZN(n537) );
  XNOR2_X1 U647 ( .A(n710), .B(G104), .ZN(n574) );
  XNOR2_X1 U648 ( .A(n730), .B(G107), .ZN(n572) );
  INV_X1 U649 ( .A(n572), .ZN(n539) );
  NAND2_X1 U650 ( .A1(n623), .A2(G224), .ZN(n540) );
  XNOR2_X1 U651 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U652 ( .A(n543), .B(n542), .ZN(n546) );
  XNOR2_X1 U653 ( .A(n447), .B(n544), .ZN(n545) );
  XNOR2_X1 U654 ( .A(n546), .B(n545), .ZN(n547) );
  INV_X1 U655 ( .A(n678), .ZN(n616) );
  NAND2_X1 U656 ( .A1(n369), .A2(n548), .ZN(n553) );
  NAND2_X1 U657 ( .A1(n553), .A2(G210), .ZN(n550) );
  INV_X1 U658 ( .A(KEYINPUT84), .ZN(n549) );
  XNOR2_X1 U659 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U660 ( .A1(n553), .A2(G214), .ZN(n555) );
  INV_X1 U661 ( .A(KEYINPUT85), .ZN(n554) );
  XNOR2_X1 U662 ( .A(n555), .B(n554), .ZN(n668) );
  INV_X1 U663 ( .A(n668), .ZN(n777) );
  INV_X1 U664 ( .A(KEYINPUT19), .ZN(n556) );
  XOR2_X1 U665 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n558) );
  XNOR2_X1 U666 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U667 ( .A1(G952), .A2(n559), .ZN(n790) );
  OR2_X1 U668 ( .A1(n790), .A2(G953), .ZN(n627) );
  NAND2_X1 U669 ( .A1(G902), .A2(n559), .ZN(n622) );
  XOR2_X1 U670 ( .A(G898), .B(KEYINPUT86), .Z(n720) );
  NAND2_X1 U671 ( .A1(G953), .A2(n720), .ZN(n724) );
  OR2_X1 U672 ( .A1(n622), .A2(n724), .ZN(n560) );
  INV_X1 U673 ( .A(KEYINPUT0), .ZN(n561) );
  INV_X1 U674 ( .A(KEYINPUT34), .ZN(n563) );
  XNOR2_X1 U675 ( .A(KEYINPUT98), .B(KEYINPUT9), .ZN(n564) );
  XNOR2_X1 U676 ( .A(n565), .B(n564), .ZN(n571) );
  NAND2_X1 U677 ( .A1(G217), .A2(n566), .ZN(n569) );
  XOR2_X1 U678 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n568) );
  XNOR2_X1 U679 ( .A(n572), .B(KEYINPUT7), .ZN(n573) );
  BUF_X1 U680 ( .A(n614), .Z(n644) );
  XNOR2_X1 U681 ( .A(n574), .B(KEYINPUT91), .ZN(n575) );
  XNOR2_X1 U682 ( .A(n801), .B(n575), .ZN(n588) );
  XOR2_X1 U683 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n577) );
  XNOR2_X1 U684 ( .A(n577), .B(n576), .ZN(n582) );
  XOR2_X1 U685 ( .A(KEYINPUT92), .B(KEYINPUT95), .Z(n580) );
  NAND2_X1 U686 ( .A1(G214), .A2(n578), .ZN(n579) );
  XNOR2_X1 U687 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U688 ( .A(n582), .B(n581), .ZN(n586) );
  XNOR2_X1 U689 ( .A(n584), .B(n583), .ZN(n585) );
  AND2_X1 U690 ( .A1(n644), .A2(n642), .ZN(n589) );
  XNOR2_X2 U691 ( .A(n591), .B(KEYINPUT101), .ZN(n779) );
  NAND2_X1 U692 ( .A1(n496), .A2(n607), .ZN(n593) );
  XNOR2_X2 U693 ( .A(n593), .B(n592), .ZN(n598) );
  BUF_X1 U694 ( .A(n594), .Z(n595) );
  INV_X1 U695 ( .A(n595), .ZN(n764) );
  AND2_X1 U696 ( .A1(n595), .A2(n629), .ZN(n596) );
  NAND2_X1 U697 ( .A1(n598), .A2(n764), .ZN(n599) );
  XNOR2_X1 U698 ( .A(n599), .B(KEYINPUT103), .ZN(n601) );
  INV_X1 U699 ( .A(n769), .ZN(n610) );
  AND2_X1 U700 ( .A1(n610), .A2(n629), .ZN(n600) );
  NAND2_X1 U701 ( .A1(n601), .A2(n600), .ZN(n715) );
  NAND2_X1 U702 ( .A1(n716), .A2(n715), .ZN(n602) );
  INV_X1 U703 ( .A(KEYINPUT79), .ZN(n603) );
  NOR2_X1 U704 ( .A1(n604), .A2(n610), .ZN(n606) );
  INV_X1 U705 ( .A(KEYINPUT90), .ZN(n605) );
  XNOR2_X1 U706 ( .A(n606), .B(n605), .ZN(n771) );
  INV_X1 U707 ( .A(n607), .ZN(n612) );
  INV_X1 U708 ( .A(KEYINPUT31), .ZN(n608) );
  NAND2_X1 U709 ( .A1(n636), .A2(n610), .ZN(n611) );
  OR2_X1 U710 ( .A1(n612), .A2(n611), .ZN(n744) );
  NAND2_X1 U711 ( .A1(n644), .A2(n613), .ZN(n743) );
  NAND2_X1 U712 ( .A1(n743), .A2(n652), .ZN(n781) );
  INV_X1 U713 ( .A(KEYINPUT102), .ZN(n615) );
  NAND2_X1 U714 ( .A1(n779), .A2(n494), .ZN(n621) );
  XNOR2_X1 U715 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n619) );
  XNOR2_X1 U716 ( .A(n619), .B(KEYINPUT41), .ZN(n620) );
  INV_X1 U717 ( .A(G900), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U719 ( .A1(n627), .A2(n626), .ZN(n635) );
  AND2_X1 U720 ( .A1(n758), .A2(n635), .ZN(n628) );
  AND2_X1 U721 ( .A1(n629), .A2(n628), .ZN(n653) );
  NAND2_X1 U722 ( .A1(n769), .A2(n653), .ZN(n630) );
  XNOR2_X1 U723 ( .A(n631), .B(KEYINPUT108), .ZN(n641) );
  INV_X1 U724 ( .A(KEYINPUT42), .ZN(n632) );
  NAND2_X1 U725 ( .A1(n769), .A2(n668), .ZN(n634) );
  INV_X1 U726 ( .A(n652), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n666), .A2(n637), .ZN(n639) );
  INV_X1 U728 ( .A(KEYINPUT40), .ZN(n638) );
  XNOR2_X1 U729 ( .A(n640), .B(KEYINPUT46), .ZN(n663) );
  OR2_X2 U730 ( .A1(n641), .A2(n406), .ZN(n751) );
  AND2_X1 U731 ( .A1(n671), .A2(n642), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n644), .A2(n643), .ZN(n646) );
  OR2_X1 U733 ( .A1(n646), .A2(n645), .ZN(n648) );
  INV_X1 U734 ( .A(KEYINPUT107), .ZN(n647) );
  XNOR2_X1 U735 ( .A(n648), .B(n647), .ZN(n815) );
  NAND2_X1 U736 ( .A1(n649), .A2(n815), .ZN(n650) );
  XNOR2_X1 U737 ( .A(n650), .B(KEYINPUT73), .ZN(n661) );
  INV_X1 U738 ( .A(KEYINPUT105), .ZN(n651) );
  XNOR2_X1 U739 ( .A(n652), .B(n651), .ZN(n708) );
  INV_X1 U740 ( .A(n653), .ZN(n654) );
  OR2_X1 U741 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U742 ( .A(KEYINPUT80), .B(KEYINPUT36), .ZN(n658) );
  INV_X1 U743 ( .A(KEYINPUT111), .ZN(n659) );
  AND2_X1 U744 ( .A1(n348), .A2(n817), .ZN(n660) );
  AND2_X1 U745 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U746 ( .A1(n663), .A2(n662), .ZN(n665) );
  XNOR2_X1 U747 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n665), .B(n664), .ZN(n674) );
  INV_X1 U749 ( .A(n743), .ZN(n748) );
  NAND2_X1 U750 ( .A1(n666), .A2(n748), .ZN(n707) );
  NAND2_X1 U751 ( .A1(n668), .A2(n667), .ZN(n669) );
  OR2_X1 U752 ( .A1(n595), .A2(n669), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(KEYINPUT43), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(n415), .ZN(n712) );
  AND2_X1 U755 ( .A1(n707), .A2(n712), .ZN(n673) );
  NAND2_X2 U756 ( .A1(n674), .A2(n673), .ZN(n683) );
  XNOR2_X2 U757 ( .A(n683), .B(KEYINPUT77), .ZN(n754) );
  XOR2_X1 U758 ( .A(KEYINPUT76), .B(n678), .Z(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(KEYINPUT2), .ZN(n680) );
  INV_X1 U760 ( .A(KEYINPUT2), .ZN(n682) );
  NOR2_X1 U761 ( .A1(n683), .A2(n682), .ZN(n686) );
  XNOR2_X1 U762 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n688) );
  XOR2_X1 U763 ( .A(n688), .B(KEYINPUT55), .Z(n689) );
  XNOR2_X1 U764 ( .A(n690), .B(n689), .ZN(n691) );
  INV_X1 U765 ( .A(G952), .ZN(n692) );
  NAND2_X1 U766 ( .A1(n692), .A2(G953), .ZN(n735) );
  INV_X1 U767 ( .A(KEYINPUT56), .ZN(n693) );
  XOR2_X1 U768 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n695) );
  XNOR2_X1 U769 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n694) );
  XOR2_X1 U770 ( .A(n695), .B(n694), .Z(n696) );
  XNOR2_X1 U771 ( .A(n446), .B(n696), .ZN(n698) );
  INV_X1 U772 ( .A(KEYINPUT120), .ZN(n699) );
  XNOR2_X1 U773 ( .A(KEYINPUT66), .B(KEYINPUT121), .ZN(n700) );
  XOR2_X1 U774 ( .A(n700), .B(KEYINPUT59), .Z(n701) );
  XNOR2_X1 U775 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U776 ( .A1(n704), .A2(n735), .ZN(n706) );
  XNOR2_X1 U777 ( .A(n706), .B(n705), .ZN(G60) );
  XNOR2_X1 U778 ( .A(n707), .B(G134), .ZN(G36) );
  BUF_X1 U779 ( .A(n708), .Z(n752) );
  NOR2_X1 U780 ( .A1(n752), .A2(n744), .ZN(n709) );
  XOR2_X1 U781 ( .A(G104), .B(n709), .Z(G6) );
  NOR2_X1 U782 ( .A1(n713), .A2(n752), .ZN(n711) );
  XNOR2_X1 U783 ( .A(n711), .B(n710), .ZN(G15) );
  XNOR2_X1 U784 ( .A(n712), .B(G140), .ZN(G42) );
  NOR2_X1 U785 ( .A1(n713), .A2(n743), .ZN(n714) );
  XOR2_X1 U786 ( .A(G116), .B(n714), .Z(G18) );
  XNOR2_X1 U787 ( .A(n715), .B(G110), .ZN(G12) );
  XNOR2_X1 U788 ( .A(n716), .B(G119), .ZN(G21) );
  INV_X1 U789 ( .A(n685), .ZN(n717) );
  NOR2_X1 U790 ( .A1(n717), .A2(G953), .ZN(n722) );
  NAND2_X1 U791 ( .A1(G953), .A2(G224), .ZN(n718) );
  XOR2_X1 U792 ( .A(KEYINPUT61), .B(n718), .Z(n719) );
  NOR2_X1 U793 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U795 ( .A1(n723), .A2(n724), .ZN(n725) );
  XNOR2_X1 U796 ( .A(n726), .B(n725), .ZN(G69) );
  XOR2_X1 U797 ( .A(G131), .B(n727), .Z(G33) );
  XNOR2_X1 U798 ( .A(G101), .B(KEYINPUT112), .ZN(n728) );
  XNOR2_X1 U799 ( .A(n729), .B(n728), .ZN(G3) );
  XOR2_X1 U800 ( .A(KEYINPUT82), .B(KEYINPUT62), .Z(n731) );
  BUF_X1 U801 ( .A(n448), .Z(n737) );
  NAND2_X1 U802 ( .A1(n737), .A2(G217), .ZN(n734) );
  XNOR2_X1 U803 ( .A(n734), .B(n733), .ZN(n736) );
  INV_X1 U804 ( .A(n735), .ZN(n741) );
  NOR2_X1 U805 ( .A1(n736), .A2(n741), .ZN(G66) );
  NAND2_X1 U806 ( .A1(n737), .A2(G478), .ZN(n740) );
  XOR2_X1 U807 ( .A(KEYINPUT122), .B(n738), .Z(n739) );
  XNOR2_X1 U808 ( .A(n740), .B(n739), .ZN(n742) );
  NOR2_X1 U809 ( .A1(n742), .A2(n741), .ZN(G63) );
  XOR2_X1 U810 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n746) );
  NOR2_X1 U811 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U812 ( .A(n746), .B(n745), .Z(n747) );
  XNOR2_X1 U813 ( .A(G107), .B(n747), .ZN(G9) );
  XOR2_X1 U814 ( .A(G128), .B(KEYINPUT29), .Z(n750) );
  NAND2_X1 U815 ( .A1(n349), .A2(n748), .ZN(n749) );
  XNOR2_X1 U816 ( .A(n750), .B(n749), .ZN(G30) );
  OR2_X1 U817 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U818 ( .A(n753), .B(G146), .ZN(G48) );
  AND2_X1 U819 ( .A1(n805), .A2(n685), .ZN(n755) );
  NOR2_X1 U820 ( .A1(n755), .A2(KEYINPUT2), .ZN(n757) );
  NOR2_X1 U821 ( .A1(n757), .A2(n756), .ZN(n796) );
  NOR2_X1 U822 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U823 ( .A(KEYINPUT113), .B(n760), .Z(n761) );
  XNOR2_X1 U824 ( .A(KEYINPUT49), .B(n761), .ZN(n768) );
  INV_X1 U825 ( .A(n762), .ZN(n763) );
  NAND2_X1 U826 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U827 ( .A(n765), .B(KEYINPUT114), .ZN(n766) );
  XNOR2_X1 U828 ( .A(KEYINPUT50), .B(n766), .ZN(n767) );
  NAND2_X1 U829 ( .A1(n768), .A2(n767), .ZN(n770) );
  OR2_X1 U830 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U831 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U832 ( .A(n773), .B(KEYINPUT115), .Z(n774) );
  XNOR2_X1 U833 ( .A(KEYINPUT51), .B(n774), .ZN(n775) );
  NOR2_X1 U834 ( .A1(n792), .A2(n775), .ZN(n787) );
  NAND2_X1 U835 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U836 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U837 ( .A1(n494), .A2(n781), .ZN(n782) );
  NAND2_X1 U838 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U839 ( .A1(n791), .A2(n784), .ZN(n785) );
  XOR2_X1 U840 ( .A(KEYINPUT116), .B(n785), .Z(n786) );
  NOR2_X1 U841 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U842 ( .A(n788), .B(KEYINPUT52), .ZN(n789) );
  NOR2_X1 U843 ( .A1(n790), .A2(n789), .ZN(n794) );
  NOR2_X1 U844 ( .A1(n792), .A2(n351), .ZN(n793) );
  OR2_X1 U845 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U846 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U847 ( .A(n797), .B(KEYINPUT117), .ZN(n798) );
  NOR2_X1 U848 ( .A1(G953), .A2(n798), .ZN(n799) );
  XNOR2_X1 U849 ( .A(KEYINPUT53), .B(n799), .ZN(G75) );
  XNOR2_X1 U850 ( .A(n800), .B(KEYINPUT124), .ZN(n802) );
  XNOR2_X1 U851 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U852 ( .A(n451), .B(n803), .ZN(n808) );
  XNOR2_X1 U853 ( .A(n805), .B(n808), .ZN(n806) );
  NOR2_X1 U854 ( .A1(n806), .A2(G953), .ZN(n807) );
  XNOR2_X1 U855 ( .A(KEYINPUT125), .B(n807), .ZN(n813) );
  XNOR2_X1 U856 ( .A(n808), .B(G227), .ZN(n809) );
  XNOR2_X1 U857 ( .A(n809), .B(KEYINPUT126), .ZN(n810) );
  NAND2_X1 U858 ( .A1(n810), .A2(G900), .ZN(n811) );
  NAND2_X1 U859 ( .A1(n811), .A2(G953), .ZN(n812) );
  NAND2_X1 U860 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U861 ( .A(KEYINPUT127), .B(n814), .Z(G72) );
  XNOR2_X1 U862 ( .A(G143), .B(n815), .ZN(G45) );
  XOR2_X1 U863 ( .A(G125), .B(KEYINPUT37), .Z(n816) );
  XNOR2_X1 U864 ( .A(n817), .B(n816), .ZN(G27) );
  XOR2_X1 U865 ( .A(G137), .B(n818), .Z(G39) );
endmodule

