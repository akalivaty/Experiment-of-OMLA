//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT27), .ZN(new_n214));
  AOI21_X1  g013(.A(G190gat), .B1(new_n214), .B2(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT28), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT68), .B1(new_n215), .B2(new_n220), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n223), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n217), .A3(new_n221), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n213), .A2(new_n224), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n231), .A2(new_n233), .A3(new_n205), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n227), .A2(KEYINPUT24), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n227), .A2(KEYINPUT24), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n231), .A2(new_n233), .A3(new_n205), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n244), .B2(KEYINPUT65), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n245), .A2(new_n234), .A3(new_n235), .A4(new_n239), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n243), .B2(new_n246), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n228), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G113gat), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  INV_X1    g056(.A(new_n251), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT71), .B(G113gat), .Z(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(G120gat), .B2(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n253), .A2(new_n257), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n250), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n253), .A2(new_n257), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n260), .A2(new_n256), .ZN(new_n264));
  OAI221_X1 g063(.A(new_n228), .B1(new_n263), .B2(new_n264), .C1(new_n248), .C2(new_n249), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n204), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n265), .A3(new_n204), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT34), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT32), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n267), .B2(KEYINPUT32), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(KEYINPUT32), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT34), .ZN(new_n274));
  INV_X1    g073(.A(new_n266), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n269), .ZN(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G71gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(G99gat), .Z(new_n279));
  INV_X1    g078(.A(new_n267), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT33), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n272), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n272), .B2(new_n276), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n202), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n288), .B(new_n202), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n276), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n281), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT36), .A3(new_n283), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n292), .A2(new_n295), .A3(KEYINPUT36), .A4(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(KEYINPUT76), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n250), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n228), .A2(new_n246), .A3(new_n243), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n299), .ZN(new_n306));
  XOR2_X1   g105(.A(G197gat), .B(G204gat), .Z(new_n307));
  AOI21_X1  g106(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G211gat), .B(G218gat), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n309), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n250), .A2(new_n304), .ZN(new_n315));
  INV_X1    g114(.A(new_n299), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n315), .A2(new_n300), .B1(new_n316), .B2(new_n303), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n313), .B(KEYINPUT75), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n314), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT78), .ZN(new_n322));
  INV_X1    g121(.A(G64gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G92gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT30), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n300), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n303), .A2(new_n316), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n319), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n314), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT77), .B(new_n314), .C1(new_n317), .C2(new_n319), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n330), .B1(new_n338), .B2(new_n327), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n329), .B1(new_n339), .B2(new_n328), .ZN(new_n340));
  INV_X1    g139(.A(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G141gat), .ZN(new_n342));
  INV_X1    g141(.A(G141gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n345), .A2(new_n346), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT79), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(KEYINPUT80), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(new_n344), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n346), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n351), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT81), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n347), .A2(new_n349), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n351), .A2(new_n353), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n355), .A2(new_n354), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n261), .B1(new_n363), .B2(KEYINPUT3), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n350), .A2(new_n356), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n261), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n261), .A2(new_n365), .A3(KEYINPUT82), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n261), .A2(new_n365), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n368), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  INV_X1    g178(.A(new_n363), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n374), .B1(new_n380), .B2(new_n261), .ZN(new_n381));
  INV_X1    g180(.A(new_n377), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n364), .A2(new_n367), .B1(new_n370), .B2(new_n375), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n382), .A2(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n370), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n368), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(KEYINPUT86), .A3(new_n382), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n385), .B2(new_n377), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT39), .B1(new_n381), .B2(new_n382), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT39), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n393), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT40), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n403), .A2(KEYINPUT40), .A3(new_n393), .A4(new_n405), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n340), .A2(new_n395), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G228gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n367), .A2(new_n304), .ZN(new_n414));
  INV_X1    g213(.A(new_n313), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n309), .ZN(new_n417));
  INV_X1    g216(.A(new_n310), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n309), .A2(new_n310), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT3), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n416), .B1(new_n421), .B2(new_n365), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n366), .B1(new_n415), .B2(KEYINPUT29), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n318), .A2(new_n414), .B1(new_n363), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n413), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G78gat), .B(G106gat), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G22gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n427), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n428), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n320), .A2(KEYINPUT37), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n327), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(KEYINPUT37), .B2(new_n338), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n328), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND4_X1   g239(.A1(KEYINPUT84), .A2(new_n384), .A3(new_n393), .A4(new_n387), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n378), .A2(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT84), .B1(new_n442), .B2(new_n393), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n395), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n395), .A2(new_n446), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n384), .A2(new_n393), .A3(new_n387), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n442), .A2(KEYINPUT84), .A3(new_n393), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n395), .A3(new_n453), .A4(new_n446), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT87), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n317), .A2(new_n319), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n313), .B1(new_n302), .B2(new_n306), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT37), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n436), .A2(new_n458), .A3(new_n439), .A4(new_n327), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n447), .A2(new_n449), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n410), .B(new_n435), .C1(new_n440), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n395), .B(KEYINPUT85), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n452), .A2(new_n446), .A3(new_n453), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n448), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n434), .B1(new_n465), .B2(new_n340), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n298), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n434), .A2(new_n284), .A3(new_n285), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n449), .A3(new_n455), .ZN(new_n469));
  INV_X1    g268(.A(new_n340), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n284), .A2(new_n285), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n435), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n474), .A2(new_n465), .A3(new_n340), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n472), .B1(new_n475), .B2(new_n471), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT88), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n467), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G197gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT11), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(new_n229), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(G1gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(G1gat), .B2(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G8gat), .ZN(new_n492));
  INV_X1    g291(.A(G8gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n490), .B(new_n493), .C1(G1gat), .C2(new_n487), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT93), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT93), .B1(new_n492), .B2(new_n494), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500));
  INV_X1    g299(.A(G43gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(G50gat), .ZN(new_n502));
  INV_X1    g301(.A(G50gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(G43gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(G43gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(G50gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT15), .ZN(new_n508));
  NOR2_X1   g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT14), .ZN(new_n510));
  INV_X1    g309(.A(new_n509), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT14), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n505), .A2(new_n508), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT15), .ZN(new_n516));
  INV_X1    g315(.A(new_n510), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(KEYINPUT14), .B2(new_n512), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT90), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n499), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT93), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n495), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n521), .B(new_n523), .C1(new_n527), .C2(new_n498), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT92), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT13), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n521), .B2(new_n523), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n522), .B1(new_n515), .B2(new_n519), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT15), .B1(new_n506), .B2(new_n507), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n516), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n518), .A2(new_n517), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT90), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n537), .A2(new_n541), .A3(KEYINPUT17), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n496), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n544));
  INV_X1    g343(.A(new_n531), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n521), .A2(new_n535), .A3(new_n523), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT17), .B1(new_n537), .B2(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n496), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n544), .A2(new_n525), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n534), .B1(new_n552), .B2(KEYINPUT18), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n486), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n549), .B1(new_n548), .B2(new_n496), .ZN(new_n556));
  AOI211_X1 g355(.A(KEYINPUT91), .B(new_n495), .C1(new_n546), .C2(new_n547), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n525), .A4(new_n545), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n553), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n555), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n563), .B(new_n553), .C1(new_n554), .C2(new_n486), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n478), .A2(new_n480), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT21), .ZN(new_n569));
  INV_X1    g368(.A(G57gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(G64gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n323), .A2(G57gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT9), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  OR2_X1    g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT96), .B1(new_n323), .B2(G57gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n570), .A3(G64gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n578), .B1(new_n582), .B2(new_n571), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  OAI22_X1  g383(.A1(new_n527), .A2(new_n498), .B1(new_n569), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n569), .ZN(new_n586));
  INV_X1    g385(.A(G127gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT97), .B(G155gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n593), .B1(new_n589), .B2(new_n594), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n596), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G162gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT8), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(G99gat), .B2(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(G85gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT99), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(G85gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n611), .B1(new_n616), .B2(new_n325), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT98), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(G85gat), .A3(G92gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n619), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n621), .A2(new_n623), .A3(new_n619), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n617), .B(new_n618), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n622), .B1(G85gat), .B2(G92gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n620), .A2(KEYINPUT98), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT7), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n623), .A3(new_n619), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n618), .B1(new_n632), .B2(new_n617), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n609), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n617), .B1(new_n624), .B2(new_n625), .ZN(new_n635));
  INV_X1    g434(.A(new_n618), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(KEYINPUT100), .A3(new_n626), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n548), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n524), .A3(new_n638), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(G134gat), .ZN(new_n644));
  INV_X1    g443(.A(G134gat), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n640), .A2(new_n645), .A3(new_n641), .A4(new_n642), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n644), .B2(new_n646), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n608), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n547), .A2(new_n546), .B1(new_n634), .B2(new_n638), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n634), .A2(new_n524), .A3(new_n638), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n645), .B1(new_n654), .B2(new_n641), .ZN(new_n655));
  INV_X1    g454(.A(new_n646), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n607), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n605), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n230), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G204gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT103), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n618), .A2(KEYINPUT101), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n576), .A2(new_n583), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n627), .B2(new_n633), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n637), .A3(new_n626), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n584), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n634), .A2(new_n638), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n669), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n667), .B1(new_n672), .B2(new_n674), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n666), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n667), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n672), .A2(new_n674), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(G230gat), .A3(G233gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n665), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n681), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n662), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n568), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT85), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n395), .B(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n449), .B1(new_n693), .B2(new_n463), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(new_n488), .ZN(G1324gat));
  NOR2_X1   g499(.A1(new_n691), .A2(new_n470), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT16), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n702), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(G8gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(G8gat), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n706), .B(new_n707), .C1(KEYINPUT42), .C2(new_n701), .ZN(G1325gat));
  INV_X1    g507(.A(new_n691), .ZN(new_n709));
  INV_X1    g508(.A(new_n298), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n709), .A2(G15gat), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(G15gat), .B1(new_n709), .B2(new_n473), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n691), .A2(new_n435), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NAND4_X1  g515(.A1(new_n478), .A2(KEYINPUT44), .A3(new_n660), .A4(new_n480), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n649), .A2(new_n650), .A3(new_n608), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n607), .B1(new_n657), .B2(new_n658), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n467), .B2(new_n476), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n722));
  INV_X1    g521(.A(new_n567), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(new_n604), .A3(new_n689), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n717), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n698), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n478), .A2(new_n660), .A3(new_n480), .A4(new_n724), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(G29gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n729), .B2(new_n697), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n728), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n698), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n726), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT106), .Z(G1328gat));
  NOR3_X1   g532(.A1(new_n728), .A2(G36gat), .A3(new_n470), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G36gat), .B1(new_n725), .B2(new_n470), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(G1329gat));
  NAND2_X1  g538(.A1(new_n473), .A2(new_n501), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n717), .A2(new_n722), .A3(new_n710), .A4(new_n724), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n744), .A2(KEYINPUT107), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT107), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n744), .A2(KEYINPUT108), .A3(new_n745), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n743), .B2(KEYINPUT47), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n750), .ZN(G1330gat));
  OAI21_X1  g550(.A(G50gat), .B1(new_n725), .B2(new_n435), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n434), .A2(new_n503), .ZN(new_n753));
  OAI221_X1 g552(.A(new_n752), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n728), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1331gat));
  AOI21_X1  g555(.A(new_n567), .B1(new_n467), .B2(new_n476), .ZN(new_n757));
  INV_X1    g556(.A(new_n689), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n662), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n697), .B(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G57gat), .ZN(G1332gat));
  INV_X1    g562(.A(new_n760), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n470), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n760), .A2(G71gat), .A3(new_n710), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT111), .Z(new_n771));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n473), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n434), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n567), .A2(new_n604), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n721), .A2(KEYINPUT51), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n721), .B2(new_n779), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n781), .A2(KEYINPUT113), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(KEYINPUT113), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n697), .A2(new_n616), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n689), .A4(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n567), .A2(new_n604), .A3(new_n758), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n717), .A2(new_n722), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT112), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n717), .A2(new_n722), .A3(new_n790), .A4(new_n787), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n698), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n792), .B2(new_n616), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n786), .B(new_n795), .C1(new_n792), .C2(new_n616), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1336gat));
  AND2_X1   g596(.A1(new_n783), .A2(new_n784), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n470), .A2(G92gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n689), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n788), .B2(new_n470), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n789), .A2(new_n791), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n325), .B1(new_n804), .B2(new_n340), .ZN(new_n805));
  INV_X1    g604(.A(new_n782), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n780), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n689), .A3(new_n799), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n807), .A2(new_n810), .A3(new_n689), .A4(new_n799), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n803), .A2(new_n813), .ZN(G1337gat));
  NAND2_X1  g613(.A1(new_n804), .A2(new_n710), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n804), .A2(KEYINPUT116), .A3(new_n710), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(G99gat), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n773), .A2(G99gat), .A3(new_n758), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(G1338gat));
  NOR2_X1   g622(.A1(new_n435), .A2(G106gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n689), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g625(.A(G106gat), .B1(new_n788), .B2(new_n435), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(G106gat), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n829), .B1(new_n804), .B2(new_n434), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n807), .A2(new_n689), .A3(new_n824), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT53), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n828), .A2(new_n832), .ZN(G1339gat));
  OAI211_X1 g632(.A(new_n683), .B(KEYINPUT54), .C1(new_n682), .C2(new_n668), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI211_X1 g634(.A(KEYINPUT118), .B(new_n665), .C1(new_n679), .C2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n682), .A2(new_n835), .A3(new_n668), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n666), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n686), .B(KEYINPUT102), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT55), .B(new_n834), .C1(new_n836), .C2(new_n839), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n563), .A2(new_n553), .A3(new_n486), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n545), .B1(new_n558), .B2(new_n525), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n529), .A2(new_n532), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n484), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n660), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n845), .B1(new_n566), .B2(new_n565), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n846), .A2(new_n689), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n720), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n605), .B(new_n851), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n723), .A2(new_n661), .A3(new_n758), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n855), .A2(KEYINPUT119), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT119), .B1(new_n855), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n474), .A2(new_n340), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n697), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n723), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n761), .A2(new_n859), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n860), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n723), .A2(new_n259), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  OAI21_X1  g666(.A(G120gat), .B1(new_n861), .B2(new_n758), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n689), .A2(new_n255), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n865), .B2(new_n869), .ZN(G1341gat));
  NOR3_X1   g669(.A1(new_n861), .A2(new_n587), .A3(new_n605), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n864), .A2(new_n604), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n587), .ZN(G1342gat));
  NOR3_X1   g672(.A1(new_n865), .A2(G134gat), .A3(new_n720), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT120), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n861), .B2(new_n720), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n710), .A2(new_n435), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n761), .A2(new_n859), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT123), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(KEYINPUT123), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n470), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n723), .A2(G141gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n845), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n854), .B1(new_n567), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n851), .A2(new_n605), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n856), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n855), .A2(KEYINPUT119), .A3(new_n856), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n434), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(KEYINPUT121), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT121), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n892), .A2(new_n434), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n697), .A2(new_n298), .A3(new_n470), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n902), .A2(new_n723), .A3(new_n903), .ZN(new_n904));
  OAI221_X1 g703(.A(new_n881), .B1(new_n886), .B2(new_n888), .C1(new_n343), .C2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n883), .A2(new_n340), .A3(new_n888), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n857), .A2(new_n858), .A3(new_n435), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  INV_X1    g710(.A(new_n901), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n896), .A2(KEYINPUT121), .A3(new_n897), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n903), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(KEYINPUT122), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n908), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n567), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n906), .B1(new_n918), .B2(G141gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n905), .B1(new_n919), .B2(new_n881), .ZN(G1344gat));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n897), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n896), .B2(new_n897), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n689), .A3(new_n915), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n914), .A2(KEYINPUT122), .A3(new_n915), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT122), .B1(new_n914), .B2(new_n915), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n689), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n341), .A2(KEYINPUT59), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n886), .A2(G148gat), .A3(new_n758), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  INV_X1    g732(.A(new_n931), .ZN(new_n934));
  INV_X1    g733(.A(new_n929), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n935), .B1(new_n917), .B2(new_n689), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n933), .B(new_n934), .C1(new_n936), .C2(new_n925), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n937), .ZN(G1345gat));
  NOR2_X1   g737(.A1(new_n605), .A2(G155gat), .ZN(new_n939));
  AND4_X1   g738(.A1(new_n470), .A2(new_n884), .A3(new_n885), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n604), .B1(new_n926), .B2(new_n927), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(G155gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI211_X1 g743(.A(KEYINPUT125), .B(new_n940), .C1(new_n941), .C2(G155gat), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1346gat));
  NOR2_X1   g745(.A1(new_n886), .A2(new_n720), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n917), .A2(new_n660), .ZN(new_n948));
  MUX2_X1   g747(.A(new_n947), .B(new_n948), .S(G162gat), .Z(G1347gat));
  INV_X1    g748(.A(new_n761), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n474), .A2(new_n470), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n859), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n723), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT126), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n857), .A2(new_n858), .A3(new_n697), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n951), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n229), .A3(new_n567), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n954), .A2(new_n958), .ZN(G1348gat));
  NOR3_X1   g758(.A1(new_n952), .A2(new_n230), .A3(new_n758), .ZN(new_n960));
  AOI21_X1  g759(.A(G176gat), .B1(new_n957), .B2(new_n689), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1349gat));
  OAI21_X1  g761(.A(G183gat), .B1(new_n952), .B2(new_n605), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n957), .B(new_n604), .C1(KEYINPUT27), .C2(new_n219), .ZN(new_n964));
  INV_X1    g763(.A(new_n220), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g766(.A(G190gat), .B1(new_n952), .B2(new_n720), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT61), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n957), .A2(new_n237), .A3(new_n660), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1351gat));
  AND3_X1   g770(.A1(new_n955), .A2(new_n340), .A3(new_n882), .ZN(new_n972));
  INV_X1    g771(.A(G197gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n973), .A3(new_n567), .ZN(new_n974));
  AND4_X1   g773(.A1(new_n340), .A2(new_n923), .A3(new_n950), .A4(new_n298), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n975), .A2(new_n567), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n976), .B2(new_n973), .ZN(G1352gat));
  INV_X1    g776(.A(G204gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n972), .A2(new_n978), .A3(new_n689), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n950), .A2(new_n340), .A3(new_n298), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n923), .A2(new_n689), .ZN(new_n982));
  OAI21_X1  g781(.A(G204gat), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n980), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT127), .ZN(G1353gat));
  INV_X1    g785(.A(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n987), .B1(new_n975), .B2(new_n604), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT63), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n987), .A3(new_n604), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n972), .B2(new_n660), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n660), .A2(G218gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n975), .B2(new_n993), .ZN(G1355gat));
endmodule


