//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  OAI22_X1  g009(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT71), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n214), .A2(KEYINPUT70), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(KEYINPUT70), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n207), .B(new_n205), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n208), .A2(new_n209), .ZN(new_n218));
  INV_X1    g017(.A(G120gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G113gat), .ZN(new_n220));
  INV_X1    g019(.A(G113gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G120gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n217), .A2(new_n218), .A3(new_n225), .A4(KEYINPUT72), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n213), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n207), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n206), .A2(G127gat), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT79), .ZN(new_n236));
  XNOR2_X1  g035(.A(G155gat), .B(G162gat), .ZN(new_n237));
  OR3_X1    g036(.A1(new_n234), .A2(KEYINPUT79), .A3(G141gat), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT80), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G162gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G155gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT2), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n233), .A2(new_n235), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n237), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n239), .A2(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND4_X1   g050(.A1(new_n202), .A2(new_n227), .A3(new_n231), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n227), .A2(new_n231), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n250), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n248), .B1(new_n244), .B2(G155gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n238), .A3(new_n237), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n257), .B2(new_n256), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n230), .B1(new_n213), .B2(new_n226), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n202), .B1(new_n262), .B2(new_n251), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n252), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n264), .A2(KEYINPUT5), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT1), .B1(new_n220), .B2(new_n222), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n205), .A2(new_n207), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT72), .B1(new_n273), .B2(new_n218), .ZN(new_n274));
  AND4_X1   g073(.A1(KEYINPUT72), .A2(new_n217), .A3(new_n218), .A4(new_n225), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n231), .B(new_n251), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n258), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(KEYINPUT4), .C1(new_n277), .C2(new_n262), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n202), .A3(new_n251), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n269), .B1(new_n280), .B2(new_n265), .ZN(new_n281));
  AOI211_X1 g080(.A(KEYINPUT81), .B(new_n266), .C1(new_n278), .C2(new_n279), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT82), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n253), .A2(new_n259), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n265), .B1(new_n285), .B2(new_n276), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n276), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n262), .A2(new_n251), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n266), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n268), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT81), .B1(new_n264), .B2(new_n266), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n269), .A3(new_n265), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n286), .A2(new_n284), .A3(new_n287), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT82), .B1(new_n291), .B2(KEYINPUT5), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n300), .A3(KEYINPUT83), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n267), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT0), .ZN(new_n304));
  XNOR2_X1  g103(.A(G57gat), .B(G85gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  AOI21_X1  g105(.A(KEYINPUT6), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n302), .B2(KEYINPUT87), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT87), .ZN(new_n310));
  AOI211_X1 g109(.A(new_n310), .B(new_n267), .C1(new_n294), .C2(new_n301), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT24), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n316), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT25), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n320), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(KEYINPUT64), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT64), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n336), .A2(KEYINPUT23), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n325), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n330), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n325), .B(new_n339), .C1(new_n318), .C2(new_n334), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT66), .A3(new_n330), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n329), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n348), .A2(KEYINPUT28), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT28), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n317), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  OR3_X1    g152(.A1(new_n353), .A2(new_n321), .A3(KEYINPUT68), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n322), .A2(KEYINPUT26), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT68), .B1(new_n353), .B2(new_n321), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n346), .A2(new_n347), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n329), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n344), .A2(KEYINPUT66), .A3(new_n330), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT66), .B1(new_n344), .B2(new_n330), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n359), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT78), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n314), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n314), .A2(KEYINPUT29), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n350), .A2(new_n351), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n317), .A4(new_n357), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT69), .B1(new_n352), .B2(new_n358), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT67), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n346), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n374), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n368), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G197gat), .B(G204gat), .Z(new_n379));
  AOI21_X1  g178(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT77), .ZN(new_n382));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n367), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n347), .B1(new_n346), .B2(new_n359), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n364), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n368), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n390), .A2(new_n314), .A3(new_n376), .A4(new_n373), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT37), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(KEYINPUT88), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n389), .A2(new_n391), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n384), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n367), .A2(new_n378), .A3(new_n385), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n404), .B2(new_n396), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT38), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n401), .A2(new_n385), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n367), .A2(new_n378), .A3(new_n384), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT37), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT38), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n402), .A2(new_n403), .A3(new_n396), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n302), .A2(new_n306), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(KEYINPUT6), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n312), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n384), .B1(new_n420), .B2(new_n258), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(G228gat), .B2(G233gat), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT85), .B1(new_n379), .B2(new_n380), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n383), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n381), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n420), .B1(new_n423), .B2(new_n383), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n255), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n259), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n384), .A2(new_n420), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n251), .B1(new_n431), .B2(new_n255), .ZN(new_n432));
  OAI211_X1 g231(.A(G228gat), .B(G233gat), .C1(new_n432), .C2(new_n421), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT31), .B(G50gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n434), .B(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G22gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n437), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n267), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n283), .A2(new_n268), .A3(new_n293), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT83), .B1(new_n297), .B2(new_n300), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n310), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n302), .A2(KEYINPUT87), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n308), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n402), .A2(new_n403), .A3(new_n448), .A4(new_n396), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n397), .B1(new_n386), .B2(new_n392), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n285), .A2(new_n265), .A3(new_n276), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT39), .B(new_n452), .C1(new_n280), .C2(new_n265), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n278), .A2(new_n454), .A3(new_n266), .A4(new_n279), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n455), .A2(KEYINPUT86), .A3(new_n306), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT86), .B1(new_n455), .B2(new_n306), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n453), .B(KEYINPUT40), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  AND4_X1   g260(.A1(new_n449), .A2(new_n451), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n440), .B1(new_n447), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n418), .A2(new_n419), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n419), .B1(new_n418), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n449), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n444), .A2(new_n469), .A3(new_n308), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT84), .B1(new_n302), .B2(new_n306), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n307), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n308), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n440), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT76), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n262), .B1(new_n375), .B2(new_n377), .ZN(new_n478));
  INV_X1    g277(.A(G227gat), .ZN(new_n479));
  INV_X1    g278(.A(G233gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n390), .A2(new_n253), .A3(new_n376), .A4(new_n373), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT73), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT73), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  XOR2_X1   g287(.A(G15gat), .B(G43gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT74), .ZN(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n483), .B2(KEYINPUT32), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n486), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n481), .B1(new_n478), .B2(new_n482), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT34), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n483), .B(KEYINPUT32), .C1(new_n484), .C2(new_n492), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n494), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n477), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(KEYINPUT75), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n494), .A2(new_n497), .ZN(new_n504));
  INV_X1    g303(.A(new_n496), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n503), .B1(new_n508), .B2(new_n477), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n503), .B1(new_n498), .B2(new_n499), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n502), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n476), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n472), .A2(new_n473), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n508), .A2(new_n440), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n467), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n506), .A2(KEYINPUT90), .A3(new_n507), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n312), .A2(new_n473), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n468), .A2(KEYINPUT35), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n521), .A2(new_n475), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n466), .A2(new_n513), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G197gat), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT11), .B(G169gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT12), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(G1gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G1gat), .B2(new_n531), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(G8gat), .Z(new_n535));
  INV_X1    g334(.A(G50gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT15), .B1(new_n536), .B2(G43gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(G43gat), .B2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT94), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT92), .B(KEYINPUT15), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n536), .B2(G43gat), .ZN(new_n544));
  INV_X1    g343(.A(G43gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(G50gat), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n543), .A2(new_n536), .A3(G43gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(KEYINPUT91), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(KEYINPUT14), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n539), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n538), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT95), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT17), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n535), .B(new_n558), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n534), .B(G8gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n530), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n564), .A2(KEYINPUT18), .A3(new_n565), .A4(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n559), .A2(KEYINPUT96), .A3(new_n566), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n535), .A2(new_n557), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(KEYINPUT97), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(KEYINPUT97), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n574), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n565), .B(KEYINPUT13), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n570), .A2(new_n573), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n572), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n568), .A2(new_n569), .B1(new_n580), .B2(new_n581), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT98), .B1(new_n568), .B2(new_n569), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n585), .B(new_n573), .C1(new_n586), .C2(new_n530), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n525), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n472), .A2(new_n473), .ZN(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT102), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n593), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n558), .B(new_n602), .C1(new_n561), .C2(new_n563), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n559), .A2(new_n601), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n606), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G64gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  OR2_X1    g418(.A1(G71gat), .A2(G78gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT9), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n624));
  AND2_X1   g423(.A1(G57gat), .A2(G64gat), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n619), .B(new_n620), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n566), .B1(KEYINPUT21), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G155gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n631), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G127gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n634), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n616), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT104), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n601), .A2(new_n628), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n593), .A2(new_n600), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n593), .A2(new_n600), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n627), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n651), .B1(new_n653), .B2(new_n657), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n650), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT105), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT103), .B(new_n652), .C1(new_n658), .C2(new_n659), .ZN(new_n666));
  INV_X1    g465(.A(new_n649), .ZN(new_n667));
  OR4_X1    g466(.A1(new_n665), .A2(new_n666), .A3(new_n661), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n646), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n590), .A2(new_n591), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT106), .B(G1gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND4_X1  g473(.A1(new_n590), .A2(new_n468), .A3(new_n670), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n512), .ZN(new_n676));
  INV_X1    g475(.A(new_n415), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n408), .A2(new_n473), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n441), .B(new_n306), .C1(new_n442), .C2(new_n443), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT6), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n306), .B1(new_n444), .B2(new_n310), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n446), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n462), .B1(new_n311), .B2(new_n309), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n475), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT89), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n440), .B1(new_n591), .B2(new_n468), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n418), .A2(new_n419), .A3(new_n463), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n676), .A2(new_n687), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n517), .A2(new_n524), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n692), .A2(new_n588), .A3(new_n468), .A4(new_n670), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G8gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT42), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n675), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1325gat));
  NAND2_X1  g502(.A1(new_n590), .A2(new_n670), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n704), .B2(new_n676), .ZN(new_n705));
  INV_X1    g504(.A(G15gat), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n590), .A2(new_n706), .A3(new_n521), .A4(new_n670), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n704), .A2(new_n475), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(new_n669), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n644), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n616), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT108), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n514), .A2(G29gat), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n692), .A2(new_n588), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n525), .B2(new_n616), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n615), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n713), .A2(new_n589), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n721), .A2(new_n722), .A3(new_n591), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G29gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1328gat));
  NAND2_X1  g527(.A1(new_n590), .A2(new_n715), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(G36gat), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n468), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n721), .A2(new_n722), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n468), .A3(new_n723), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G36gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(G1329gat));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n722), .A3(new_n512), .A4(new_n723), .ZN(new_n740));
  INV_X1    g539(.A(new_n521), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  AOI22_X1  g541(.A1(G43gat), .A2(new_n740), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n744));
  OAI21_X1  g543(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n744), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n740), .A2(G43gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n729), .A2(G43gat), .A3(new_n741), .ZN(new_n748));
  OAI211_X1 g547(.A(KEYINPUT113), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(G1330gat));
  NAND3_X1  g550(.A1(new_n730), .A2(new_n536), .A3(new_n440), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n721), .A2(new_n722), .A3(new_n440), .A4(new_n723), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1331gat));
  NOR3_X1   g556(.A1(new_n525), .A2(new_n588), .A3(new_n646), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n669), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n514), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g560(.A1(new_n467), .A2(new_n712), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT49), .B(G64gat), .Z(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n676), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n758), .A2(new_n669), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n758), .A2(new_n771), .A3(new_n669), .A4(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n767), .B1(new_n759), .B2(new_n741), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n759), .A2(new_n475), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g579(.A1(new_n645), .A2(new_n588), .A3(new_n712), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n735), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n514), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n645), .A2(new_n588), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT76), .B1(new_n506), .B2(new_n507), .ZN(new_n785));
  OAI211_X1 g584(.A(KEYINPUT36), .B(new_n510), .C1(new_n785), .C2(new_n503), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n502), .C1(new_n474), .C2(new_n475), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n787), .A2(new_n464), .A3(new_n465), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n517), .A2(new_n524), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n615), .B(new_n784), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n616), .B1(new_n690), .B2(new_n691), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n712), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n597), .A3(new_n591), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n783), .A2(new_n796), .ZN(G1336gat));
  NAND4_X1  g596(.A1(new_n721), .A2(new_n722), .A3(new_n468), .A4(new_n781), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n790), .A2(new_n791), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n793), .B2(new_n784), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n598), .B(new_n762), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n782), .B2(new_n676), .ZN(new_n805));
  INV_X1    g604(.A(new_n795), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n741), .A2(G99gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(G1338gat));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n721), .A2(new_n722), .A3(new_n440), .A4(new_n781), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n475), .A2(G106gat), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n669), .B(new_n812), .C1(new_n800), .C2(new_n801), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n814));
  AND4_X1   g613(.A1(new_n809), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n795), .A2(new_n812), .B1(new_n810), .B2(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n809), .B1(new_n816), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n811), .A2(new_n813), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n815), .B1(new_n817), .B2(new_n819), .ZN(G1339gat));
  NAND3_X1  g619(.A1(new_n585), .A2(new_n530), .A3(new_n573), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n580), .A2(new_n581), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n565), .B1(new_n564), .B2(new_n567), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n529), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n669), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n658), .A2(new_n652), .A3(new_n659), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n665), .A2(new_n666), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n649), .B1(new_n660), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n660), .B(new_n664), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT55), .B(new_n832), .C1(new_n835), .C2(new_n829), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n836), .A3(new_n668), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n826), .B1(new_n589), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n616), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n834), .A2(new_n836), .A3(new_n668), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n615), .A2(new_n825), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n645), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n646), .A2(new_n588), .A3(new_n669), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n440), .A3(new_n741), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n591), .A3(new_n467), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n221), .A3(new_n589), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n844), .A2(new_n514), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n515), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n467), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n588), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n847), .B1(new_n851), .B2(new_n221), .ZN(G1340gat));
  NOR3_X1   g651(.A1(new_n846), .A2(new_n219), .A3(new_n712), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n669), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n219), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n204), .A3(new_n645), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n846), .B2(new_n644), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  NAND4_X1  g657(.A1(new_n849), .A2(new_n206), .A3(new_n467), .A4(new_n615), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(KEYINPUT56), .A3(new_n861), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n846), .B2(new_n616), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n844), .B2(new_n475), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n837), .A2(KEYINPUT119), .B1(new_n584), .B2(new_n587), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n834), .A2(new_n836), .A3(new_n871), .A4(new_n668), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n615), .B1(new_n873), .B2(new_n826), .ZN(new_n874));
  INV_X1    g673(.A(new_n841), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n644), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n843), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n475), .A2(new_n868), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n869), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n512), .A2(new_n514), .A3(new_n468), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n232), .B1(new_n883), .B2(new_n588), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n512), .A2(new_n475), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n848), .A2(new_n467), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G141gat), .A3(new_n589), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT58), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(KEYINPUT120), .A3(new_n588), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n881), .A2(new_n882), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n589), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n891), .A2(G141gat), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n890), .B2(new_n895), .ZN(G1344gat));
  NOR2_X1   g695(.A1(new_n234), .A2(KEYINPUT59), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n883), .B2(new_n669), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n870), .A2(new_n872), .B1(new_n669), .B2(new_n825), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n841), .B1(new_n901), .B2(new_n615), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n843), .B1(new_n902), .B2(new_n644), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n868), .B1(new_n903), .B2(new_n475), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n879), .B1(new_n842), .B2(new_n843), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n712), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n234), .B1(new_n906), .B2(new_n882), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n475), .B1(new_n876), .B2(new_n877), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n669), .A3(new_n882), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G148gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n899), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n887), .A2(G148gat), .A3(new_n712), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT122), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n897), .B1(new_n893), .B2(new_n712), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT121), .B1(new_n913), .B2(KEYINPUT59), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n900), .B(new_n908), .C1(new_n912), .C2(G148gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  INV_X1    g721(.A(new_n916), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n917), .A2(new_n924), .ZN(G1345gat));
  AOI21_X1  g724(.A(G155gat), .B1(new_n886), .B2(new_n645), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n645), .A2(G155gat), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n883), .B2(new_n928), .ZN(G1346gat));
  NAND4_X1  g728(.A1(new_n886), .A2(new_n241), .A3(new_n243), .A4(new_n615), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n883), .A2(KEYINPUT124), .A3(new_n615), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n244), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT124), .B1(new_n883), .B2(new_n615), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n844), .A2(new_n591), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n468), .A3(new_n515), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n588), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n591), .A2(new_n467), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n845), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n845), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n589), .A2(new_n337), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n938), .B1(new_n944), .B2(new_n945), .ZN(G1348gat));
  AOI21_X1  g745(.A(G176gat), .B1(new_n937), .B2(new_n669), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n712), .B1(new_n336), .B2(new_n338), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n944), .B2(new_n948), .ZN(G1349gat));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n645), .A3(new_n943), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G183gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n937), .A2(new_n348), .A3(new_n645), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n349), .A3(new_n615), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n944), .A2(new_n615), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(G190gat), .ZN(new_n958));
  AOI211_X1 g757(.A(KEYINPUT61), .B(new_n349), .C1(new_n944), .C2(new_n615), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NAND3_X1  g759(.A1(new_n935), .A2(new_n468), .A3(new_n885), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n588), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n676), .A2(new_n939), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT126), .Z(new_n965));
  AOI21_X1  g764(.A(new_n965), .B1(new_n904), .B2(new_n905), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n588), .A2(G197gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n935), .A2(new_n969), .A3(new_n762), .A4(new_n885), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  INV_X1    g770(.A(new_n906), .ZN(new_n972));
  OAI21_X1  g771(.A(G204gat), .B1(new_n972), .B2(new_n965), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1353gat));
  INV_X1    g773(.A(G211gat), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n964), .A2(new_n644), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n911), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT63), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n975), .A3(new_n645), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1354gat));
  AOI21_X1  g779(.A(G218gat), .B1(new_n962), .B2(new_n615), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n615), .A2(G218gat), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n982), .A2(new_n983), .B1(new_n966), .B2(new_n984), .ZN(G1355gat));
endmodule


