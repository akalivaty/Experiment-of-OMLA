//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n540, new_n541, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n589, new_n592, new_n593, new_n595, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT67), .ZN(new_n477));
  MUX2_X1   g052(.A(G100), .B(G112), .S(G2105), .Z(new_n478));
  AOI22_X1  g053(.A1(G136), .A2(new_n467), .B1(new_n478), .B2(G2104), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(G162));
  NAND3_X1  g055(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(G114), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G102), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n481), .A2(KEYINPUT68), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT68), .B1(new_n481), .B2(new_n485), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n467), .B2(G138), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n468), .C1(new_n459), .C2(new_n460), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  OAI22_X1  g066(.A1(new_n486), .A2(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  AND2_X1   g068(.A1(KEYINPUT6), .A2(G651), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT6), .A2(G651), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G50), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n495), .B2(new_n494), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n497), .A2(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n504), .A2(new_n507), .ZN(G166));
  NAND3_X1  g083(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n509));
  INV_X1    g084(.A(G51), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n497), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n496), .A2(new_n501), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G89), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT69), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT7), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n513), .A2(new_n517), .A3(KEYINPUT70), .A4(new_n518), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(G168));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n497), .A2(new_n524), .B1(new_n502), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n506), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n526), .A2(new_n528), .ZN(G301));
  INV_X1    g104(.A(G301), .ZN(G171));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT71), .B(G81), .Z(new_n532));
  OAI22_X1  g107(.A1(new_n497), .A2(new_n531), .B1(new_n502), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n506), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  AND3_X1   g112(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G36), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G188));
  AOI22_X1  g117(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n506), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n512), .A2(G91), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n496), .A2(G53), .A3(G543), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n546), .A2(KEYINPUT9), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(KEYINPUT9), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n544), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(G299));
  NAND2_X1  g124(.A1(new_n521), .A2(new_n522), .ZN(new_n550));
  INV_X1    g125(.A(new_n511), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G286));
  INV_X1    g127(.A(G166), .ZN(G303));
  INV_X1    g128(.A(new_n497), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G49), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n512), .A2(G87), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(G288));
  OAI211_X1 g133(.A(G48), .B(G543), .C1(new_n494), .C2(new_n495), .ZN(new_n559));
  INV_X1    g134(.A(G86), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n502), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n499), .B2(new_n500), .ZN(new_n563));
  AND2_X1   g138(.A1(G73), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G305));
  INV_X1    g143(.A(G47), .ZN(new_n569));
  INV_X1    g144(.A(G85), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n497), .A2(new_n569), .B1(new_n502), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n506), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  INV_X1    g150(.A(G92), .ZN(new_n576));
  XOR2_X1   g151(.A(KEYINPUT72), .B(KEYINPUT10), .Z(new_n577));
  OR3_X1    g152(.A1(new_n502), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n502), .B2(new_n576), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n501), .A2(G66), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n506), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(G54), .B2(new_n554), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  MUX2_X1   g161(.A(G301), .B(new_n585), .S(new_n586), .Z(G284));
  MUX2_X1   g162(.A(G301), .B(new_n585), .S(new_n586), .Z(G321));
  NOR2_X1   g163(.A1(G299), .A2(G868), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g165(.A(new_n589), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g166(.A(new_n585), .ZN(new_n592));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(G860), .ZN(G148));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n536), .A2(new_n586), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT11), .Z(G282));
  INV_X1    g173(.A(new_n597), .ZN(G323));
  MUX2_X1   g174(.A(G99), .B(G111), .S(G2105), .Z(new_n600));
  AOI22_X1  g175(.A1(new_n475), .A2(G123), .B1(G2104), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G135), .ZN(new_n602));
  INV_X1    g177(.A(new_n467), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT75), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(G2096), .Z(new_n606));
  NAND2_X1  g181(.A1(new_n467), .A2(G2104), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n608), .A2(new_n609), .B1(KEYINPUT74), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n608), .B2(new_n609), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n612), .A2(KEYINPUT74), .A3(new_n610), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(KEYINPUT74), .B2(new_n610), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n606), .A2(new_n613), .A3(new_n614), .ZN(G156));
  INV_X1    g190(.A(G14), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT14), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT15), .B(G2435), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2427), .ZN(new_n620));
  INV_X1    g195(.A(G2430), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n620), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n616), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n623), .B2(new_n629), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT76), .Z(G401));
  XOR2_X1   g207(.A(G2084), .B(G2090), .Z(new_n633));
  XNOR2_X1  g208(.A(G2072), .B(G2078), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n633), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n634), .A2(KEYINPUT17), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n635), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n633), .A2(new_n635), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n634), .B1(new_n644), .B2(KEYINPUT17), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n638), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2096), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT78), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  OR2_X1    g234(.A1(new_n652), .A2(new_n654), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(new_n657), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n657), .A3(new_n655), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT23), .ZN(new_n673));
  INV_X1    g248(.A(G299), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n671), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1956), .ZN(new_n676));
  NOR2_X1   g251(.A1(G171), .A2(new_n671), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G5), .B2(new_n671), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n605), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n679), .A2(G1961), .B1(new_n680), .B2(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n682), .A2(new_n683), .B1(new_n469), .B2(G105), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n683), .B2(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n467), .A2(G141), .ZN(new_n686));
  INV_X1    g261(.A(G129), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n474), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n690), .B2(G32), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT27), .B(G1996), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G2084), .ZN(new_n696));
  INV_X1    g271(.A(G34), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(KEYINPUT24), .ZN(new_n698));
  AOI21_X1  g273(.A(G29), .B1(new_n697), .B2(KEYINPUT24), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(KEYINPUT89), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(KEYINPUT89), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n471), .B2(new_n690), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n693), .A2(new_n695), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G2078), .ZN(new_n704));
  NAND2_X1  g279(.A1(G164), .A2(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G27), .B2(G29), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n681), .B(new_n703), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  AOI211_X1 g282(.A(new_n676), .B(new_n707), .C1(new_n704), .C2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G11), .ZN(new_n709));
  INV_X1    g284(.A(G28), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n710), .B2(KEYINPUT30), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT91), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n713), .A2(new_n710), .A3(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(new_n710), .B2(KEYINPUT30), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n709), .B1(new_n712), .B2(new_n717), .C1(new_n679), .C2(G1961), .ZN(new_n718));
  NOR2_X1   g293(.A1(G29), .A2(G33), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n469), .A2(G103), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT25), .Z(new_n722));
  INV_X1    g297(.A(G139), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n603), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n468), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n720), .B1(new_n728), .B2(new_n690), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G2072), .Z(new_n730));
  NOR2_X1   g305(.A1(new_n693), .A2(new_n695), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n702), .A2(new_n696), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n718), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n592), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT85), .B(G1348), .Z(new_n736));
  XOR2_X1   g311(.A(new_n735), .B(new_n736), .Z(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n536), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1341), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n690), .A2(G26), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT86), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n467), .A2(G140), .ZN(new_n744));
  MUX2_X1   g319(.A(G104), .B(G116), .S(G2105), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G2104), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n473), .A2(G128), .A3(G2105), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n690), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2067), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n737), .A2(new_n740), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n671), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n671), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(G1966), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n708), .A2(new_n733), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G162), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2090), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n752), .A2(new_n753), .B1(G1966), .B2(new_n755), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n757), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n671), .A2(G23), .ZN(new_n766));
  INV_X1    g341(.A(G288), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n671), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT33), .B(G1976), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G22), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G166), .B2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1971), .Z(new_n773));
  NOR2_X1   g348(.A1(G6), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n567), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n770), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT34), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(KEYINPUT34), .ZN(new_n780));
  INV_X1    g355(.A(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT81), .B1(new_n781), .B2(G16), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n781), .A2(KEYINPUT81), .A3(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n574), .B(KEYINPUT82), .Z(new_n784));
  OAI211_X1 g359(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n671), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT83), .B(G1986), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n467), .A2(G131), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT80), .Z(new_n789));
  MUX2_X1   g364(.A(G95), .B(G107), .S(G2105), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n475), .A2(G119), .B1(G2104), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G25), .B(new_n792), .S(G29), .Z(new_n793));
  XOR2_X1   g368(.A(KEYINPUT35), .B(G1991), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n779), .A2(new_n780), .A3(new_n787), .A4(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT84), .B(KEYINPUT36), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n765), .A2(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  AOI22_X1  g375(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(new_n506), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n512), .A2(G93), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT94), .B(G55), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n496), .A2(new_n805), .A3(G543), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n806), .B1(new_n808), .B2(new_n502), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(KEYINPUT95), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n802), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G860), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  INV_X1    g388(.A(new_n536), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n536), .B(new_n802), .C1(new_n807), .C2(new_n810), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n585), .A2(new_n593), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT96), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT97), .Z(new_n824));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n825));
  AOI21_X1  g400(.A(G860), .B1(new_n821), .B2(new_n822), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n825), .B1(new_n824), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n813), .B1(new_n827), .B2(new_n828), .ZN(G145));
  XOR2_X1   g404(.A(new_n605), .B(G162), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n471), .B(KEYINPUT99), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n830), .B(new_n831), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n481), .A2(new_n485), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n473), .A2(new_n488), .A3(G138), .A4(new_n468), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n748), .ZN(new_n842));
  INV_X1    g417(.A(new_n689), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n749), .B(new_n835), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT100), .B1(new_n489), .B2(new_n491), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n749), .B1(new_n851), .B2(new_n835), .ZN(new_n852));
  AOI211_X1 g427(.A(new_n834), .B(new_n748), .C1(new_n849), .C2(new_n850), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n689), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT101), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n727), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n728), .A3(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n475), .A2(G130), .B1(G142), .B2(new_n467), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n864), .B(new_n865), .C1(G118), .C2(new_n468), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(new_n608), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n792), .ZN(new_n869));
  OAI211_X1 g444(.A(KEYINPUT102), .B(new_n727), .C1(new_n848), .C2(new_n856), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n860), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n860), .B2(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI211_X1 g449(.A(KEYINPUT104), .B(new_n869), .C1(new_n860), .C2(new_n870), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n833), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g453(.A(KEYINPUT105), .B(new_n833), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n832), .B(new_n871), .C1(new_n872), .C2(KEYINPUT106), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n872), .A2(KEYINPUT106), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT40), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n887));
  AOI211_X1 g462(.A(new_n887), .B(new_n884), .C1(new_n878), .C2(new_n879), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n886), .A2(new_n888), .ZN(G395));
  NOR2_X1   g464(.A1(new_n811), .A2(G868), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n585), .A2(G299), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n585), .A2(G299), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT41), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n674), .A2(new_n580), .A3(new_n584), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n892), .A2(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n592), .A2(new_n593), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n817), .B(new_n900), .ZN(new_n901));
  MUX2_X1   g476(.A(new_n898), .B(new_n899), .S(new_n901), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT42), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n574), .B(G288), .Z(new_n904));
  XNOR2_X1  g479(.A(G166), .B(new_n567), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n903), .B(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n890), .B1(new_n907), .B2(G868), .ZN(G295));
  AOI21_X1  g483(.A(new_n890), .B1(new_n907), .B2(G868), .ZN(G331));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(G286), .A2(G301), .ZN(new_n911));
  NAND2_X1  g486(.A1(G168), .A2(G171), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n815), .A3(new_n816), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(G168), .A2(G171), .ZN(new_n914));
  AOI211_X1 g489(.A(new_n511), .B(G301), .C1(new_n521), .C2(new_n522), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n817), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n913), .A2(new_n916), .A3(new_n899), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n916), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n898), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n906), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n897), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n895), .A2(new_n891), .A3(KEYINPUT108), .A4(new_n896), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n894), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT109), .B1(new_n918), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(new_n917), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n924), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n906), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI211_X1 g505(.A(KEYINPUT110), .B(new_n906), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n906), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n919), .A2(KEYINPUT107), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n919), .A2(KEYINPUT107), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n920), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n910), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n930), .B2(new_n931), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(KEYINPUT43), .A3(new_n920), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT44), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n939), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT45), .B1(new_n841), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n464), .A2(G40), .A3(new_n470), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(G1996), .A3(new_n843), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT111), .Z(new_n950));
  NOR2_X1   g525(.A1(new_n947), .A2(G1996), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n748), .B(G2067), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n951), .A2(new_n689), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n792), .B(new_n794), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n947), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n574), .B(G1986), .Z(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT115), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n492), .A2(new_n944), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n962));
  NAND3_X1  g537(.A1(new_n841), .A2(new_n944), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n946), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n964), .B2(G2084), .ZN(new_n965));
  INV_X1    g540(.A(new_n946), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n967), .A2(KEYINPUT115), .A3(new_n696), .A4(new_n963), .ZN(new_n968));
  INV_X1    g543(.A(G1966), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n946), .B1(new_n960), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n971), .B2(new_n945), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G8), .B1(new_n973), .B2(G286), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT51), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n973), .B2(G286), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT62), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n975), .B(new_n980), .C1(new_n974), .C2(new_n977), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT55), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n966), .B1(new_n960), .B2(new_n970), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n841), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n986));
  AOI21_X1  g561(.A(G1971), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n946), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n841), .A2(new_n944), .ZN(new_n989));
  INV_X1    g564(.A(new_n962), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n991), .B2(new_n762), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n964), .A2(G2090), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n983), .B(G8), .C1(new_n995), .C2(new_n987), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n512), .A2(G86), .ZN(new_n997));
  INV_X1    g572(.A(G1981), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n565), .A4(new_n559), .ZN(new_n999));
  OAI21_X1  g574(.A(G1981), .B1(new_n561), .B2(new_n566), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(KEYINPUT114), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(G1981), .C1(new_n561), .C2(new_n566), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n841), .A2(new_n946), .A3(new_n944), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n767), .A2(G1976), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(KEYINPUT113), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1010), .A2(new_n1007), .A3(G8), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  NAND3_X1  g589(.A1(G288), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(new_n1007), .A3(G8), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(KEYINPUT113), .B2(new_n1011), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1009), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n994), .A2(new_n996), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n985), .A2(new_n986), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(G2078), .ZN(new_n1023));
  INV_X1    g598(.A(G1961), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n964), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n704), .A2(KEYINPUT53), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n971), .A2(new_n945), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G171), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1020), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n979), .A2(new_n981), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n1032));
  INV_X1    g607(.A(new_n996), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1008), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n767), .A2(new_n1014), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n999), .B1(new_n1009), .B2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1033), .A2(new_n1019), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G286), .A2(new_n993), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n973), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n973), .A2(KEYINPUT116), .A3(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1019), .A2(new_n996), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1022), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n989), .A2(new_n990), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n946), .C1(KEYINPUT50), .C2(new_n960), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1046), .A2(G1971), .B1(new_n1048), .B2(G2090), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n983), .B1(new_n1049), .B2(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1038), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n995), .B2(new_n987), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n984), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1054), .A2(KEYINPUT63), .A3(new_n1019), .A4(new_n996), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1032), .B(new_n1037), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1046), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1048), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(KEYINPUT119), .ZN(new_n1064));
  MUX2_X1   g639(.A(new_n1062), .B(new_n1064), .S(G299), .Z(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1059), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G2067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1007), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n964), .A2(new_n736), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n585), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1065), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1067), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1066), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT58), .B(G1341), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1022), .A2(G1996), .B1(new_n1069), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n536), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n1083));
  NAND2_X1  g658(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n536), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1070), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(new_n592), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1071), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n585), .ZN(new_n1090));
  AND4_X1   g665(.A1(new_n1079), .A2(new_n1086), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1067), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1074), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n1067), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1075), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n704), .A2(KEYINPUT124), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n704), .A2(KEYINPUT124), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT53), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n463), .B(KEYINPUT122), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G2105), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(G40), .A3(new_n470), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1103), .B2(KEYINPUT123), .ZN(new_n1104));
  INV_X1    g679(.A(new_n945), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(new_n1106), .A3(G40), .A4(new_n470), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1104), .A2(new_n986), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(G301), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1109), .A2(KEYINPUT125), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(KEYINPUT125), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1029), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1023), .A2(new_n1027), .A3(G301), .A4(new_n1025), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1108), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n1118), .B2(G171), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1020), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(new_n1120), .A3(new_n978), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1031), .B(new_n1057), .C1(new_n1097), .C2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1032), .B1(new_n1123), .B2(new_n1037), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n958), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n954), .A2(new_n789), .A3(new_n791), .A4(new_n794), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n749), .A2(new_n1068), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n947), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n948), .B1(new_n843), .B2(new_n952), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT47), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n947), .A2(G1986), .A3(G290), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT48), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n956), .B2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1125), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g713(.A1(new_n631), .A2(new_n649), .A3(G319), .ZN(new_n1140));
  NAND2_X1  g714(.A1(new_n669), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n1142));
  XNOR2_X1  g716(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  NAND3_X1  g717(.A1(new_n940), .A2(new_n1143), .A3(new_n941), .ZN(new_n1144));
  AOI21_X1  g718(.A(new_n884), .B1(new_n878), .B2(new_n879), .ZN(new_n1145));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n1145), .ZN(G308));
  OR2_X1    g720(.A1(new_n1144), .A2(new_n1145), .ZN(G225));
endmodule


