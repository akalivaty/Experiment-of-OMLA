//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n204));
  INV_X1    g0004(.A(G87), .ZN(new_n205));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n203), .B1(new_n210), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n203), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(new_n213), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n219), .A2(new_n222), .A3(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(G270), .Z(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  OAI211_X1 g0047(.A(G1), .B(G13), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT5), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT77), .B1(new_n249), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT77), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(new_n247), .A3(KEYINPUT5), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n249), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(G270), .B(new_n248), .C1(new_n253), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT80), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n250), .A2(new_n252), .A3(new_n256), .A4(new_n255), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT80), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(G270), .A4(new_n248), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G45), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n267), .A2(G274), .A3(new_n250), .A4(new_n252), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n269));
  OR2_X1    g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT81), .B(G303), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G264), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n208), .B2(G1698), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n268), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n263), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n226), .A3(G1), .ZN(new_n285));
  INV_X1    g0085(.A(G116), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n227), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n265), .A2(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G116), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(G20), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G283), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n226), .C1(G33), .C2(new_n207), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT20), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AND4_X1   g0097(.A1(KEYINPUT20), .A2(new_n296), .A3(new_n289), .A4(new_n293), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n287), .B(new_n292), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  AND4_X1   g0099(.A1(KEYINPUT21), .A2(new_n283), .A3(G169), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n263), .B2(new_n282), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT21), .B1(new_n302), .B2(new_n299), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT82), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n263), .A2(G179), .A3(new_n282), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n299), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n263), .A2(new_n282), .A3(G190), .ZN(new_n308));
  INV_X1    g0108(.A(new_n299), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n281), .B1(new_n259), .B2(new_n262), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n283), .A2(G169), .A3(new_n299), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT21), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n302), .A2(KEYINPUT21), .A3(new_n299), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n307), .A3(new_n312), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT82), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  OAI211_X1 g0121(.A(G244), .B(new_n321), .C1(new_n275), .C2(new_n276), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT76), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n272), .A2(G244), .A3(new_n321), .A4(new_n324), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n295), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n269), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n260), .A2(G257), .A3(new_n248), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n268), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n290), .A2(new_n291), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n207), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT7), .B1(new_n277), .B2(new_n226), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  NOR4_X1   g0137(.A1(new_n275), .A2(new_n276), .A3(new_n337), .A4(G20), .ZN(new_n338));
  OAI21_X1  g0138(.A(G107), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G20), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n215), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT6), .ZN(new_n344));
  INV_X1    g0144(.A(G107), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n207), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G97), .A2(G107), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(KEYINPUT6), .A3(G97), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n339), .B(new_n343), .C1(new_n226), .C2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n335), .B1(new_n351), .B2(new_n289), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n285), .A2(new_n207), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n330), .A2(new_n331), .A3(G190), .A4(new_n268), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n333), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT78), .A2(G250), .ZN(new_n356));
  INV_X1    g0156(.A(G274), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n255), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT78), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n266), .A2(new_n360), .A3(G250), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n248), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G116), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n270), .A2(new_n271), .B1(new_n216), .B2(G1698), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n214), .A2(new_n321), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n363), .B(G190), .C1(new_n368), .C2(new_n248), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n347), .A2(new_n205), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n226), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT19), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n226), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT19), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n371), .B2(G20), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n377), .A2(new_n289), .B1(new_n285), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n216), .A2(G1698), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n367), .B(new_n380), .C1(new_n275), .C2(new_n276), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n248), .B1(new_n381), .B2(new_n364), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n269), .B1(new_n359), .B2(new_n361), .ZN(new_n383));
  OAI21_X1  g0183(.A(G200), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n290), .A2(G87), .A3(new_n291), .ZN(new_n385));
  AND4_X1   g0185(.A1(new_n369), .A2(new_n379), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n382), .A2(new_n383), .ZN(new_n387));
  INV_X1    g0187(.A(G179), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT79), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT79), .ZN(new_n390));
  NOR4_X1   g0190(.A1(new_n382), .A2(new_n383), .A3(new_n390), .A4(G179), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n334), .A2(new_n378), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n363), .B1(new_n368), .B2(new_n248), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n379), .A2(new_n393), .B1(new_n394), .B2(new_n301), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n386), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n332), .A2(new_n301), .ZN(new_n397));
  INV_X1    g0197(.A(new_n335), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n270), .A2(new_n226), .A3(new_n271), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n337), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n271), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n345), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n226), .B1(new_n348), .B2(new_n349), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n402), .A2(new_n403), .A3(new_n342), .ZN(new_n404));
  INV_X1    g0204(.A(new_n289), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n353), .B(new_n398), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n330), .A2(new_n331), .A3(new_n388), .A4(new_n268), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n355), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n334), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G107), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n285), .A2(new_n345), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT85), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT24), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT83), .B1(new_n364), .B2(G20), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT83), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n420), .A2(new_n226), .A3(G33), .A4(G116), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT23), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n226), .B2(G107), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n345), .A2(KEYINPUT23), .A3(G20), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n422), .A2(KEYINPUT84), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT84), .B1(new_n422), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n226), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT22), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n418), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(new_n426), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT84), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n422), .A2(KEYINPUT84), .A3(new_n426), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n418), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n430), .B(KEYINPUT22), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n417), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n411), .B(new_n414), .C1(new_n442), .C2(new_n405), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n206), .A2(new_n321), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n208), .A2(G1698), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(new_n275), .C2(new_n276), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G294), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n269), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n260), .A2(G264), .A3(new_n248), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n450), .A2(new_n268), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G190), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(G200), .B2(new_n452), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n409), .B1(new_n444), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(G169), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n388), .B2(new_n452), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n443), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n320), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n265), .A2(G20), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT67), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G50), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(KEYINPUT68), .A3(G50), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n290), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(G20), .B1(new_n224), .B2(G50), .ZN(new_n469));
  INV_X1    g0269(.A(G150), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT8), .B(G58), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n226), .A2(G33), .ZN(new_n472));
  OAI221_X1 g0272(.A(new_n469), .B1(new_n470), .B2(new_n341), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G50), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n473), .A2(new_n289), .B1(new_n474), .B2(new_n285), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT9), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n321), .A2(G222), .ZN(new_n478));
  INV_X1    g0278(.A(G223), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n272), .B(new_n478), .C1(new_n479), .C2(new_n321), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n269), .C1(G77), .C2(new_n272), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(new_n357), .ZN(new_n483));
  INV_X1    g0283(.A(G226), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n248), .A2(new_n482), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n486), .A2(new_n453), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(G200), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT70), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT10), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(KEYINPUT70), .A3(G200), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n477), .A2(new_n487), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n476), .A2(KEYINPUT9), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT9), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n468), .B2(new_n475), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n487), .B(new_n488), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT10), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n486), .A2(G179), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n486), .A2(new_n301), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n476), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT16), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n213), .B1(new_n400), .B2(new_n401), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n223), .A2(new_n213), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G58), .A2(G68), .ZN(new_n506));
  OAI21_X1  g0306(.A(G20), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n340), .A2(G159), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n503), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(G68), .B1(new_n336), .B2(new_n338), .ZN(new_n511));
  INV_X1    g0311(.A(new_n509), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(KEYINPUT16), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n513), .A3(new_n289), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n471), .A2(new_n285), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n463), .A2(new_n290), .ZN(new_n516));
  INV_X1    g0316(.A(new_n471), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n479), .A2(new_n321), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n484), .A2(G1698), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n275), .C2(new_n276), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n269), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n248), .A2(G232), .A3(new_n482), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(new_n388), .A3(new_n526), .A4(new_n483), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT74), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n482), .A2(new_n357), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n524), .B2(new_n269), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n526), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n301), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n519), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n519), .A2(new_n529), .A3(new_n533), .A4(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT17), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n531), .A2(G190), .A3(new_n526), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n514), .A2(new_n540), .A3(new_n515), .A4(new_n518), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(KEYINPUT17), .A3(new_n542), .A4(new_n540), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n538), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n502), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G238), .A2(G1698), .ZN(new_n549));
  INV_X1    g0349(.A(G232), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n272), .B(new_n549), .C1(new_n550), .C2(G1698), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n551), .B(new_n269), .C1(G107), .C2(new_n272), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n483), .C1(new_n216), .C2(new_n485), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n517), .A2(new_n340), .B1(G20), .B2(G77), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n472), .B2(new_n378), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n289), .B1(G77), .B2(new_n516), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n285), .A2(new_n215), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT69), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n553), .A2(new_n453), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n553), .A2(G200), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT69), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n558), .A4(new_n557), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n516), .A2(G68), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT73), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n284), .A2(G1), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n226), .A2(G68), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n341), .A2(new_n474), .B1(new_n472), .B2(new_n215), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n289), .B1(new_n572), .B2(new_n569), .ZN(new_n573));
  XOR2_X1   g0373(.A(KEYINPUT72), .B(KEYINPUT11), .Z(new_n574));
  XNOR2_X1  g0374(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n550), .A2(G1698), .ZN(new_n577));
  OAI221_X1 g0377(.A(new_n577), .B1(G226), .B2(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n371), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n269), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n248), .A2(new_n482), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n530), .B1(new_n581), .B2(G238), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT13), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT71), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n248), .B1(new_n578), .B2(new_n371), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n483), .B1(new_n485), .B2(new_n214), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT13), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT71), .A4(new_n583), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(G169), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT14), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT14), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n589), .A2(new_n593), .A3(G169), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n584), .A2(new_n588), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n388), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n576), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n589), .A2(G200), .A3(new_n590), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n596), .A2(new_n453), .ZN(new_n600));
  OR3_X1    g0400(.A1(new_n576), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n553), .A2(G179), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n553), .A2(new_n301), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n559), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n598), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n565), .A4(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT75), .ZN(new_n608));
  INV_X1    g0408(.A(new_n501), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n492), .B2(new_n497), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n546), .A2(new_n544), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n610), .A2(new_n612), .A3(new_n538), .A4(new_n565), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n608), .B1(new_n613), .B2(new_n605), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n460), .B1(new_n607), .B2(new_n614), .ZN(G372));
  NAND2_X1  g0415(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  INV_X1    g0416(.A(new_n455), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n443), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n393), .A2(new_n379), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n394), .A2(new_n301), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n387), .A2(new_n388), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n369), .A2(new_n379), .A3(new_n384), .A4(new_n385), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n355), .A2(new_n624), .A3(new_n408), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT87), .B1(new_n618), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n459), .A2(new_n307), .A3(new_n304), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n355), .A2(new_n624), .A3(new_n408), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n429), .A2(new_n418), .A3(new_n432), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n415), .B2(new_n416), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n289), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n411), .A3(new_n414), .A4(new_n455), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n622), .B(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n622), .A2(new_n623), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n408), .A2(KEYINPUT26), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n397), .A2(new_n407), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n406), .A3(new_n396), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n637), .B(new_n639), .C1(KEYINPUT26), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n616), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n538), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n536), .A2(KEYINPUT89), .A3(new_n537), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n604), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n601), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n598), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n651), .B2(new_n611), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n609), .B1(new_n652), .B2(new_n498), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(G369));
  XNOR2_X1  g0454(.A(new_n318), .B(new_n305), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n568), .A2(new_n226), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT27), .ZN(new_n658));
  INV_X1    g0458(.A(G213), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n656), .B2(KEYINPUT27), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n657), .B1(new_n656), .B2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(new_n309), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n304), .A2(new_n307), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT91), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(KEYINPUT91), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n633), .B1(new_n444), .B2(new_n665), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n459), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n443), .A2(new_n458), .A3(new_n665), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n668), .A2(new_n665), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n676), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n220), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G1), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n347), .A2(new_n205), .A3(new_n286), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n688), .A2(new_n689), .B1(new_n225), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n664), .B1(new_n636), .B2(new_n642), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n622), .B(KEYINPUT88), .Z(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT26), .B1(new_n408), .B2(new_n638), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n696), .C1(new_n641), .C2(KEYINPUT26), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n618), .A2(new_n625), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n627), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n664), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT94), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n330), .A2(new_n331), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n452), .B1(new_n705), .B2(new_n268), .ZN(new_n706));
  AOI21_X1  g0506(.A(G179), .B1(new_n263), .B2(new_n282), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT93), .B1(new_n707), .B2(new_n394), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT93), .ZN(new_n709));
  NOR4_X1   g0509(.A1(new_n311), .A2(new_n709), .A3(G179), .A4(new_n387), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n706), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n330), .A2(new_n331), .A3(new_n387), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(KEYINPUT92), .A2(KEYINPUT30), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n306), .A3(new_n452), .A4(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n452), .A2(G179), .A3(new_n263), .A4(new_n282), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n716), .A2(new_n712), .B1(KEYINPUT92), .B2(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n704), .A2(new_n719), .A3(KEYINPUT31), .A4(new_n664), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n711), .B2(new_n718), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n704), .B1(new_n722), .B2(new_n664), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n355), .A2(new_n408), .A3(new_n396), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(new_n633), .A3(new_n459), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n726), .B2(new_n320), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n664), .B1(new_n719), .B2(KEYINPUT31), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n724), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n703), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n691), .B1(new_n733), .B2(G1), .ZN(G364));
  OR3_X1    g0534(.A1(KEYINPUT95), .A2(G13), .A3(G33), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT95), .B1(G13), .B2(G33), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n671), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n453), .A2(G20), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n388), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n388), .A2(new_n310), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G317), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT33), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n751), .A2(KEYINPUT33), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n743), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G329), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n742), .A2(G179), .A3(new_n310), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n754), .B(new_n758), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n226), .B1(new_n755), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n747), .B(new_n762), .C1(G294), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n226), .A2(new_n453), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n744), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G322), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n310), .A2(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G303), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n766), .A2(new_n748), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n272), .B1(new_n775), .B2(G326), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n765), .A2(new_n769), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n272), .B1(new_n205), .B2(new_n771), .C1(new_n761), .C2(new_n345), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n768), .A2(G58), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n749), .A2(new_n213), .B1(new_n745), .B2(new_n215), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G50), .B2(new_n775), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n764), .A2(G97), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n757), .A2(G159), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n777), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n227), .B1(G20), .B2(new_n301), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n272), .A2(G355), .A3(new_n220), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n241), .A2(new_n254), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n685), .A2(new_n272), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n225), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n790), .B1(G116), .B2(new_n220), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n739), .A2(new_n788), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n284), .A2(G20), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n688), .B1(G45), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n741), .A2(new_n789), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n671), .B2(G330), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G330), .B2(new_n671), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n559), .A2(new_n664), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n565), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n604), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n604), .A2(new_n664), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n737), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n737), .A2(new_n788), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n215), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n783), .B1(new_n345), .B2(new_n771), .C1(new_n812), .C2(new_n774), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n761), .A2(new_n205), .B1(new_n756), .B2(new_n746), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n277), .B1(new_n745), .B2(new_n286), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n759), .B2(new_n749), .C1(new_n817), .C2(new_n767), .ZN(new_n818));
  INV_X1    g0618(.A(new_n745), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G159), .B1(new_n768), .B2(G143), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n774), .C1(new_n470), .C2(new_n749), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n822), .A2(new_n823), .B1(G58), .B2(new_n764), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n772), .A2(G50), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n761), .A2(new_n213), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n272), .B1(new_n756), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT97), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n818), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n788), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n809), .A2(new_n798), .A3(new_n811), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n649), .B1(new_n565), .B2(new_n803), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n806), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n692), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(new_n731), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n839), .B2(new_n798), .ZN(G384));
  NOR2_X1   g0640(.A1(new_n598), .A2(new_n664), .ZN(new_n841));
  INV_X1    g0641(.A(new_n662), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n519), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n536), .A2(new_n537), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n611), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n545), .A2(new_n662), .B1(new_n541), .B2(new_n543), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n519), .A2(new_n533), .A3(new_n529), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n545), .A2(new_n542), .A3(new_n540), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n534), .A4(new_n843), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n846), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT39), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  AOI221_X4 g0658(.A(new_n858), .B1(new_n849), .B2(new_n852), .C1(new_n547), .C2(new_n844), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n611), .B1(new_n646), .B2(new_n647), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(KEYINPUT99), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT99), .B1(new_n849), .B2(new_n852), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n860), .A2(new_n843), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n859), .B1(new_n864), .B2(new_n858), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n841), .B(new_n857), .C1(new_n865), .C2(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n643), .A2(new_n665), .A3(new_n837), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n806), .B(KEYINPUT98), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n855), .A2(new_n856), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n576), .A2(new_n664), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n598), .A2(new_n601), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n598), .B2(new_n601), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n648), .A2(new_n842), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n866), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n616), .B1(new_n694), .B2(new_n702), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n653), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n879), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n837), .B1(new_n872), .B2(new_n873), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n725), .A2(new_n633), .A3(new_n459), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT31), .B1(new_n655), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n728), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n722), .A2(new_n664), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT99), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n853), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n861), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n536), .A2(KEYINPUT89), .A3(new_n537), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT89), .B1(new_n536), .B2(new_n537), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n612), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n844), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n888), .B(KEYINPUT40), .C1(new_n896), .C2(new_n859), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n598), .A2(new_n601), .A3(new_n871), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n598), .A2(new_n601), .ZN(new_n900));
  INV_X1    g0700(.A(new_n871), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n808), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n729), .B1(new_n460), .B2(KEYINPUT31), .ZN(new_n904));
  INV_X1    g0704(.A(new_n887), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n859), .A2(new_n854), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n898), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n886), .A2(new_n887), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n616), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(G330), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n882), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n265), .B2(new_n797), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n226), .B(new_n227), .C1(new_n350), .C2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(G116), .C1(new_n916), .C2(new_n350), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  OAI21_X1  g0719(.A(G77), .B1(new_n223), .B2(new_n213), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n225), .A2(new_n920), .B1(G50), .B2(new_n213), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n284), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(G367));
  NAND2_X1  g0723(.A1(new_n797), .A2(G45), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G1), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT104), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n640), .A2(new_n406), .A3(new_n664), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n406), .A2(new_n664), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n355), .A2(new_n408), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n683), .A2(KEYINPUT44), .A3(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n675), .B(new_n930), .C1(new_n674), .C2(new_n681), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT45), .Z(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT44), .B1(new_n683), .B2(new_n930), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(new_n680), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n677), .A2(new_n682), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n671), .A2(G330), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n671), .B2(G330), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT103), .B1(new_n678), .B2(new_n681), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n938), .B2(new_n939), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n732), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n686), .B(KEYINPUT41), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n926), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n677), .A2(new_n682), .A3(new_n930), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n408), .B1(new_n459), .B2(new_n929), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n665), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT101), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n949), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n950), .B(new_n952), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n379), .A2(new_n385), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n664), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n624), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n695), .B2(new_n959), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT100), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT102), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n957), .A2(new_n963), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n957), .A2(KEYINPUT102), .A3(new_n963), .A4(new_n964), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n679), .A2(new_n930), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n971), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n967), .A2(new_n973), .A3(new_n968), .A4(new_n969), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n948), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n961), .A2(new_n740), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n277), .B1(new_n763), .B2(new_n345), .ZN(new_n977));
  INV_X1    g0777(.A(new_n273), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n978), .A2(new_n767), .B1(new_n756), .B2(new_n751), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(G97), .C2(new_n760), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n775), .A2(G311), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n772), .A2(G116), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT46), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n819), .A2(G283), .B1(new_n750), .B2(G294), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n980), .A2(new_n981), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n756), .A2(new_n821), .B1(new_n771), .B2(new_n223), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n277), .B(new_n986), .C1(G159), .C2(new_n750), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n775), .A2(G143), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n819), .A2(G50), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n767), .A2(new_n470), .B1(new_n763), .B2(new_n213), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT106), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n761), .A2(new_n215), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n788), .ZN(new_n996));
  INV_X1    g0796(.A(new_n792), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n795), .B1(new_n220), .B2(new_n378), .C1(new_n237), .C2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT105), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n976), .A2(new_n996), .A3(new_n798), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n975), .A2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n926), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n944), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n772), .A2(G77), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n378), .B2(new_n763), .C1(new_n474), .C2(new_n767), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n757), .A2(G150), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n761), .A2(new_n207), .B1(new_n213), .B2(new_n745), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n517), .B2(new_n750), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n277), .B1(new_n775), .B2(G159), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n978), .A2(new_n745), .B1(new_n751), .B2(new_n767), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT108), .Z(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT109), .B(G322), .Z(new_n1014));
  OAI22_X1  g0814(.A1(new_n774), .A2(new_n1014), .B1(new_n749), .B2(new_n746), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n759), .B2(new_n763), .C1(new_n817), .C2(new_n771), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n760), .A2(G116), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n757), .A2(G326), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n277), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1011), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n788), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n678), .A2(new_n739), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n234), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n792), .B1(new_n1029), .B2(new_n254), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n272), .A2(new_n689), .A3(new_n220), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n213), .A2(new_n215), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n689), .A2(G45), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n471), .A2(G50), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT107), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT50), .Z(new_n1036));
  AOI22_X1  g0836(.A1(new_n1030), .A2(new_n1031), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n220), .A2(G107), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n795), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1027), .A2(new_n1028), .A3(new_n798), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n686), .B1(new_n944), .B2(new_n733), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n732), .B1(new_n942), .B2(new_n943), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1003), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(G393));
  INV_X1    g0843(.A(new_n1042), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT113), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n935), .B(new_n679), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT113), .B1(new_n936), .B2(new_n1042), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n936), .A2(new_n1042), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n686), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n936), .A2(new_n1002), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n761), .A2(new_n345), .B1(new_n756), .B2(new_n1014), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n774), .A2(new_n751), .B1(new_n767), .B2(new_n746), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT111), .Z(new_n1054));
  AOI211_X1 g0854(.A(new_n272), .B(new_n1052), .C1(new_n1054), .C2(KEYINPUT52), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n819), .A2(G294), .B1(G116), .B2(new_n764), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n978), .B2(new_n749), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT112), .Z(new_n1058));
  AND2_X1   g0858(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(KEYINPUT52), .B2(new_n1054), .C1(new_n759), .C2(new_n771), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n763), .A2(new_n215), .ZN(new_n1061));
  INV_X1    g0861(.A(G159), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n774), .A2(new_n470), .B1(new_n767), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n757), .A2(G143), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n277), .B1(new_n760), .B2(G87), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n745), .A2(new_n471), .B1(new_n771), .B2(new_n213), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G50), .B2(new_n750), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1060), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n788), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n927), .A2(new_n929), .A3(new_n739), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n795), .B1(new_n207), .B2(new_n220), .C1(new_n244), .C2(new_n997), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1071), .A2(new_n798), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1050), .A2(new_n1051), .A3(new_n1074), .ZN(G390));
  NAND4_X1  g0875(.A1(new_n730), .A2(G330), .A3(new_n837), .A4(new_n875), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n861), .A2(new_n890), .B1(new_n894), .B2(new_n844), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n856), .B1(new_n1078), .B2(KEYINPUT38), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n699), .A2(new_n664), .A3(new_n836), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n875), .B1(new_n1080), .B2(new_n806), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n841), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT39), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n859), .A2(new_n854), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n841), .B1(new_n869), .B2(new_n875), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1077), .B(new_n1083), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n857), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n868), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n692), .B2(new_n837), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1082), .B1(new_n1091), .B2(new_n874), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n865), .A2(new_n841), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1089), .A2(new_n1092), .B1(new_n1093), .B2(new_n1081), .ZN(new_n1094));
  INV_X1    g0894(.A(G330), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1095), .B(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1002), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT115), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1089), .A2(new_n737), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n810), .A2(new_n471), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n749), .A2(new_n345), .B1(new_n745), .B2(new_n207), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT116), .Z(new_n1104));
  NAND2_X1  g0904(.A1(new_n757), .A2(G294), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n277), .B1(new_n771), .B2(new_n205), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT117), .Z(new_n1107));
  NAND2_X1  g0907(.A1(new_n775), .A2(G283), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n767), .A2(new_n286), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1109), .A2(new_n827), .A3(new_n1061), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n764), .A2(G159), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n768), .A2(G132), .B1(new_n760), .B2(G50), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1113), .B1(new_n821), .B2(new_n749), .C1(new_n745), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n772), .A2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n277), .B1(new_n757), .B2(G125), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n774), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1116), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1111), .B1(new_n1112), .B2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT118), .Z(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n788), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1101), .A2(new_n798), .A3(new_n1102), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1100), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n616), .A2(G330), .A3(new_n910), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n880), .A2(new_n653), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1080), .A2(new_n806), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1076), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(G330), .B(new_n837), .C1(new_n904), .C2(new_n905), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n874), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT114), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT114), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1135), .A3(new_n874), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1095), .B1(new_n886), .B2(new_n724), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n875), .B1(new_n1138), .B2(new_n837), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n869), .B1(new_n1139), .B2(new_n1096), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1129), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1097), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1097), .A2(new_n1141), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1142), .A2(new_n686), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1127), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(G378));
  INV_X1    g0946(.A(new_n1129), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n476), .A2(new_n842), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n610), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n610), .A2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n502), .A2(new_n1150), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n610), .A2(new_n1151), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1155), .A2(new_n476), .A3(new_n842), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1095), .B1(new_n1158), .B2(KEYINPUT122), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n897), .A2(new_n908), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT122), .B1(new_n1158), .B2(KEYINPUT121), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1161), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(new_n897), .A3(new_n908), .A4(new_n1159), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1162), .A2(new_n879), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n877), .B1(new_n1086), .B2(new_n841), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1162), .A2(new_n1164), .B1(new_n1166), .B2(new_n876), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1148), .A2(new_n1168), .A3(KEYINPUT57), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT123), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1148), .A2(new_n1168), .A3(KEYINPUT123), .A4(KEYINPUT57), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n686), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT124), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT124), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1175), .A3(new_n686), .A4(new_n1172), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT57), .B1(new_n1148), .B2(new_n1168), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT125), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n767), .A2(new_n345), .B1(new_n763), .B2(new_n213), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G41), .B(new_n272), .C1(new_n760), .C2(G58), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n1004), .C1(new_n759), .C2(new_n756), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT119), .Z(new_n1183));
  AOI211_X1 g0983(.A(new_n1180), .B(new_n1183), .C1(G97), .C2(new_n750), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n286), .B2(new_n774), .C1(new_n378), .C2(new_n745), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT58), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n474), .B1(new_n275), .B2(G41), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n745), .A2(new_n821), .B1(new_n767), .B2(new_n1120), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1115), .A2(new_n771), .B1(new_n470), .B2(new_n763), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G125), .C2(new_n775), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n830), .B2(new_n749), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT59), .Z(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n757), .C2(G124), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n1062), .C2(new_n761), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1186), .A2(new_n1187), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(new_n788), .B1(new_n474), .B2(new_n810), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1158), .A2(new_n737), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n798), .A3(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT120), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1168), .B2(new_n1002), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1179), .A2(new_n1200), .ZN(G375));
  NOR2_X1   g1001(.A1(new_n767), .A2(new_n821), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n761), .A2(new_n223), .B1(new_n830), .B2(new_n774), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G50), .C2(new_n764), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n272), .B1(new_n745), .B2(new_n470), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G159), .B2(new_n772), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n1120), .C2(new_n756), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n750), .B2(new_n1114), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n756), .A2(new_n812), .B1(new_n378), .B2(new_n763), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n761), .A2(new_n215), .B1(new_n207), .B2(new_n771), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G294), .C2(new_n775), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n272), .B1(new_n819), .B2(G107), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n759), .C2(new_n767), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G116), .B2(new_n750), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n788), .B1(new_n1208), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n798), .B(new_n1215), .C1(new_n875), .C2(new_n738), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n213), .B2(new_n810), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n1002), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1137), .A2(new_n1140), .A3(new_n1129), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n946), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1221), .B2(new_n1141), .ZN(G381));
  NAND3_X1  g1022(.A1(new_n1179), .A2(new_n1145), .A3(new_n1200), .ZN(new_n1223));
  OR2_X1    g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1223), .A2(G387), .A3(G390), .A4(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G381), .A2(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(G407));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  NAND4_X1  g1028(.A1(G387), .A2(new_n1051), .A3(new_n1050), .A4(new_n1074), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(G390), .A2(new_n975), .A3(new_n1000), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(G393), .B(G396), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT127), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1229), .A2(new_n1233), .A3(new_n1230), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1145), .B1(new_n1179), .B2(new_n1200), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n686), .B1(new_n1220), .B2(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(new_n1141), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1220), .A2(new_n1241), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1219), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(G384), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n659), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1148), .A2(new_n1168), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(new_n947), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1249), .A2(new_n1252), .A3(new_n947), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1145), .B(new_n1200), .C1(new_n1251), .C2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(new_n1240), .A2(new_n1247), .A3(new_n1248), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT62), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1240), .A2(new_n1248), .A3(new_n1255), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1248), .A2(G2897), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1246), .B(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1256), .A2(new_n1257), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1248), .B1(G375), .B2(G378), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1262), .A2(new_n1257), .A3(new_n1246), .A4(new_n1254), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1239), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1237), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1230), .A2(new_n1229), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1264), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1256), .B2(KEYINPUT63), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1262), .A2(new_n1254), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1260), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1270), .B1(new_n1274), .B2(new_n1256), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1275), .ZN(G405));
  INV_X1    g1076(.A(new_n1240), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1223), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1239), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1238), .A2(new_n1223), .A3(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1247), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1246), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(G402));
endmodule


