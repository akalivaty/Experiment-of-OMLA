//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n187), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n196), .A2(new_n198), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT19), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g025(.A(G125), .B(G140), .Z(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT72), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT72), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI211_X1 g030(.A(G146), .B(new_n211), .C1(new_n216), .C2(new_n210), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT18), .A2(G131), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT86), .B1(new_n194), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT86), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n193), .A2(new_n220), .A3(KEYINPUT18), .A4(G131), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n194), .A2(new_n218), .ZN(new_n223));
  AOI21_X1  g037(.A(G146), .B1(new_n213), .B2(new_n215), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n206), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n209), .A2(new_n217), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n200), .A2(new_n234), .A3(new_n202), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n193), .A2(KEYINPUT17), .A3(new_n201), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n236), .A2(KEYINPUT87), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n207), .B(new_n225), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(KEYINPUT87), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n216), .A2(new_n225), .ZN(new_n241));
  INV_X1    g055(.A(new_n226), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n223), .A3(new_n219), .A4(new_n221), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n244), .A3(new_n231), .ZN(new_n245));
  AOI21_X1  g059(.A(G475), .B1(new_n233), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n247));
  INV_X1    g061(.A(G902), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT88), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n246), .A2(new_n248), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT88), .A3(new_n247), .ZN(new_n254));
  INV_X1    g068(.A(new_n245), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n231), .B1(new_n240), .B2(new_n244), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n248), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n252), .A2(new_n254), .B1(G475), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(G234), .A2(G237), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(G952), .A3(new_n188), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT21), .B(G898), .Z(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(G902), .A3(G953), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G116), .B(G122), .ZN(new_n264));
  INV_X1    g078(.A(G107), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT14), .A3(G122), .ZN(new_n268));
  XOR2_X1   g082(.A(G116), .B(G122), .Z(new_n269));
  OAI211_X1 g083(.A(G107), .B(new_n268), .C1(new_n269), .C2(KEYINPUT14), .ZN(new_n270));
  INV_X1    g084(.A(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT89), .B1(new_n271), .B2(G143), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n190), .A3(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(G143), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n266), .B(new_n270), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(KEYINPUT9), .A2(G234), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT9), .A2(G234), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT75), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n285), .A2(G217), .A3(new_n188), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT13), .B1(new_n272), .B2(new_n274), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT13), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(new_n277), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n276), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n269), .A2(G107), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n266), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n278), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n281), .B(new_n289), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT13), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n275), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n291), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n290), .A2(KEYINPUT90), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n298), .B1(new_n304), .B2(G134), .ZN(new_n305));
  INV_X1    g119(.A(new_n281), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n288), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n248), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n309), .B(new_n311), .Z(new_n312));
  NAND3_X1  g126(.A1(new_n258), .A2(new_n263), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  XOR2_X1   g128(.A(G110), .B(G122), .Z(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT8), .Z(new_n316));
  NOR2_X1   g130(.A1(new_n230), .A2(G107), .ZN(new_n317));
  AND2_X1   g131(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n318));
  NOR2_X1   g132(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n317), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n265), .A2(G104), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n317), .B(KEYINPUT77), .C1(new_n319), .C2(new_n318), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n322), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n329));
  OAI21_X1  g143(.A(G101), .B1(new_n317), .B2(new_n324), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n328), .B2(new_n330), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G116), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(KEYINPUT83), .ZN(new_n336));
  XNOR2_X1  g150(.A(G116), .B(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT5), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(KEYINPUT83), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n336), .A2(new_n338), .A3(G113), .A4(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT2), .B(G113), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n331), .A2(new_n332), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n328), .A2(new_n330), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n316), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n225), .A2(G143), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT65), .B1(new_n190), .B2(G146), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n225), .A3(G143), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT0), .A2(G128), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n190), .A2(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n225), .A2(G143), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT0), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n271), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n352), .A2(new_n353), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n204), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n354), .A2(new_n355), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n271), .B1(new_n355), .B2(KEYINPUT1), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n350), .B1(G143), .B2(new_n225), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n190), .A2(KEYINPUT65), .A3(G146), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n367), .B(new_n354), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n352), .A2(new_n372), .A3(new_n367), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n366), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n363), .B1(new_n374), .B2(new_n204), .ZN(new_n375));
  INV_X1    g189(.A(G224), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G953), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n378), .A2(KEYINPUT7), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(KEYINPUT84), .ZN(new_n380));
  OR3_X1    g194(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n322), .A2(new_n325), .A3(new_n327), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n328), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n385), .A3(G101), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT2), .B(G113), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n267), .A2(G119), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n334), .A2(G116), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n342), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n345), .A2(KEYINPUT79), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n394));
  INV_X1    g208(.A(new_n343), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n315), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n379), .B1(new_n375), .B2(new_n380), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n347), .A2(new_n381), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n248), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n396), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n315), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n375), .B(new_n378), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n407), .A3(new_n315), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT85), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n402), .B2(new_n409), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n314), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n313), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n285), .A2(new_n287), .ZN(new_n418));
  OAI21_X1  g232(.A(G221), .B1(new_n418), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n331), .A2(new_n332), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n374), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n372), .B1(new_n352), .B2(new_n367), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n425), .A2(new_n426), .B1(new_n352), .B2(new_n365), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n328), .A3(new_n330), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n422), .A2(new_n424), .B1(new_n428), .B2(new_n423), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT11), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n276), .B2(G137), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n276), .A2(G137), .ZN(new_n432));
  INV_X1    g246(.A(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT11), .A3(G134), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G131), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n199), .A2(new_n432), .A3(new_n434), .A4(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n328), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n386), .A2(new_n362), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n384), .A2(KEYINPUT78), .A3(new_n386), .A4(new_n362), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n429), .A2(new_n439), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G140), .ZN(new_n446));
  INV_X1    g260(.A(G227), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n446), .B(new_n448), .Z(new_n449));
  AND3_X1   g263(.A1(new_n445), .A2(KEYINPUT80), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n428), .A2(new_n423), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n424), .A2(new_n393), .A3(new_n394), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n443), .A2(new_n451), .A3(new_n452), .A4(new_n444), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT81), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n429), .A2(new_n455), .A3(new_n443), .A4(new_n444), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n439), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT80), .B1(new_n445), .B2(new_n449), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n450), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n366), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n425), .B2(new_n426), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n428), .B1(new_n422), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n438), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT12), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n462), .B2(new_n438), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n445), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n449), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n421), .B1(new_n459), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n456), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n438), .ZN(new_n472));
  INV_X1    g286(.A(new_n458), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n445), .A2(KEYINPUT80), .A3(new_n449), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n467), .A2(new_n468), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(KEYINPUT82), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n420), .B1(new_n470), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n445), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n468), .B1(new_n457), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n445), .B(new_n449), .C1(new_n465), .C2(new_n466), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n420), .A3(new_n248), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n420), .A2(new_n248), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n417), .B(new_n419), .C1(new_n478), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n475), .A2(KEYINPUT82), .A3(new_n476), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT82), .B1(new_n475), .B2(new_n476), .ZN(new_n491));
  OAI21_X1  g305(.A(G469), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n480), .B2(new_n481), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n484), .B1(new_n493), .B2(new_n420), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n419), .A4(new_n417), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT22), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n433), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(G119), .B(G128), .Z(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT71), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n271), .A2(G119), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT23), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(G119), .B2(new_n271), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n241), .B(new_n208), .C1(new_n504), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n238), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n502), .A2(new_n503), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(G110), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT73), .B1(new_n509), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n500), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n499), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT25), .B1(new_n520), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(G217), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(G234), .B2(new_n248), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n518), .A2(new_n524), .A3(new_n519), .A4(new_n248), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n523), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n518), .A2(new_n529), .A3(new_n519), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(G101), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n435), .A2(new_n201), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n433), .A2(G134), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n195), .B1(new_n432), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n461), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n391), .B1(new_n438), .B2(new_n362), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT68), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n537), .A2(new_n539), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(KEYINPUT68), .C1(new_n374), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n536), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT69), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n438), .A2(new_n362), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n541), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n549), .B1(new_n541), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n391), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n374), .A2(new_n544), .ZN(new_n556));
  INV_X1    g370(.A(new_n542), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n545), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n536), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT31), .ZN(new_n563));
  INV_X1    g377(.A(new_n536), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n541), .A2(new_n550), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n391), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n565), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT28), .B1(new_n541), .B2(new_n542), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n548), .A2(new_n571), .A3(new_n561), .A4(new_n554), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n563), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT70), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n563), .A2(new_n575), .A3(new_n570), .A4(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n582));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n554), .A2(new_n559), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT29), .B1(new_n584), .B2(new_n564), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n568), .A2(new_n569), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n536), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(KEYINPUT29), .A3(new_n536), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n581), .A2(new_n582), .A3(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n489), .A2(new_n496), .A3(new_n532), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  OAI21_X1  g408(.A(new_n419), .B1(new_n478), .B2(new_n486), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n583), .A2(KEYINPUT92), .ZN(new_n596));
  AOI211_X1 g410(.A(G902), .B(new_n596), .C1(new_n574), .C2(new_n576), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n574), .B2(new_n576), .ZN(new_n598));
  INV_X1    g412(.A(new_n596), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n595), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n601), .A2(new_n532), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT97), .B(G478), .Z(new_n603));
  NAND2_X1  g417(.A1(new_n309), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n288), .B(KEYINPUT94), .ZN(new_n607));
  OAI211_X1 g421(.A(KEYINPUT95), .B(new_n607), .C1(new_n305), .C2(new_n306), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(new_n299), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n305), .B2(new_n306), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n606), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n299), .A2(new_n307), .A3(new_n606), .ZN(new_n614));
  OAI211_X1 g428(.A(G478), .B(new_n248), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n610), .A2(new_n611), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n299), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n614), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n310), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(KEYINPUT96), .A3(new_n248), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n605), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT98), .B1(new_n624), .B2(new_n258), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT96), .B1(new_n622), .B2(new_n248), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n612), .A2(new_n299), .A3(new_n608), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n614), .B1(new_n627), .B2(KEYINPUT33), .ZN(new_n628));
  NOR4_X1   g442(.A1(new_n628), .A2(new_n616), .A3(new_n310), .A4(G902), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n604), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n252), .A2(new_n254), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n257), .A2(G475), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n625), .A2(new_n635), .A3(new_n263), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n411), .B1(new_n637), .B2(new_n401), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(KEYINPUT93), .A3(new_n413), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT93), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n415), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n639), .A2(new_n314), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n602), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n230), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(G6));
  XNOR2_X1  g460(.A(new_n253), .B(new_n247), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n632), .ZN(new_n648));
  INV_X1    g462(.A(new_n263), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n648), .A2(new_n649), .A3(new_n312), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n602), .A2(new_n642), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n600), .A2(new_n597), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n514), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n528), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT100), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n526), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n489), .A2(new_n496), .A3(new_n654), .A4(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT37), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G110), .ZN(G12));
  OAI211_X1 g476(.A(new_n419), .B(new_n659), .C1(new_n478), .C2(new_n486), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n260), .B(KEYINPUT101), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(G900), .B2(new_n262), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n648), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n312), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n664), .A2(new_n592), .A3(new_n642), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  INV_X1    g488(.A(new_n419), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n492), .B2(new_n494), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n667), .B(KEYINPUT102), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT40), .Z(new_n680));
  INV_X1    g494(.A(new_n562), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n536), .B1(new_n559), .B2(new_n567), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n248), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G472), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n581), .A2(new_n582), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n659), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n414), .A2(new_n415), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT38), .Z(new_n689));
  NOR2_X1   g503(.A1(new_n258), .A2(new_n312), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n680), .A2(new_n314), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  NAND3_X1  g507(.A1(new_n630), .A2(new_n633), .A3(new_n667), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n639), .A2(new_n314), .A3(new_n641), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n694), .B2(new_n695), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n664), .A2(new_n592), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  AOI21_X1  g515(.A(new_n420), .B1(new_n482), .B2(new_n248), .ZN(new_n702));
  AOI211_X1 g516(.A(G469), .B(G902), .C1(new_n480), .C2(new_n481), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n695), .A2(new_n702), .A3(new_n703), .A4(new_n675), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n592), .A2(new_n532), .A3(new_n704), .A4(new_n636), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT104), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n592), .A2(new_n532), .A3(new_n704), .A4(new_n650), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  INV_X1    g524(.A(new_n659), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n313), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n592), .A2(new_n704), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NAND2_X1  g528(.A1(new_n573), .A2(new_n578), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n532), .B(new_n715), .C1(new_n598), .C2(new_n583), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n704), .A3(new_n263), .A4(new_n690), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  OAI211_X1 g533(.A(new_n659), .B(new_n715), .C1(new_n598), .C2(new_n583), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n694), .A2(new_n695), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n702), .A2(new_n703), .A3(new_n675), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n702), .A2(new_n703), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n624), .A2(new_n258), .A3(new_n668), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n642), .A3(new_n727), .A4(new_n419), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT105), .B1(new_n728), .B2(new_n720), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  NOR2_X1   g545(.A1(new_n459), .A2(KEYINPUT106), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n475), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(G469), .B(new_n476), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n675), .B1(new_n735), .B2(new_n494), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n688), .A2(new_n314), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n694), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n592), .A2(new_n532), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT107), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n735), .A2(new_n494), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(new_n419), .A3(new_n738), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n532), .A4(new_n592), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n740), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT32), .B1(new_n577), .B2(new_n578), .ZN(new_n748));
  INV_X1    g562(.A(new_n578), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n580), .B(new_n749), .C1(new_n574), .C2(new_n576), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n748), .A2(new_n750), .A3(new_n590), .ZN(new_n751));
  INV_X1    g565(.A(new_n532), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n592), .A2(KEYINPUT108), .A3(new_n532), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(KEYINPUT42), .A3(new_n743), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  AND2_X1   g571(.A1(new_n736), .A2(new_n672), .ZN(new_n758));
  INV_X1    g572(.A(new_n737), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n592), .A3(new_n532), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  OAI211_X1 g575(.A(KEYINPUT45), .B(new_n476), .C1(new_n732), .C2(new_n734), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n470), .A2(new_n477), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n762), .B(G469), .C1(KEYINPUT45), .C2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n485), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n483), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n773));
  NOR2_X1   g587(.A1(new_n624), .A2(new_n633), .ZN(new_n774));
  MUX2_X1   g588(.A(new_n772), .B(new_n773), .S(new_n774), .Z(new_n775));
  INV_X1    g589(.A(new_n654), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n659), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n770), .A2(new_n419), .A3(new_n678), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n759), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  AND3_X1   g599(.A1(new_n751), .A2(new_n752), .A3(new_n738), .ZN(new_n786));
  INV_X1    g600(.A(new_n769), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n419), .B1(new_n767), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(G952), .A2(G953), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT120), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n775), .A2(new_n665), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n775), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n717), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n689), .A2(new_n314), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n724), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT50), .B1(new_n806), .B2(KEYINPUT117), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(KEYINPUT117), .B2(KEYINPUT50), .ZN(new_n808));
  INV_X1    g622(.A(new_n724), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n810), .B2(new_n805), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n737), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n801), .A2(new_n721), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT118), .ZN(new_n814));
  INV_X1    g628(.A(new_n812), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n815), .A2(new_n260), .A3(new_n752), .A4(new_n685), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n258), .A3(new_n624), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n807), .A2(new_n811), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n802), .A2(new_n737), .ZN(new_n820));
  INV_X1    g634(.A(new_n792), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n790), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n726), .A2(new_n675), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT115), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n790), .A3(new_n823), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(new_n820), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n826), .A2(new_n827), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n751), .A2(new_n663), .A3(new_n697), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n832), .A2(new_n699), .B1(new_n725), .B2(new_n729), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n675), .B(new_n668), .C1(new_n735), .C2(new_n494), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n695), .A2(new_n312), .A3(new_n258), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n685), .A3(new_n711), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(KEYINPUT112), .A3(new_n673), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n730), .A2(new_n673), .A3(new_n700), .A4(new_n836), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n838), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  MUX2_X1   g658(.A(new_n630), .B(new_n670), .S(new_n258), .Z(new_n845));
  NOR2_X1   g659(.A1(new_n416), .A2(new_n649), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n601), .A2(new_n532), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n593), .A3(new_n660), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n705), .A2(new_n709), .A3(new_n718), .A4(new_n713), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n664), .A2(new_n312), .A3(new_n592), .A4(new_n669), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n737), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n743), .A2(new_n721), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n760), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n746), .B2(new_n755), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n852), .B2(new_n856), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n831), .B(new_n844), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n855), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n756), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n489), .A2(new_n496), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n751), .A2(new_n752), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n676), .A2(new_n654), .A3(new_n532), .A4(new_n846), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n862), .A2(new_n863), .B1(new_n864), .B2(new_n845), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n705), .A2(new_n709), .A3(new_n713), .A4(new_n718), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n850), .A2(new_n737), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n660), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT111), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n838), .A2(new_n839), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n838), .A2(new_n839), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT52), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n842), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n859), .B(KEYINPUT54), .C1(new_n874), .C2(new_n831), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n844), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n856), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n876), .B(new_n877), .C1(new_n874), .C2(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT113), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n803), .A2(new_n704), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n625), .A2(new_n635), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n816), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(G952), .A3(new_n188), .A4(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT119), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n830), .A2(new_n880), .A3(new_n882), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n753), .A2(new_n754), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n801), .A2(new_n890), .A3(new_n812), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT48), .Z(new_n892));
  OAI21_X1  g706(.A(new_n796), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n726), .B(KEYINPUT49), .Z(new_n894));
  NOR4_X1   g708(.A1(new_n894), .A2(new_n675), .A3(new_n752), .A4(new_n689), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n314), .A3(new_n686), .A4(new_n774), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(G75));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n877), .B1(new_n874), .B2(KEYINPUT53), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(G902), .A3(new_n411), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT121), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n405), .A2(new_n408), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n406), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n637), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND4_X1   g719(.A1(new_n898), .A2(new_n901), .A3(new_n900), .A4(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n188), .A2(G952), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n901), .A2(new_n905), .B1(new_n898), .B2(new_n900), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n878), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n484), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n485), .A2(KEYINPUT57), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n482), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n899), .A2(G902), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(new_n764), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n907), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND4_X1  g732(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n233), .A2(new_n245), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n907), .ZN(G60));
  INV_X1    g737(.A(new_n628), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n911), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n907), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n880), .B2(new_n882), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT122), .B1(new_n931), .B2(new_n924), .ZN(new_n932));
  INV_X1    g746(.A(new_n882), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n881), .B1(new_n875), .B2(new_n878), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n936), .A3(new_n628), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n930), .B1(new_n932), .B2(new_n937), .ZN(G63));
  XNOR2_X1  g752(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n899), .A2(new_n656), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n929), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n899), .A2(new_n942), .B1(new_n527), .B2(new_n530), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT125), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n899), .A2(new_n942), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n527), .A2(new_n530), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n950), .A3(new_n929), .A4(new_n943), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT61), .B1(new_n946), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  INV_X1    g768(.A(new_n261), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n955), .B2(new_n376), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n848), .A2(new_n849), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n902), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(G898), .B2(new_n188), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  NOR2_X1   g775(.A1(new_n552), .A2(new_n553), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n211), .B1(new_n216), .B2(new_n210), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G227), .A2(G953), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n833), .A2(new_n673), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n692), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT62), .Z(new_n968));
  INV_X1    g782(.A(new_n679), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n863), .A2(new_n969), .A3(new_n759), .A4(new_n845), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n784), .A3(new_n793), .A4(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n964), .B(new_n965), .C1(new_n971), .C2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(G900), .B1(new_n964), .B2(new_n447), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(G953), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n966), .B1(new_n780), .B2(new_n783), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(KEYINPUT126), .B(new_n966), .C1(new_n780), .C2(new_n783), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n793), .A2(new_n756), .A3(new_n760), .ZN(new_n980));
  INV_X1    g794(.A(new_n788), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(new_n678), .A3(new_n890), .A4(new_n835), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n979), .A2(new_n980), .A3(new_n188), .A4(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n972), .B(new_n974), .C1(new_n983), .C2(new_n964), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  INV_X1    g800(.A(new_n957), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n971), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n536), .A3(new_n584), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n681), .B1(new_n564), .B2(new_n584), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n859), .B(new_n986), .C1(new_n874), .C2(new_n831), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n989), .B(new_n929), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n979), .A2(new_n980), .A3(new_n957), .A4(new_n982), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n993), .A2(new_n994), .A3(new_n986), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n993), .B2(new_n986), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n536), .ZN(new_n997));
  INV_X1    g811(.A(new_n584), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n992), .B1(new_n997), .B2(new_n998), .ZN(G57));
endmodule


