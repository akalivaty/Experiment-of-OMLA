//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT0), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(G143), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n198), .A2(new_n192), .B1(KEYINPUT0), .B2(G128), .ZN(new_n199));
  OR3_X1    g013(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n194), .A2(new_n197), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT11), .B1(new_n205), .B2(G134), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(G137), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT11), .A2(G134), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n205), .B2(G134), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT67), .A3(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n204), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n205), .A2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(new_n208), .ZN(new_n219));
  INV_X1    g033(.A(new_n206), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n204), .A2(new_n214), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n203), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(KEYINPUT70), .A2(G116), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT70), .A2(G116), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(G119), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(KEYINPUT69), .A2(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT69), .A2(G119), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(G116), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT2), .B(G113), .Z(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n209), .A2(new_n204), .A3(new_n214), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n198), .A2(new_n192), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n189), .A2(new_n191), .A3(new_n237), .A4(new_n192), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n205), .A2(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n207), .B2(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n232), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n222), .A2(new_n231), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n222), .A2(KEYINPUT71), .A3(new_n231), .A4(new_n243), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT74), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n249), .A2(KEYINPUT74), .A3(new_n250), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n222), .A2(new_n243), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n255), .A2(new_n231), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n247), .B1(new_n257), .B2(KEYINPUT28), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT29), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n222), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n214), .A2(new_n219), .A3(new_n220), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n232), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n203), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n231), .B1(new_n276), .B2(new_n243), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT28), .B1(new_n277), .B2(new_n251), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n264), .B(KEYINPUT73), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n246), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n255), .A2(KEYINPUT30), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n229), .B(new_n230), .Z(new_n282));
  INV_X1    g096(.A(new_n243), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n271), .B2(new_n275), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n281), .B(new_n282), .C1(new_n284), .C2(KEYINPUT30), .ZN(new_n285));
  INV_X1    g099(.A(new_n251), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n265), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n280), .A2(new_n288), .A3(new_n266), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n268), .A2(new_n269), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n249), .A2(new_n250), .A3(new_n264), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n249), .A2(new_n295), .A3(new_n250), .A4(new_n264), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n285), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n294), .A2(new_n285), .A3(KEYINPUT31), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n279), .B1(new_n278), .B2(new_n246), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n292), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n307));
  INV_X1    g121(.A(new_n305), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(KEYINPUT32), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n291), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G140), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n260), .A2(G227), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n193), .A2(new_n234), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n238), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n316), .B2(G107), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n318));
  INV_X1    g132(.A(G107), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G104), .ZN(new_n320));
  INV_X1    g134(.A(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(G107), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n317), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n316), .A2(G107), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n319), .A2(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(G101), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n326), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n236), .A3(new_n238), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n274), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT12), .B1(new_n331), .B2(new_n274), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n202), .A2(new_n199), .ZN(new_n335));
  INV_X1    g149(.A(new_n197), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n193), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n317), .A2(new_n320), .A3(new_n322), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT82), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n317), .A2(new_n320), .A3(new_n340), .A4(new_n322), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(G101), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n321), .B1(new_n338), .B2(KEYINPUT82), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(new_n236), .B2(new_n238), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n327), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n329), .B1(new_n238), .B2(new_n314), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(KEYINPUT10), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n347), .A2(new_n352), .A3(new_n274), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n313), .B1(new_n334), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n345), .A2(new_n341), .B1(KEYINPUT4), .B2(new_n323), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n203), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n274), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n328), .A2(new_n348), .B1(new_n327), .B2(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n361));
  INV_X1    g175(.A(new_n313), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n274), .B1(new_n347), .B2(new_n352), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n361), .B1(new_n360), .B2(new_n362), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n354), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n354), .B(new_n369), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT85), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n370), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT83), .B1(new_n353), .B2(new_n313), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n363), .A3(new_n364), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n369), .B1(new_n376), .B2(new_n354), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n269), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G469), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n362), .B1(new_n364), .B2(new_n360), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT86), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n360), .B(new_n362), .C1(new_n332), .C2(new_n333), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n381), .A2(KEYINPUT86), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n372), .B(new_n269), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n385), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n382), .A3(new_n383), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n372), .A4(new_n269), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n373), .A2(new_n380), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n226), .A2(G128), .A3(new_n227), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT75), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n226), .A2(new_n227), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n196), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n401), .A3(KEYINPUT23), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(KEYINPUT76), .A3(new_n196), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n396), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G110), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT24), .B(G110), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n196), .A2(G119), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n394), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT16), .ZN(new_n411));
  INV_X1    g225(.A(G140), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(G125), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT80), .ZN(new_n414));
  INV_X1    g228(.A(G125), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT78), .B1(new_n415), .B2(KEYINPUT77), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n412), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT78), .B(G140), .C1(new_n415), .C2(KEYINPUT77), .ZN(new_n418));
  AND2_X1   g232(.A1(G125), .A2(G140), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n416), .A2(new_n412), .B1(new_n420), .B2(new_n419), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT16), .A4(new_n418), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n414), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G146), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n190), .B(new_n414), .C1(new_n423), .C2(new_n426), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n407), .B(new_n410), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G110), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n404), .A2(new_n431), .A3(new_n405), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n408), .B1(new_n409), .B2(new_n394), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n427), .A2(G146), .ZN(new_n437));
  NOR2_X1   g251(.A1(G125), .A2(G140), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n419), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G146), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT22), .B(G137), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n443), .B(new_n444), .Z(new_n445));
  AND3_X1   g259(.A1(new_n430), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n430), .B2(new_n442), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT25), .A3(new_n269), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n430), .A2(new_n442), .ZN(new_n450));
  INV_X1    g264(.A(new_n445), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n430), .A2(new_n442), .A3(new_n445), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n269), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(G234), .B2(new_n269), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G902), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n457), .A2(new_n459), .B1(new_n448), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT5), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT5), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n226), .A2(new_n464), .A3(G116), .A4(new_n227), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G113), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n462), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n230), .A2(new_n225), .A3(new_n228), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT5), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n469), .A2(KEYINPUT88), .A3(G113), .A4(new_n465), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n467), .A2(new_n468), .A3(new_n327), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT89), .ZN(new_n472));
  INV_X1    g286(.A(new_n468), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(G113), .A3(new_n465), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n462), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n327), .A4(new_n470), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n282), .B1(new_n356), .B2(new_n355), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n472), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n472), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n484));
  OR3_X1    g298(.A1(new_n203), .A2(KEYINPUT90), .A3(new_n415), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n236), .A2(new_n415), .A3(new_n238), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n337), .A2(G125), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n260), .A2(G224), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT92), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n495), .A3(new_n481), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n484), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n475), .A2(new_n329), .A3(new_n470), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n480), .B(KEYINPUT8), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n474), .A2(new_n468), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n498), .B(new_n499), .C1(new_n329), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n488), .A2(new_n489), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n492), .A2(KEYINPUT7), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n488), .A2(new_n485), .A3(new_n490), .A4(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n507), .B2(new_n483), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G210), .B1(G237), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT93), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n497), .A2(new_n512), .A3(new_n508), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(G104), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n188), .ZN(new_n520));
  AND2_X1   g334(.A1(KEYINPUT18), .A2(G131), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n424), .A2(new_n418), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n440), .B1(new_n523), .B2(G146), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n518), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n424), .A2(KEYINPUT19), .A3(new_n418), .ZN(new_n526));
  INV_X1    g340(.A(new_n439), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(KEYINPUT19), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n520), .A2(G131), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n519), .A2(new_n188), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n519), .A2(new_n188), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n204), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n528), .A2(new_n190), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n525), .B1(new_n533), .B2(new_n437), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n522), .A2(new_n524), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n428), .A2(new_n429), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n539), .A3(new_n532), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n520), .A2(KEYINPUT17), .A3(G131), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n537), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n535), .B(new_n536), .C1(new_n543), .C2(new_n518), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT20), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n423), .A2(new_n426), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n190), .B1(new_n546), .B2(new_n414), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(new_n542), .A3(new_n437), .ZN(new_n548));
  INV_X1    g362(.A(new_n537), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n518), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n534), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n536), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n518), .A2(KEYINPUT94), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n548), .A2(new_n557), .A3(new_n549), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n269), .A3(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n545), .A2(new_n554), .B1(G475), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G128), .B(G143), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(new_n212), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n223), .A2(G122), .A3(new_n224), .ZN(new_n563));
  INV_X1    g377(.A(G122), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G116), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n319), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT14), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n563), .A2(new_n567), .A3(new_n565), .ZN(new_n568));
  OAI21_X1  g382(.A(G107), .B1(new_n563), .B2(new_n567), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n562), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n561), .A2(KEYINPUT13), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n196), .A2(KEYINPUT13), .A3(G143), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n212), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n571), .A2(new_n573), .B1(new_n212), .B2(new_n561), .ZN(new_n574));
  INV_X1    g388(.A(new_n566), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n319), .B1(new_n563), .B2(new_n565), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT9), .B(G234), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n578), .A2(new_n458), .A3(G953), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n570), .B2(new_n577), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n269), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT95), .ZN(new_n583));
  INV_X1    g397(.A(G478), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT95), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n269), .C1(new_n580), .C2(new_n581), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n582), .A2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G234), .ZN(new_n592));
  OAI211_X1 g406(.A(G902), .B(G953), .C1(new_n592), .C2(new_n259), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT96), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT21), .B(G898), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n260), .A2(G952), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n592), .B2(new_n259), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G221), .B1(new_n578), .B2(G902), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G214), .B1(G237), .B2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n560), .A2(new_n591), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n516), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n310), .A2(new_n393), .A3(new_n461), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND2_X1  g422(.A1(new_n368), .A2(new_n370), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n372), .B1(new_n609), .B2(new_n269), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n610), .A2(new_n379), .B1(new_n388), .B2(new_n391), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n601), .B1(new_n611), .B2(new_n373), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n509), .A2(new_n511), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n497), .A2(new_n510), .A3(new_n508), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n603), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n304), .A2(new_n305), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n307), .B2(G902), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n461), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n623), .B(KEYINPUT33), .C1(new_n580), .C2(new_n581), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n570), .A2(new_n577), .ZN(new_n625));
  INV_X1    g439(.A(new_n579), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n627), .B(new_n621), .C1(new_n622), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n584), .A2(G902), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n620), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n631), .ZN(new_n633));
  AOI211_X1 g447(.A(KEYINPUT98), .B(new_n633), .C1(new_n624), .C2(new_n629), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n560), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n599), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NOR2_X1   g455(.A1(new_n543), .A2(new_n557), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n558), .A2(new_n269), .ZN(new_n643));
  OAI21_X1  g457(.A(G475), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n553), .B1(new_n552), .B2(new_n536), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n518), .B1(new_n548), .B2(new_n549), .ZN(new_n646));
  INV_X1    g460(.A(new_n536), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n646), .A2(KEYINPUT20), .A3(new_n534), .A4(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n644), .B(new_n590), .C1(new_n645), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n599), .B(KEYINPUT99), .Z(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n619), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT35), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT100), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  AND2_X1   g469(.A1(new_n616), .A2(new_n617), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT25), .B1(new_n448), .B2(new_n269), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n446), .A2(new_n447), .A3(new_n455), .A4(G902), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n459), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n451), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n450), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n460), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n393), .A2(new_n656), .A3(new_n606), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  NAND3_X1  g480(.A1(new_n304), .A2(new_n292), .A3(new_n305), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT32), .B1(new_n307), .B2(new_n308), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n667), .A2(new_n668), .B1(G472), .B2(new_n290), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n615), .A2(new_n663), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n594), .A2(KEYINPUT101), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n598), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT101), .B1(new_n594), .B2(new_n671), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT102), .B1(new_n649), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n677));
  INV_X1    g491(.A(new_n675), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n560), .A2(new_n677), .A3(new_n590), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n669), .A2(new_n670), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n612), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n675), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n612), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT104), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n514), .A2(new_n515), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT38), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n667), .A2(new_n668), .ZN(new_n692));
  INV_X1    g506(.A(new_n279), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n257), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n694), .A2(new_n297), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n560), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n590), .A3(new_n602), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n691), .A2(new_n698), .A3(new_n663), .A4(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT103), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n688), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  NOR2_X1   g518(.A1(new_n669), .A2(new_n670), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n560), .A2(new_n636), .A3(new_n675), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n612), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NAND2_X1  g522(.A1(new_n390), .A2(new_n269), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n388), .A2(new_n391), .B1(G469), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n600), .A3(new_n615), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n669), .ZN(new_n712));
  INV_X1    g526(.A(new_n461), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n638), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NOR2_X1   g531(.A1(new_n669), .A2(new_n713), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n649), .A2(new_n651), .ZN(new_n719));
  INV_X1    g533(.A(new_n711), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n718), .A2(new_n720), .A3(KEYINPUT105), .A4(new_n719), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NOR2_X1   g540(.A1(new_n699), .A2(new_n590), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n599), .A3(new_n663), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n712), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n712), .A2(KEYINPUT106), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  INV_X1    g548(.A(new_n710), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n601), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n301), .B1(new_n279), .B2(new_n258), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n305), .B(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n617), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n713), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n700), .B1(new_n614), .B2(new_n613), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n736), .A2(new_n741), .A3(new_n650), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND4_X1  g558(.A1(new_n706), .A2(new_n739), .A3(new_n663), .A4(new_n617), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n711), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n415), .ZN(G27));
  NAND2_X1  g561(.A1(new_n367), .A2(new_n269), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n601), .B1(new_n392), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n689), .A2(new_n603), .ZN(new_n751));
  AND4_X1   g565(.A1(KEYINPUT42), .A2(new_n750), .A3(new_n706), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n692), .A2(KEYINPUT109), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n667), .A2(new_n754), .A3(new_n668), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n291), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n461), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n758));
  NAND4_X1  g572(.A1(new_n310), .A2(new_n461), .A3(new_n750), .A4(new_n751), .ZN(new_n759));
  INV_X1    g573(.A(new_n706), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n680), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n676), .A2(new_n679), .A3(KEYINPUT110), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT111), .B(G134), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G36));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n367), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n609), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n372), .A2(new_n269), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n775), .A2(new_n776), .B1(new_n388), .B2(new_n391), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n601), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n684), .ZN(new_n780));
  INV_X1    g594(.A(new_n663), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n656), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n560), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n636), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n560), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n787), .A3(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT44), .B1(new_n782), .B2(new_n787), .ZN(new_n789));
  INV_X1    g603(.A(new_n751), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n780), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(G137), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G39));
  XOR2_X1   g608(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n795));
  OR2_X1    g609(.A1(new_n779), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n779), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n310), .A2(new_n790), .A3(new_n461), .A4(new_n760), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NOR3_X1   g615(.A1(new_n790), .A2(new_n735), .A3(new_n601), .ZN(new_n802));
  INV_X1    g616(.A(new_n598), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n461), .A3(new_n803), .A4(new_n698), .ZN(new_n804));
  INV_X1    g618(.A(new_n637), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n787), .A2(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n741), .ZN(new_n807));
  OAI221_X1 g621(.A(new_n597), .B1(new_n804), .B2(new_n805), .C1(new_n807), .C2(new_n711), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT121), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n756), .A2(new_n461), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n806), .A3(new_n802), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT48), .Z(new_n812));
  NOR2_X1   g626(.A1(new_n808), .A2(KEYINPUT121), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n809), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n804), .A2(new_n699), .A3(new_n785), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n806), .A2(new_n802), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n781), .A3(new_n740), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n691), .A2(new_n736), .A3(new_n603), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n807), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n807), .B2(new_n819), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n815), .B(new_n817), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n807), .A2(new_n790), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n796), .A2(new_n798), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n735), .A2(new_n600), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n826), .B2(KEYINPUT120), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n814), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n715), .A2(new_n743), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n725), .A2(new_n733), .A3(new_n762), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n746), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n663), .A2(new_n675), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n742), .A2(new_n697), .A3(new_n750), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n682), .A2(new_n707), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT52), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n746), .B1(new_n681), .B2(new_n612), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n707), .A4(new_n837), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n751), .A2(new_n663), .A3(new_n678), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n310), .A2(new_n393), .A3(new_n727), .A4(new_n600), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n750), .A2(new_n637), .A3(new_n617), .A4(new_n739), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n649), .B1(new_n560), .B2(new_n636), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n651), .A2(new_n603), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(new_n689), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n618), .A2(new_n849), .A3(new_n393), .A4(new_n600), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n607), .A3(new_n664), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n846), .A2(new_n851), .A3(new_n768), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n839), .A2(new_n842), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n725), .A2(new_n733), .A3(new_n762), .A4(new_n831), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n834), .A2(KEYINPUT53), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n857));
  NAND3_X1  g671(.A1(new_n839), .A2(new_n852), .A3(new_n842), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n854), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n862), .B(new_n857), .C1(new_n858), .C2(new_n854), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n856), .A2(new_n860), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n857), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n853), .A2(new_n832), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n858), .B2(new_n854), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT117), .B1(new_n869), .B2(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n871), .B(new_n861), .C1(new_n866), .C2(new_n868), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n864), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n830), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n461), .A2(new_n604), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT115), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n697), .A2(new_n786), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n710), .B(KEYINPUT49), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n691), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n874), .A2(new_n879), .ZN(G75));
  NAND3_X1  g694(.A1(new_n856), .A2(new_n860), .A3(new_n863), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(G902), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n884), .A3(G902), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n511), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n484), .A2(new_n496), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n494), .Z(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n260), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(G210), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n887), .B1(new_n882), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n892), .A2(new_n896), .ZN(G51));
  INV_X1    g711(.A(new_n885), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n884), .B1(new_n881), .B2(G902), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n773), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n881), .B(new_n861), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n774), .B(KEYINPUT57), .Z(new_n903));
  OAI21_X1  g717(.A(new_n390), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n893), .B1(new_n901), .B2(new_n904), .ZN(G54));
  AND2_X1   g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n552), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n883), .A2(new_n552), .A3(new_n885), .A4(new_n906), .ZN(new_n908));
  INV_X1    g722(.A(new_n893), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n907), .A2(new_n910), .ZN(G60));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n630), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n909), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n853), .B2(new_n832), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n858), .A2(new_n854), .A3(new_n857), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n871), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n869), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n913), .B1(new_n922), .B2(new_n864), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT123), .B1(new_n923), .B2(new_n630), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n873), .A2(new_n914), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n926));
  INV_X1    g740(.A(new_n630), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n916), .B1(new_n924), .B2(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n881), .A2(new_n661), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n881), .A2(new_n931), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n909), .B(new_n932), .C1(new_n933), .C2(new_n448), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G66));
  INV_X1    g750(.A(G224), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n595), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n725), .A2(new_n733), .A3(new_n831), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n851), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n888), .B1(G898), .B2(new_n260), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  AND2_X1   g757(.A1(new_n840), .A2(new_n707), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n703), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n703), .B(new_n944), .C1(new_n946), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n800), .A2(new_n792), .ZN(new_n951));
  INV_X1    g765(.A(new_n686), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n718), .A2(new_n751), .A3(new_n847), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n948), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n260), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n281), .B1(new_n284), .B2(KEYINPUT30), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n528), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n768), .B1(new_n757), .B2(new_n761), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT125), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n780), .A2(new_n742), .A3(new_n810), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n944), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n961), .A2(new_n951), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n260), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n958), .B1(G900), .B2(G953), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n968), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n959), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n969), .ZN(new_n974));
  INV_X1    g788(.A(new_n958), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n955), .B2(new_n260), .ZN(new_n976));
  OAI211_X1 g790(.A(KEYINPUT126), .B(new_n974), .C1(new_n976), .C2(new_n967), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n973), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n869), .ZN(new_n982));
  AOI211_X1 g796(.A(new_n981), .B(new_n982), .C1(new_n297), .C2(new_n288), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n287), .A2(new_n264), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n948), .A2(new_n940), .A3(new_n950), .A4(new_n954), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n980), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n964), .B2(new_n940), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n285), .A2(new_n286), .A3(new_n265), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n909), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n983), .B(new_n986), .C1(new_n991), .C2(new_n992), .ZN(G57));
endmodule


