//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(new_n456), .B2(G2106), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n469), .B2(KEYINPUT69), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT69), .A3(G125), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n476), .A2(new_n478), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT70), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n476), .B2(new_n478), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  AOI211_X1 g067(.A(new_n485), .B(new_n492), .C1(G136), .C2(new_n477), .ZN(G162));
  OAI211_X1 g068(.A(G138), .B(new_n478), .C1(new_n475), .C2(new_n466), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n478), .A3(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT71), .B1(new_n476), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n496), .A2(new_n478), .A3(G138), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n471), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n495), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n486), .B2(G126), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  OAI221_X1 g094(.A(new_n519), .B1(new_n515), .B2(new_n516), .C1(new_n513), .C2(new_n514), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n509), .B(G543), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n518), .A2(new_n520), .B1(G651), .B2(new_n524), .ZN(G166));
  AND2_X1   g100(.A1(new_n512), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n511), .A2(G89), .A3(new_n512), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n522), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n538), .B2(new_n537), .ZN(new_n540));
  INV_X1    g115(.A(new_n513), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT75), .B(G52), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n541), .A2(G90), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n534), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n513), .A2(new_n547), .B1(new_n548), .B2(new_n516), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT76), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n526), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n522), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n541), .A2(G91), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n540), .A2(new_n543), .ZN(G301));
  OR3_X1    g139(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT77), .B1(new_n531), .B2(new_n532), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  OR2_X1    g144(.A1(new_n511), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(G49), .B2(new_n526), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n541), .A2(new_n572), .A3(G87), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n572), .B1(new_n541), .B2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n522), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n526), .B2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n541), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G305));
  XNOR2_X1  g156(.A(KEYINPUT80), .B(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n513), .A2(new_n582), .B1(new_n583), .B2(new_n516), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT81), .Z(new_n585));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n522), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n534), .B1(new_n588), .B2(KEYINPUT79), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(KEYINPUT79), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n585), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n511), .A2(G92), .A3(new_n512), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n522), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n526), .B2(G54), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G321));
  NOR2_X1   g177(.A1(G299), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n567), .ZN(G297));
  AOI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n567), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(new_n606), .B2(G860), .ZN(G148));
  NOR2_X1   g182(.A1(new_n599), .A2(G559), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT82), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(KEYINPUT82), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n611), .B(new_n612), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n471), .A2(new_n479), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n478), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(G123), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n619), .B1(new_n620), .B2(new_n621), .C1(new_n490), .C2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n618), .A2(G2100), .B1(G2096), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n624), .B(new_n625), .C1(G2100), .C2(new_n618), .ZN(G156));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n632), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G14), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n644), .A2(new_n646), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(new_n647), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n644), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT84), .ZN(new_n658));
  OAI22_X1  g233(.A1(new_n657), .A2(KEYINPUT84), .B1(new_n647), .B2(new_n651), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT87), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n665), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  NAND2_X1  g260(.A1(G162), .A2(G29), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G29), .B2(G35), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT29), .B(G2090), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G1966), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NOR2_X1   g266(.A1(G168), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(G21), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n689), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n690), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(G171), .A2(new_n691), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G5), .B2(new_n691), .ZN(new_n697));
  INV_X1    g272(.A(G1961), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT100), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT30), .B(G28), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OR2_X1    g277(.A1(KEYINPUT31), .A2(G11), .ZN(new_n703));
  NAND2_X1  g278(.A1(KEYINPUT31), .A2(G11), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n701), .A2(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n705), .B1(new_n702), .B2(new_n623), .C1(new_n687), .C2(new_n688), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(G27), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G164), .B2(new_n702), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2078), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n691), .A2(G4), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n600), .B2(new_n691), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1348), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n691), .A2(G20), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT23), .Z(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G299), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1956), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n695), .A2(new_n700), .A3(new_n710), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G105), .B2(new_n479), .ZN(new_n724));
  INV_X1    g299(.A(G141), .ZN(new_n725));
  INV_X1    g300(.A(new_n477), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n491), .A2(G129), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(new_n702), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n702), .B2(G32), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n702), .B1(new_n733), .B2(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n733), .B2(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G160), .B2(G29), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n731), .A2(new_n732), .B1(G2084), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n698), .B2(new_n697), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT101), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n731), .A2(new_n732), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(G2084), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n702), .A2(G33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G139), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n726), .B2(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n478), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n742), .B1(new_n750), .B2(new_n702), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G2072), .Z(new_n752));
  NAND3_X1  g327(.A1(new_n740), .A2(new_n741), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n550), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT96), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G1341), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n702), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n762));
  INV_X1    g337(.A(G128), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n490), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n487), .A2(KEYINPUT97), .A3(new_n489), .A4(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n767));
  INV_X1    g342(.A(G116), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G2105), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n477), .B2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n761), .B1(new_n772), .B2(new_n702), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G2067), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n753), .A2(new_n754), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n755), .A2(new_n759), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n720), .A2(new_n739), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n691), .A2(G23), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G288), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT93), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n780), .B(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G22), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G166), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1971), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n691), .A2(G6), .ZN(new_n790));
  INV_X1    g365(.A(G305), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n691), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n783), .A2(new_n785), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n785), .B1(new_n783), .B2(new_n795), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n691), .A2(G24), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G290), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT90), .B(G1986), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n702), .A2(G25), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n487), .A2(G119), .A3(new_n489), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT89), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n478), .A2(G107), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n806), .A2(new_n807), .A3(new_n805), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n808), .A2(new_n809), .B1(new_n477), .B2(G131), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n804), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n803), .B1(new_n811), .B2(new_n702), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n801), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n796), .A2(KEYINPUT95), .A3(new_n797), .A4(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n777), .B1(new_n819), .B2(KEYINPUT36), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n796), .A2(new_n797), .A3(new_n816), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT36), .B1(new_n821), .B2(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n818), .B2(new_n817), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(G311));
  INV_X1    g399(.A(G311), .ZN(G150));
  NAND2_X1  g400(.A1(new_n600), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n534), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n513), .A2(new_n830), .B1(new_n831), .B2(new_n516), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n550), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n546), .A2(new_n549), .B1(new_n829), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n827), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n833), .A2(new_n840), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(G160), .B(new_n623), .ZN(new_n846));
  XNOR2_X1  g421(.A(G162), .B(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n766), .A2(G164), .A3(new_n770), .ZN(new_n848));
  AOI21_X1  g423(.A(G164), .B1(new_n766), .B2(new_n770), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n729), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n771), .A2(new_n507), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n727), .A2(new_n728), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n766), .A2(G164), .A3(new_n770), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n850), .A2(new_n854), .A3(new_n750), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n750), .B1(new_n850), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n477), .A2(G142), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(G2105), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n490), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n616), .A2(new_n804), .A3(new_n810), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n616), .B1(new_n810), .B2(new_n804), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n847), .B1(new_n857), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n871), .A2(KEYINPUT102), .A3(new_n872), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT102), .B1(new_n871), .B2(new_n872), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n855), .B2(new_n856), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n880));
  INV_X1    g455(.A(new_n750), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n848), .A2(new_n849), .A3(new_n729), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n850), .A2(new_n854), .A3(new_n750), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n875), .A2(new_n876), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT104), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n884), .A2(new_n889), .A3(new_n886), .A4(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n877), .B(new_n891), .C1(new_n855), .C2(new_n856), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n880), .A2(new_n888), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(new_n847), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n893), .B2(new_n847), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n879), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n899), .B(new_n879), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(G395));
  INV_X1    g478(.A(G868), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n836), .B(KEYINPUT107), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n609), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n599), .A2(G299), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n599), .A2(G299), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n906), .B(new_n608), .ZN(new_n917));
  INV_X1    g492(.A(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n905), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G290), .B(G303), .ZN(new_n922));
  XNOR2_X1  g497(.A(G288), .B(new_n791), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n916), .A2(new_n919), .A3(new_n905), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n924), .ZN(new_n927));
  INV_X1    g502(.A(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n920), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n904), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n833), .A2(G868), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n930), .A2(KEYINPUT108), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT108), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  OR2_X1    g509(.A1(new_n930), .A2(new_n931), .ZN(G331));
  NAND2_X1  g510(.A1(new_n567), .A2(G171), .ZN(new_n936));
  INV_X1    g511(.A(G168), .ZN(new_n937));
  NAND2_X1  g512(.A1(G301), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(new_n836), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n836), .B1(new_n936), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n911), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n936), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n837), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n936), .A2(new_n836), .A3(new_n938), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n911), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n946), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(KEYINPUT110), .A3(new_n914), .A4(new_n912), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n912), .A2(new_n944), .A3(new_n914), .A4(new_n945), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n927), .A2(new_n949), .A3(new_n951), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n951), .A2(new_n954), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(KEYINPUT112), .A3(new_n927), .A4(new_n949), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n952), .A2(new_n941), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n924), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT113), .A4(new_n961), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n951), .A2(new_n954), .ZN(new_n967));
  INV_X1    g542(.A(new_n949), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n924), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n957), .A2(new_n959), .A3(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(KEYINPUT44), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(KEYINPUT43), .B2(new_n962), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(KEYINPUT126), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n507), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n474), .A2(G40), .A3(new_n480), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n852), .A2(new_n984), .A3(G1996), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT114), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n771), .B(G2067), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n852), .A2(G1996), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n811), .A2(new_n813), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n811), .A2(new_n813), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n984), .ZN(new_n995));
  XOR2_X1   g570(.A(G290), .B(G1986), .Z(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n502), .B2(new_n506), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n982), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n980), .A2(KEYINPUT115), .A3(new_n981), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n983), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n980), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n474), .A2(G40), .A3(new_n480), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(KEYINPUT50), .B2(new_n980), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n717), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT57), .B1(new_n558), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(G299), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1007), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n983), .B1(KEYINPUT50), .B2(new_n980), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1348), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT116), .B1(new_n507), .B2(new_n979), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1006), .B(G1384), .C1(new_n502), .C2(new_n506), .ZN(new_n1023));
  NOR4_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n983), .A4(G2067), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1018), .B1(new_n599), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1004), .A2(new_n1016), .A3(new_n1012), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT121), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1004), .A2(new_n1012), .A3(new_n1016), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1018), .A2(KEYINPUT61), .A3(new_n1027), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n599), .B1(new_n1025), .B2(KEYINPUT60), .ZN(new_n1036));
  NOR4_X1   g611(.A1(new_n1021), .A2(new_n1024), .A3(new_n1034), .A4(new_n600), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n1039));
  INV_X1    g614(.A(G1996), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1010), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n981), .B(G1384), .C1(new_n502), .C2(new_n506), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1043), .A2(new_n1044), .A3(KEYINPUT115), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1001), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT58), .B(G1341), .Z(new_n1048));
  NAND2_X1  g623(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n983), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1041), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1048), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n1010), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT122), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1039), .B1(new_n1058), .B2(new_n550), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n546), .A2(new_n549), .ZN(new_n1060));
  AOI211_X1 g635(.A(KEYINPUT59), .B(new_n1060), .C1(new_n1052), .C2(new_n1057), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1033), .B(new_n1038), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT61), .B1(new_n1031), .B2(new_n1018), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1032), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT123), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n1032), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1010), .B1(new_n981), .B2(new_n980), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1049), .B2(new_n981), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1069), .A2(G1966), .B1(new_n1070), .B2(G2084), .ZN(new_n1071));
  OAI21_X1  g646(.A(G8), .B1(new_n1071), .B2(new_n937), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1044), .A2(new_n983), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1055), .B2(KEYINPUT45), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1073), .A2(new_n1074), .B1(new_n1076), .B2(new_n690), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G168), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1077), .B2(G168), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G303), .A2(G8), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT55), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1002), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1088));
  INV_X1    g663(.A(G2090), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1087), .A2(new_n788), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1090), .B2(new_n1080), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1080), .B1(new_n1055), .B2(new_n1010), .ZN(new_n1092));
  INV_X1    g667(.A(G1976), .ZN(new_n1093));
  OR2_X1    g668(.A1(G288), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT52), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1981), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n579), .A2(new_n1099), .A3(new_n580), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT118), .B(G86), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n541), .A2(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n579), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1103), .B2(new_n1099), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1100), .B(KEYINPUT49), .C1(new_n1103), .C2(new_n1099), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1096), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1085), .B(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1002), .A2(G1971), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1070), .A2(G2090), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1111), .B(G8), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1091), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1087), .B2(G2078), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1070), .A2(new_n698), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(G301), .B(KEYINPUT54), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT124), .B(G2078), .Z(new_n1121));
  NOR3_X1   g696(.A1(new_n1043), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1075), .B2(new_n1122), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1076), .A2(new_n1116), .A3(G2078), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1117), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1119), .A2(new_n1123), .B1(new_n1125), .B2(new_n1120), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1084), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1065), .A2(new_n1067), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1071), .A2(new_n937), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1082), .B1(new_n1081), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1072), .A2(KEYINPUT51), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT62), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1079), .A2(new_n1134), .A3(new_n1083), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1125), .A2(G171), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1133), .A2(new_n1135), .A3(new_n1115), .A4(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1077), .A2(new_n1080), .A3(G286), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1091), .A2(new_n1114), .A3(new_n1138), .A4(new_n1109), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(G8), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1086), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(new_n1138), .A3(KEYINPUT63), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1114), .A2(new_n1109), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1092), .B(KEYINPUT119), .Z(new_n1147));
  NOR2_X1   g722(.A1(G288), .A2(G1976), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1108), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1100), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1114), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1109), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1137), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n997), .B1(new_n1129), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n995), .A2(G290), .A3(G1986), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n994), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n984), .B1(new_n987), .B2(new_n852), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n984), .A2(new_n1040), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT46), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n771), .A2(G2067), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n990), .B2(new_n992), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n995), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n978), .B1(new_n1154), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1137), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1127), .B1(new_n1064), .B2(KEYINPUT123), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1067), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(KEYINPUT126), .B(new_n1168), .C1(new_n1173), .C2(new_n997), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1170), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g750(.A1(new_n898), .A2(new_n900), .ZN(new_n1177));
  OAI21_X1  g751(.A(G319), .B1(new_n640), .B2(new_n641), .ZN(new_n1178));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(G227), .B2(new_n1178), .ZN(new_n1179));
  OR3_X1    g753(.A1(G227), .A2(new_n1178), .A3(KEYINPUT127), .ZN(new_n1180));
  OAI211_X1 g754(.A(new_n1179), .B(new_n1180), .C1(new_n683), .C2(new_n684), .ZN(new_n1181));
  INV_X1    g755(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n974), .A3(new_n1182), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


