//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n207), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n216), .A2(new_n217), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n216), .B2(new_n217), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n203), .B2(new_n226), .C1(new_n227), .C2(new_n207), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G97), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n229), .B1(new_n202), .B2(new_n230), .C1(new_n231), .C2(new_n214), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n211), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n224), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n230), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n201), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n246), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(G1698), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT66), .B(G223), .Z(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n257), .B2(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n208), .A2(new_n267), .B1(new_n268), .B2(new_n261), .ZN(new_n269));
  XOR2_X1   g0069(.A(KEYINPUT65), .B(G226), .Z(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n262), .A3(G274), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n253), .B1(new_n264), .B2(new_n275), .ZN(new_n276));
  AOI211_X1 g0076(.A(KEYINPUT67), .B(new_n274), .C1(new_n260), .C2(new_n263), .ZN(new_n277));
  OAI21_X1  g0077(.A(G190), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n258), .A2(new_n259), .ZN(new_n279));
  OR2_X1    g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1698), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n282), .A2(G222), .B1(new_n285), .B2(G77), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n262), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT67), .B1(new_n287), .B2(new_n274), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n264), .A2(new_n253), .A3(new_n275), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(G200), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n209), .A3(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n218), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT69), .B1(new_n209), .B2(G1), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(new_n208), .A3(G20), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n201), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(new_n299), .B1(new_n201), .B2(new_n292), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n209), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n209), .A2(KEYINPUT68), .A3(G33), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G20), .A2(G33), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n294), .ZN(new_n311));
  OAI211_X1 g0111(.A(KEYINPUT9), .B(new_n300), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  INV_X1    g0113(.A(new_n300), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n307), .B2(new_n309), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n312), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n278), .A2(new_n290), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n320), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n278), .A2(new_n322), .A3(new_n290), .A4(new_n318), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT70), .B(G179), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n276), .B2(new_n277), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n288), .A2(new_n289), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n321), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT71), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n291), .A2(G1), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(G20), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n331), .A2(new_n208), .A3(G13), .A4(G20), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n294), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n296), .A2(new_n298), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G77), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G20), .A2(G77), .ZN(new_n339));
  INV_X1    g0139(.A(new_n308), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n339), .B1(new_n301), .B2(new_n340), .C1(new_n303), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n294), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n335), .A2(new_n257), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n338), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n282), .A2(G232), .ZN(new_n346));
  INV_X1    g0146(.A(G107), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n346), .B1(new_n347), .B2(new_n254), .C1(new_n258), .C2(new_n226), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n263), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n269), .A2(G244), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n273), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n345), .B1(new_n327), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n348), .B2(new_n263), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n324), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n345), .A2(KEYINPUT72), .B1(new_n353), .B2(G200), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n338), .A2(new_n343), .A3(new_n344), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n359), .A2(new_n360), .B1(new_n355), .B2(G190), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n330), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n305), .A2(G77), .A3(new_n306), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n365), .B1(new_n209), .B2(G68), .C1(new_n201), .C2(new_n340), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n294), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n336), .A2(G68), .A3(new_n337), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT12), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n335), .B2(new_n203), .ZN(new_n373));
  AND4_X1   g0173(.A1(new_n372), .A2(new_n332), .A3(G20), .A4(new_n203), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n367), .A2(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n255), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n230), .A2(G1698), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n378), .B(new_n379), .C1(new_n283), .C2(new_n284), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n263), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  INV_X1    g0184(.A(G274), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n268), .B2(new_n261), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n269), .A2(G238), .B1(new_n386), .B2(new_n272), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n262), .B1(new_n380), .B2(new_n381), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n262), .A2(G238), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n273), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT13), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(G190), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n383), .A2(new_n387), .A3(KEYINPUT74), .A4(new_n384), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n397), .A2(G200), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n376), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(G169), .A3(new_n398), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n397), .A2(KEYINPUT14), .A3(G169), .A4(new_n398), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n388), .A2(G179), .A3(new_n393), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT75), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT75), .ZN(new_n410));
  INV_X1    g0210(.A(new_n408), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n405), .C2(new_n406), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n402), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  OAI211_X1 g0214(.A(G226), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT77), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n254), .A2(KEYINPUT77), .A3(G226), .A4(G1698), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n254), .A2(G223), .A3(new_n255), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT78), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n263), .ZN(new_n424));
  INV_X1    g0224(.A(new_n324), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n262), .A2(G232), .A3(new_n390), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n262), .A2(new_n390), .A3(KEYINPUT79), .A4(G232), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n428), .A2(new_n429), .B1(new_n272), .B2(new_n386), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n327), .B1(new_n424), .B2(new_n430), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n414), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n428), .A2(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n273), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n263), .B2(new_n423), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT80), .B(new_n434), .C1(new_n437), .C2(new_n327), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT7), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n254), .B2(G20), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n203), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G58), .A2(G68), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT76), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(G58), .A3(G68), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n447), .A3(new_n220), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G20), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n308), .A2(G159), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n439), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT7), .B1(new_n285), .B2(new_n209), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n283), .A2(new_n284), .A3(new_n440), .A4(G20), .ZN(new_n454));
  OAI21_X1  g0254(.A(G68), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n448), .A2(G20), .B1(G159), .B2(new_n308), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(KEYINPUT16), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n457), .A3(new_n294), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n301), .B1(new_n298), .B2(new_n296), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(new_n295), .B1(new_n292), .B2(new_n301), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n433), .A2(new_n438), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT18), .ZN(new_n463));
  XOR2_X1   g0263(.A(KEYINPUT81), .B(G190), .Z(new_n464));
  AND3_X1   g0264(.A1(new_n424), .A2(new_n430), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(G200), .B1(new_n424), .B2(new_n430), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n458), .B(new_n460), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT17), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n424), .A2(new_n430), .A3(new_n464), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n437), .B2(G200), .ZN(new_n470));
  INV_X1    g0270(.A(new_n460), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n455), .A2(new_n456), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n311), .B1(new_n472), .B2(new_n439), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n473), .B2(new_n457), .ZN(new_n474));
  XOR2_X1   g0274(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT18), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n433), .A2(new_n438), .A3(new_n478), .A4(new_n461), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n463), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n364), .A2(new_n401), .A3(new_n413), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n484));
  OAI211_X1 g0284(.A(G244), .B(new_n255), .C1(new_n283), .C2(new_n284), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT4), .B1(new_n282), .B2(G244), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n263), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n266), .A2(G1), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G257), .A3(new_n262), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(KEYINPUT84), .A3(G257), .A4(new_n262), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n386), .B(new_n490), .C1(new_n492), .C2(new_n491), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n489), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G169), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n324), .B2(new_n500), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n292), .A2(new_n231), .ZN(new_n503));
  INV_X1    g0303(.A(G33), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n295), .B1(G1), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(new_n231), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  AND2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G97), .A2(G107), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n347), .A2(KEYINPUT6), .A3(G97), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n209), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n340), .A2(new_n257), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n514), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n347), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  XNOR2_X1  g0317(.A(G97), .B(G107), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n508), .ZN(new_n519));
  OAI211_X1 g0319(.A(KEYINPUT83), .B(new_n516), .C1(new_n519), .C2(new_n209), .ZN(new_n520));
  OAI21_X1  g0320(.A(G107), .B1(new_n453), .B2(new_n454), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n506), .B1(new_n522), .B2(new_n294), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n525), .B(new_n506), .C1(new_n522), .C2(new_n294), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n502), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n500), .A2(G200), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n489), .A2(new_n498), .A3(G190), .A4(new_n499), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n505), .ZN(new_n532));
  INV_X1    g0332(.A(new_n341), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n209), .B1(new_n381), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n510), .A2(new_n227), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n209), .B(G68), .C1(new_n283), .C2(new_n284), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n535), .B1(new_n303), .B2(new_n231), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n294), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n335), .A2(new_n341), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT87), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n534), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G238), .B(new_n255), .C1(new_n283), .C2(new_n284), .ZN(new_n547));
  OAI211_X1 g0347(.A(G244), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT86), .A2(G116), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(KEYINPUT86), .A2(G116), .ZN(new_n551));
  OAI21_X1  g0351(.A(G33), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n263), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n262), .A2(G274), .A3(new_n490), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n208), .A2(G45), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n262), .A2(G250), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(G169), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n263), .B2(new_n553), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n324), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n546), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G190), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n554), .A2(new_n564), .A3(new_n559), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G200), .B2(new_n561), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n532), .A2(G87), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n545), .C2(new_n544), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n493), .A2(G264), .A3(new_n262), .ZN(new_n569));
  INV_X1    g0369(.A(G294), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n504), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G250), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n214), .B2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(new_n254), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n499), .B(new_n569), .C1(new_n574), .C2(new_n262), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  INV_X1    g0376(.A(new_n569), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n207), .A2(new_n255), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n214), .A2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n283), .C2(new_n284), .ZN(new_n580));
  INV_X1    g0380(.A(new_n571), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n262), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT88), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT88), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n569), .C1(new_n574), .C2(new_n262), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n499), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G200), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n576), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n209), .B(G87), .C1(new_n283), .C2(new_n284), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n254), .A2(new_n591), .A3(new_n209), .A4(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT24), .ZN(new_n594));
  OR2_X1    g0394(.A1(KEYINPUT86), .A2(G116), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n504), .B1(new_n595), .B2(new_n549), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT23), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n209), .B2(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n347), .A2(KEYINPUT23), .A3(G20), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n596), .A2(new_n209), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n593), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n594), .B1(new_n593), .B2(new_n600), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n294), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n292), .A2(new_n347), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT25), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(G107), .B2(new_n532), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n563), .B(new_n568), .C1(new_n588), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n332), .A2(G20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT71), .ZN(new_n610));
  INV_X1    g0410(.A(new_n334), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n550), .A2(new_n551), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n208), .B2(G33), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n311), .B(new_n615), .C1(new_n333), .C2(new_n334), .ZN(new_n616));
  AOI21_X1  g0416(.A(G20), .B1(G33), .B2(G283), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n504), .A2(G97), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n618), .B1(new_n293), .B2(new_n218), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n595), .A2(G20), .A3(new_n549), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n619), .A2(KEYINPUT20), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT20), .B1(new_n619), .B2(new_n620), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n613), .B(new_n616), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G303), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n280), .A2(new_n624), .A3(new_n281), .ZN(new_n625));
  NOR2_X1   g0425(.A1(G257), .A2(G1698), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n215), .B2(G1698), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n263), .B(new_n625), .C1(new_n627), .C2(new_n285), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n493), .A2(G270), .A3(new_n262), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n499), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n623), .A2(KEYINPUT21), .A3(G169), .A4(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(G179), .A2(new_n628), .A3(new_n499), .A4(new_n629), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n623), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(G169), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT21), .B1(new_n636), .B2(new_n623), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n583), .A2(G179), .A3(new_n585), .A4(new_n499), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n575), .A2(G169), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n607), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n464), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n628), .A2(new_n499), .A3(new_n629), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n623), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n587), .B2(new_n644), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n638), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n482), .A2(new_n531), .A3(new_n608), .A4(new_n647), .ZN(G372));
  AND2_X1   g0448(.A1(new_n321), .A2(new_n323), .ZN(new_n649));
  INV_X1    g0449(.A(new_n477), .ZN(new_n650));
  INV_X1    g0450(.A(new_n357), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n399), .B2(new_n395), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n413), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n434), .B1(new_n437), .B2(new_n327), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n654), .A2(new_n478), .A3(new_n461), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n478), .B1(new_n654), .B2(new_n461), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n649), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n329), .ZN(new_n660));
  INV_X1    g0460(.A(new_n482), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n563), .B(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT21), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n621), .A2(new_n622), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n613), .A2(new_n616), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n667), .B2(new_n635), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n633), .A3(new_n631), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n603), .A2(new_n606), .B1(new_n639), .B2(new_n640), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n608), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n530), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n523), .B(KEYINPUT85), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n502), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n663), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(new_n523), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n502), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n563), .A2(new_n568), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n542), .A2(new_n543), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT87), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT87), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(G87), .B2(new_n532), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n686), .A2(new_n566), .B1(new_n546), .B2(new_n562), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n674), .A2(new_n502), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n681), .B1(new_n688), .B2(new_n677), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n676), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n661), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n660), .A2(new_n691), .ZN(G369));
  NOR2_X1   g0492(.A1(new_n607), .A2(new_n588), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n332), .A2(new_n209), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n603), .B2(new_n606), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n642), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n670), .A2(new_n700), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n638), .A2(new_n699), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n703), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n700), .A2(new_n667), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n669), .B(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(new_n646), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n710), .B1(new_n714), .B2(new_n704), .ZN(G399));
  NOR2_X1   g0515(.A1(new_n213), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n537), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n221), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(new_n679), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT26), .A3(new_n687), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n677), .B1(new_n527), .B2(new_n680), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n699), .B1(new_n676), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n699), .B1(new_n676), .B2(new_n689), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(KEYINPUT29), .B2(new_n728), .ZN(new_n729));
  NOR4_X1   g0529(.A1(new_n531), .A2(new_n647), .A3(new_n608), .A4(new_n699), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n583), .A2(new_n561), .A3(new_n585), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n489), .A2(new_n498), .A3(new_n499), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT30), .A4(new_n632), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n632), .A2(new_n561), .A3(new_n583), .A4(new_n585), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n735), .B2(new_n500), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n644), .A2(new_n561), .A3(new_n425), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n500), .A3(new_n586), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n699), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n730), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n729), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n721), .B1(new_n749), .B2(G1), .ZN(G364));
  NOR2_X1   g0550(.A1(new_n713), .A2(G330), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT90), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n291), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n208), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n716), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n752), .A2(new_n714), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n218), .B1(G20), .B2(new_n327), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n564), .A2(new_n587), .A3(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G179), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n254), .B1(new_n761), .B2(G329), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n763), .A2(new_n564), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n765), .A2(G303), .B1(new_n767), .B2(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n464), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n324), .A2(new_n209), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n762), .B(new_n768), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n324), .A2(new_n760), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n564), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n209), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n570), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n643), .A2(new_n770), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G326), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT93), .Z(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(new_n564), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n774), .B(new_n784), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n761), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  OR3_X1    g0590(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT32), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(new_n772), .C2(new_n202), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n775), .B(KEYINPUT92), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n257), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n764), .A2(new_n227), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G107), .B2(new_n767), .ZN(new_n798));
  INV_X1    g0598(.A(new_n779), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n285), .B1(new_n799), .B2(G97), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(new_n785), .C2(new_n203), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n781), .A2(new_n201), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n793), .A2(new_n796), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n759), .B1(new_n788), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n212), .A2(new_n254), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(KEYINPUT91), .B2(G355), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(KEYINPUT91), .B2(G355), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n251), .A2(new_n266), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n213), .A2(new_n254), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(G45), .B2(new_n221), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n807), .B1(G116), .B2(new_n212), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n759), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n757), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n814), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n804), .B(new_n816), .C1(new_n713), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n758), .A2(new_n818), .ZN(G396));
  OAI21_X1  g0619(.A(new_n254), .B1(new_n779), .B2(new_n202), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n201), .A2(new_n764), .B1(new_n766), .B2(new_n203), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT95), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G132), .C2(new_n761), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n781), .A2(new_n824), .B1(new_n785), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT94), .Z(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n772), .C1(new_n790), .C2(new_n795), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n285), .B1(new_n231), .B2(new_n779), .C1(new_n772), .C2(new_n570), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n795), .A2(new_n612), .B1(new_n624), .B2(new_n781), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n766), .A2(new_n227), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G311), .B2(new_n761), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n347), .B2(new_n764), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n785), .A2(new_n838), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n833), .A2(new_n834), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n759), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n759), .A2(new_n812), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n757), .B1(new_n257), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n357), .A2(new_n699), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n359), .A2(new_n699), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n362), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n357), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n841), .B(new_n843), .C1(new_n813), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT96), .B1(new_n728), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n728), .A2(new_n847), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n747), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n757), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(new_n747), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(G384));
  INV_X1    g0655(.A(new_n519), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(G116), .A4(new_n219), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  NAND4_X1  g0660(.A1(new_n222), .A2(G77), .A3(new_n447), .A4(new_n445), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n208), .B(G13), .C1(new_n861), .C2(new_n247), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n728), .A2(new_n847), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n844), .B(KEYINPUT97), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  INV_X1    g0668(.A(new_n697), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n461), .B2(new_n869), .ZN(new_n870));
  AOI211_X1 g0670(.A(KEYINPUT98), .B(new_n697), .C1(new_n458), .C2(new_n460), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n452), .A2(new_n457), .A3(new_n294), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n873), .A2(new_n471), .B1(new_n431), .B2(new_n432), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n467), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n470), .B2(new_n474), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n461), .A2(new_n869), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n462), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n480), .A2(new_n872), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(KEYINPUT98), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n461), .A2(new_n868), .A3(new_n869), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n874), .A2(new_n467), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n879), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT38), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(KEYINPUT18), .A2(new_n462), .B1(new_n468), .B2(new_n476), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n884), .B1(new_n889), .B2(new_n479), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n880), .A2(KEYINPUT38), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n411), .B1(new_n405), .B2(new_n406), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT75), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n402), .B(new_n699), .C1(new_n893), .C2(new_n400), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n402), .A2(new_n699), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n413), .A2(new_n401), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n867), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n657), .A2(new_n869), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n888), .A2(new_n890), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n874), .A2(KEYINPUT18), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n654), .A2(new_n478), .A3(new_n461), .ZN(new_n905));
  INV_X1    g0705(.A(new_n475), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n467), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT17), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n470), .B2(new_n474), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n904), .B(new_n905), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n878), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n874), .A2(new_n878), .A3(new_n467), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n910), .A2(new_n911), .B1(new_n913), .B2(new_n879), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n903), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT100), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n480), .A2(new_n872), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n876), .A2(new_n879), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT100), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n878), .B1(new_n657), .B2(new_n477), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n878), .A2(new_n467), .A3(new_n881), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n923), .A2(new_n462), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n919), .A2(new_n920), .A3(new_n925), .A4(new_n903), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n916), .A2(new_n926), .B1(KEYINPUT39), .B2(new_n891), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n893), .A2(KEYINPUT99), .A3(new_n402), .A4(new_n700), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n402), .B(new_n700), .C1(new_n409), .C2(new_n412), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT99), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n901), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n659), .A2(new_n329), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT29), .B1(new_n690), .B2(new_n700), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT29), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n938), .B(new_n699), .C1(new_n676), .C2(new_n725), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n936), .B1(new_n940), .B2(new_n661), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n935), .B(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n888), .A2(new_n890), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT101), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT101), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n919), .A2(new_n945), .A3(new_n925), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n846), .A2(new_n357), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n651), .A2(new_n700), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n743), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT31), .B1(new_n739), .B2(new_n699), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n647), .A2(new_n608), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n675), .A3(new_n700), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n950), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n413), .A2(new_n401), .A3(new_n895), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n895), .B1(new_n413), .B2(new_n401), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(KEYINPUT40), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n891), .A2(new_n897), .A3(new_n956), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n947), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n482), .B2(new_n745), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n661), .A3(new_n746), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(G330), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n942), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n208), .B2(new_n753), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n942), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n863), .B1(new_n969), .B2(new_n970), .ZN(G367));
  AOI21_X1  g0771(.A(new_n531), .B1(new_n678), .B2(new_n699), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT102), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n974), .A2(new_n975), .B1(new_n722), .B2(new_n699), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n714), .A2(new_n704), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT104), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n686), .A2(new_n700), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n680), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n663), .B2(new_n981), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n980), .B(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n976), .A2(new_n708), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n527), .B1(new_n976), .B2(new_n642), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT103), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n700), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n984), .B2(new_n983), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n986), .B(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n716), .B(KEYINPUT41), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n976), .A2(new_n709), .ZN(new_n997));
  XNOR2_X1  g0797(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n997), .B(new_n998), .Z(new_n999));
  INV_X1    g0799(.A(KEYINPUT109), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n978), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n977), .A2(new_n710), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n976), .B2(new_n709), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1004), .A2(new_n1006), .B1(new_n1000), .B2(new_n978), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n999), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1002), .B1(new_n999), .B2(new_n1007), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n704), .B(new_n706), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(new_n714), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n748), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(KEYINPUT108), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT108), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n996), .B1(new_n1023), .B2(new_n749), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n995), .B1(new_n1024), .B2(new_n755), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n809), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n815), .B1(new_n212), .B2(new_n341), .C1(new_n1026), .C2(new_n242), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n766), .A2(new_n257), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G58), .B2(new_n765), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n824), .B2(new_n789), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n254), .B1(new_n203), .B2(new_n779), .C1(new_n772), .C2(new_n825), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(G143), .C2(new_n782), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n794), .A2(G50), .B1(new_n786), .B2(G159), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n767), .A2(G97), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n347), .C2(new_n779), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G311), .B2(new_n782), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n612), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT46), .B1(new_n765), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(G317), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n285), .B1(new_n789), .B2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n771), .C2(G303), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n794), .A2(G283), .B1(new_n786), .B2(G294), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1040), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT47), .Z(new_n1049));
  INV_X1    g0849(.A(new_n759), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n756), .B(new_n1027), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT111), .Z(new_n1052));
  INV_X1    g0852(.A(new_n983), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n817), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1025), .A2(new_n1054), .ZN(G387));
  AOI21_X1  g0855(.A(new_n717), .B1(new_n748), .B2(new_n1013), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1019), .A2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n805), .A2(new_n718), .B1(G107), .B2(new_n212), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n239), .A2(new_n266), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n718), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n1060), .C1(G68), .C2(G77), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n301), .A2(G50), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1026), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1058), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n815), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n756), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n781), .A2(new_n773), .B1(new_n785), .B2(new_n777), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT114), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT114), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n794), .A2(G303), .B1(new_n771), .B2(G317), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n799), .A2(G283), .B1(new_n765), .B2(G294), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n285), .B1(new_n766), .B2(new_n612), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G326), .B2(new_n761), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n771), .A2(G50), .B1(new_n533), .B2(new_n799), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT113), .Z(new_n1085));
  NOR2_X1   g0885(.A1(new_n781), .A2(new_n790), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT112), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n775), .A2(G68), .B1(G150), .B2(new_n761), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n765), .A2(G77), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1088), .A2(new_n254), .A3(new_n1038), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n302), .B2(new_n786), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1085), .A2(new_n1087), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1067), .B1(new_n1093), .B2(new_n759), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1094), .A2(KEYINPUT115), .B1(new_n704), .B2(new_n814), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(KEYINPUT115), .B2(new_n1094), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1013), .A2(new_n754), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1057), .A2(new_n1099), .ZN(G393));
  NOR2_X1   g0900(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n717), .B1(new_n1101), .B2(new_n1019), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1023), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n976), .A2(new_n814), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n815), .B1(new_n231), .B2(new_n212), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n809), .B2(new_n246), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n772), .A2(new_n790), .B1(new_n781), .B2(new_n825), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n789), .A2(new_n828), .B1(new_n764), .B2(new_n203), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n779), .A2(new_n257), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n835), .A4(new_n285), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n794), .A2(new_n302), .B1(new_n786), .B2(G50), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n772), .A2(new_n777), .B1(new_n781), .B2(new_n1043), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n285), .B1(new_n766), .B2(new_n347), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n776), .A2(new_n570), .B1(new_n612), .B2(new_n779), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G303), .C2(new_n786), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n789), .A2(new_n773), .B1(new_n764), .B2(new_n838), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT116), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT117), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n757), .B(new_n1106), .C1(new_n1123), .C2(new_n759), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1011), .A2(new_n755), .B1(new_n1104), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1103), .A2(new_n1125), .ZN(G390));
  INV_X1    g0926(.A(KEYINPUT121), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n916), .A2(new_n926), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n865), .B1(new_n728), .B2(new_n847), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n957), .A2(new_n958), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n933), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n676), .A2(new_n725), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n700), .A3(new_n948), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n949), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n897), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n929), .A2(KEYINPUT118), .A3(new_n932), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT118), .B1(new_n929), .B2(new_n932), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n947), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n897), .A2(G330), .A3(new_n956), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1133), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n754), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n927), .A2(new_n812), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n842), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n756), .B1(new_n302), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT120), .Z(new_n1149));
  AOI211_X1 g0949(.A(new_n254), .B(new_n797), .C1(new_n771), .C2(G116), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1110), .B1(G68), .B2(new_n767), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n570), .C2(new_n789), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n794), .A2(G97), .B1(new_n786), .B2(G107), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n838), .B2(new_n781), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n794), .A2(new_n1156), .B1(new_n786), .B2(G137), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n779), .A2(new_n790), .B1(new_n766), .B2(new_n201), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n285), .B(new_n1158), .C1(G125), .C2(new_n761), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1157), .B(new_n1159), .C1(new_n1160), .C2(new_n781), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT53), .B1(new_n764), .B2(new_n825), .ZN(new_n1162));
  OR3_X1    g0962(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n825), .ZN(new_n1163));
  INV_X1    g0963(.A(G132), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1163), .C1(new_n772), .C2(new_n1164), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1152), .A2(new_n1154), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1149), .B1(new_n1166), .B2(new_n759), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1145), .B1(new_n1146), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1133), .A2(new_n1141), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1142), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1133), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n661), .A2(G330), .A3(new_n746), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n660), .B(new_n1173), .C1(new_n482), .C2(new_n729), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n847), .B1(new_n730), .B2(new_n744), .ZN(new_n1175));
  INV_X1    g0975(.A(G330), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n896), .B(new_n894), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1129), .B1(new_n1142), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n844), .B1(new_n726), .B2(new_n948), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1142), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1174), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1171), .A2(new_n1172), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(KEYINPUT119), .A3(new_n716), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1142), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n941), .B(new_n1173), .C1(new_n1185), .C2(new_n1178), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT119), .B1(new_n1183), .B2(new_n716), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1127), .B(new_n1168), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT119), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1143), .A2(new_n1144), .A3(new_n1186), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n717), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n1187), .A3(new_n1184), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1127), .B1(new_n1195), .B2(new_n1168), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1191), .A2(new_n1196), .ZN(G378));
  AOI21_X1  g0997(.A(new_n1175), .B1(new_n896), .B2(new_n894), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n919), .A2(new_n945), .A3(new_n925), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n945), .B1(new_n919), .B2(new_n925), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1198), .B(KEYINPUT40), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n917), .A2(new_n918), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n921), .B1(new_n876), .B2(new_n879), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1203), .A2(new_n921), .B1(new_n917), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n962), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(G330), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n326), .A2(new_n869), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n330), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n321), .A2(new_n323), .A3(new_n329), .A4(new_n1208), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1207), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n898), .B(new_n900), .C1(new_n927), .C2(new_n933), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT124), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1215), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(KEYINPUT124), .A3(new_n1213), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1201), .A2(new_n1224), .A3(G330), .A4(new_n1206), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1218), .A2(new_n1219), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1219), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n755), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n812), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n756), .B1(G50), .B2(new_n1147), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT123), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n781), .A2(new_n614), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n776), .A2(new_n341), .B1(new_n202), .B2(new_n766), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1089), .B1(new_n838), .B2(new_n789), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n285), .A2(new_n265), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n799), .B2(G68), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1235), .B(new_n1237), .C1(new_n347), .C2(new_n772), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1232), .B(new_n1238), .C1(G97), .C2(new_n786), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(KEYINPUT58), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT58), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1236), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n504), .B(new_n265), .C1(new_n766), .C2(new_n790), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n775), .A2(G137), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n765), .A2(new_n1156), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n1164), .B2(new_n785), .C1(new_n772), .C2(new_n1160), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n782), .A2(G125), .B1(G150), .B2(new_n799), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(KEYINPUT122), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(KEYINPUT122), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1248), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT59), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1244), .B(new_n1255), .C1(G124), .C2(new_n761), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(KEYINPUT59), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1243), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1229), .B(new_n1231), .C1(new_n1050), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1228), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1174), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1216), .B1(new_n963), .B2(G330), .ZN(new_n1263));
  AND4_X1   g1063(.A1(G330), .A2(new_n1201), .A3(new_n1206), .A4(new_n1224), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n935), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1218), .A2(new_n1219), .A3(new_n1225), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1262), .A2(new_n1183), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n717), .B1(new_n1267), .B2(KEYINPUT57), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1183), .A2(new_n1262), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1261), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(G375));
  NOR2_X1   g1075(.A1(new_n1185), .A2(new_n1178), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1130), .A2(new_n812), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n756), .B1(G68), .B2(new_n1147), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n254), .B(new_n1028), .C1(new_n771), .C2(G283), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n799), .A2(new_n533), .B1(G303), .B2(new_n761), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(new_n231), .C2(new_n764), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n794), .A2(G107), .B1(new_n786), .B2(new_n1041), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n570), .B2(new_n781), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n776), .A2(new_n825), .B1(new_n201), .B2(new_n779), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n789), .A2(new_n1160), .B1(new_n764), .B2(new_n790), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n285), .B1(new_n767), .B2(G58), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(new_n824), .C2(new_n772), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n781), .A2(new_n1164), .B1(new_n785), .B2(new_n1155), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n1282), .A2(new_n1284), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1279), .B1(new_n1291), .B2(new_n759), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(KEYINPUT125), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1277), .A2(new_n755), .B1(new_n1278), .B2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1277), .A2(new_n1262), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n996), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1186), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1295), .B2(new_n1297), .ZN(G381));
  NOR2_X1   g1098(.A1(G393), .A2(G396), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(G381), .A2(G384), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1103), .A2(new_n1125), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1168), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1302));
  OR4_X1    g1102(.A1(G387), .A2(new_n1301), .A3(new_n1302), .A4(G375), .ZN(G407));
  INV_X1    g1103(.A(new_n1302), .ZN(new_n1304));
  INV_X1    g1104(.A(G213), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1305), .A2(G343), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1274), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(G407), .A2(G213), .A3(new_n1307), .ZN(G409));
  AND2_X1   g1108(.A1(G393), .A2(G396), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(new_n1299), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(G390), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1103), .B(new_n1125), .C1(new_n1309), .C2(new_n1299), .ZN(new_n1312));
  AND4_X1   g1112(.A1(new_n1025), .A2(new_n1311), .A3(new_n1054), .A4(new_n1312), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1311), .A2(new_n1312), .B1(new_n1025), .B2(new_n1054), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1302), .A2(KEYINPUT121), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1274), .A2(new_n1316), .A3(new_n1190), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1269), .A2(new_n1270), .A3(new_n1296), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1267), .A2(KEYINPUT126), .A3(new_n1296), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1228), .A4(new_n1260), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1304), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1317), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1306), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1186), .A2(KEYINPUT60), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n717), .B1(new_n1326), .B2(new_n1295), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1295), .B2(new_n1326), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1294), .ZN(new_n1329));
  INV_X1    g1129(.A(G384), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(G384), .A3(new_n1294), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1324), .A2(new_n1325), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT127), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1324), .A2(new_n1337), .A3(new_n1325), .A4(new_n1334), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT62), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1306), .A2(G2897), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1331), .A2(new_n1332), .A3(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1261), .B1(new_n1319), .B2(new_n1318), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1302), .B1(new_n1344), .B2(new_n1321), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(G378), .B2(new_n1274), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1343), .B1(new_n1346), .B2(new_n1306), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  AOI211_X1 g1149(.A(new_n1306), .B(new_n1333), .C1(new_n1317), .C2(new_n1323), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1347), .B(new_n1348), .C1(new_n1349), .C2(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1315), .B1(new_n1339), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1336), .A2(new_n1353), .A3(new_n1338), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1350), .A2(KEYINPUT63), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1354), .A2(new_n1355), .A3(new_n1356), .A4(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1352), .A2(new_n1358), .ZN(G405));
  OAI21_X1  g1159(.A(new_n1317), .B1(new_n1302), .B2(new_n1274), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1333), .ZN(new_n1361));
  XNOR2_X1  g1161(.A(new_n1361), .B(new_n1356), .ZN(G402));
endmodule


