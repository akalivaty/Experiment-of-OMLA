//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT2), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n208), .A3(KEYINPUT2), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT74), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(new_n209), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n211), .A2(new_n212), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n213), .A2(new_n214), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n222), .A2(new_n224), .A3(new_n207), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n227));
  AND2_X1   g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n212), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n220), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n222), .A2(new_n207), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n223), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  INV_X1    g038(.A(G113gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G120gat), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245));
  INV_X1    g044(.A(G127gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(G134gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(G134gat), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n245), .A2(KEYINPUT1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n237), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n235), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n250), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n232), .A2(new_n231), .B1(new_n234), .B2(new_n223), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n244), .A2(new_n249), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT4), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n251), .A2(new_n254), .A3(new_n257), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n253), .A2(new_n252), .A3(new_n250), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT4), .B1(new_n255), .B2(new_n256), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT78), .A3(new_n251), .A4(new_n261), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n250), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n233), .A2(new_n235), .B1(new_n244), .B2(new_n249), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n260), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT76), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n254), .A3(new_n257), .A4(new_n259), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n260), .C1(new_n270), .C2(new_n271), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n273), .A2(new_n274), .A3(new_n258), .A4(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n206), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n269), .A2(new_n206), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n280), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n278), .B1(new_n283), .B2(KEYINPUT79), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n285), .A3(new_n280), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n281), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT26), .B1(new_n289), .B2(new_n290), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n297), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT28), .B1(new_n297), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n302), .A2(new_n304), .A3(new_n294), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n298), .A3(KEYINPUT67), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n307), .A2(new_n309), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n313), .A3(KEYINPUT25), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(new_n298), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n307), .A4(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n305), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n321), .B2(KEYINPUT66), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  AOI211_X1 g122(.A(new_n323), .B(new_n315), .C1(new_n305), .C2(new_n320), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n301), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n326), .B(KEYINPUT72), .Z(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n327), .B(new_n301), .C1(new_n322), .C2(new_n324), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT70), .ZN(new_n333));
  NAND2_X1  g132(.A1(G211gat), .A2(G218gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(new_n333), .A3(new_n335), .ZN(new_n342));
  INV_X1    g141(.A(G197gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G204gat), .ZN(new_n344));
  INV_X1    g143(.A(G204gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G197gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n339), .A2(new_n341), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT71), .B(new_n340), .C1(new_n347), .C2(new_n336), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n351), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n330), .A2(new_n353), .A3(new_n331), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n352), .A2(KEYINPUT73), .A3(new_n354), .A4(new_n357), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n352), .B2(new_n354), .ZN(new_n364));
  INV_X1    g163(.A(new_n358), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(KEYINPUT30), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n202), .B1(new_n287), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n363), .A2(new_n366), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n282), .A2(new_n285), .A3(new_n280), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n285), .B1(new_n282), .B2(new_n280), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n370), .A2(new_n371), .A3(new_n278), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n369), .B(KEYINPUT80), .C1(new_n372), .C2(new_n281), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n325), .A2(new_n250), .ZN(new_n374));
  INV_X1    g173(.A(G227gat), .ZN(new_n375));
  INV_X1    g174(.A(G233gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n256), .B(new_n301), .C1(new_n322), .C2(new_n324), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n383), .A3(new_n381), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G15gat), .B(G43gat), .Z(new_n386));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n378), .B1(new_n374), .B2(new_n379), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(KEYINPUT33), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT32), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n379), .ZN(new_n394));
  AOI221_X4 g193(.A(new_n391), .B1(KEYINPUT33), .B2(new_n388), .C1(new_n394), .C2(new_n377), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n385), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n377), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n400), .A3(new_n388), .ZN(new_n401));
  INV_X1    g200(.A(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n384), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT81), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n411), .B(KEYINPUT82), .Z(new_n412));
  NAND3_X1  g211(.A1(new_n349), .A2(new_n328), .A3(new_n350), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n255), .B1(new_n413), .B2(new_n236), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n237), .A2(new_n328), .B1(new_n350), .B2(new_n349), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n415), .A2(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n414), .A2(new_n417), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n410), .B(new_n416), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n413), .A2(new_n236), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n253), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT83), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n418), .A3(new_n419), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n410), .B1(new_n427), .B2(new_n416), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n409), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n409), .C1(new_n423), .C2(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G22gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n422), .A3(new_n408), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT85), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n435), .A2(new_n438), .A3(new_n422), .A4(new_n408), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n405), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n368), .A2(new_n373), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT35), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n283), .A2(new_n278), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n281), .ZN(new_n445));
  OR3_X1    g244(.A1(new_n445), .A2(KEYINPUT35), .A3(new_n367), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n433), .A2(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(new_n405), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n283), .A2(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(new_n279), .A3(new_n286), .ZN(new_n453));
  INV_X1    g252(.A(new_n281), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT80), .B1(new_n455), .B2(new_n369), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n287), .A2(new_n202), .A3(new_n367), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n385), .A2(new_n393), .A3(new_n395), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n403), .B1(new_n401), .B2(new_n402), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n396), .A2(new_n404), .A3(new_n459), .A4(new_n460), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n251), .A2(new_n254), .A3(new_n257), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n260), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n270), .A2(new_n271), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT39), .B1(new_n471), .B2(new_n260), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n259), .B1(new_n267), .B2(new_n251), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n206), .B(new_n470), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT87), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT86), .B1(new_n479), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n278), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n433), .A2(new_n440), .B1(new_n482), .B2(new_n367), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n352), .A2(new_n484), .A3(new_n354), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n357), .B1(new_n485), .B2(KEYINPUT89), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(KEYINPUT89), .B2(new_n485), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n352), .B2(new_n354), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT38), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n360), .A2(new_n362), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n352), .A2(new_n491), .A3(new_n354), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n353), .B1(new_n330), .B2(new_n331), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n484), .B1(new_n493), .B2(KEYINPUT88), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT38), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n486), .C1(KEYINPUT89), .C2(new_n485), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n489), .A2(new_n445), .A3(new_n490), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n467), .B1(new_n483), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n443), .A2(new_n450), .B1(new_n458), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G197gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT11), .B(G169gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n501), .B(new_n502), .Z(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT12), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g304(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  INV_X1    g309(.A(G29gat), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G43gat), .ZN(new_n515));
  INV_X1    g314(.A(G43gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G50gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT15), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT91), .B1(new_n516), .B2(G50gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(G43gat), .B2(new_n514), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(KEYINPUT91), .A3(G50gat), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT15), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n508), .ZN(new_n525));
  OAI221_X1 g324(.A(new_n518), .B1(new_n511), .B2(new_n512), .C1(new_n525), .C2(new_n506), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n520), .A2(KEYINPUT17), .A3(new_n527), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(G1gat), .B2(new_n532), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(G8gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(G8gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n539), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT92), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n530), .A2(new_n531), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT93), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n542), .A2(new_n540), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n531), .A4(new_n530), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n541), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n544), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n528), .A2(new_n554), .A3(new_n541), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n528), .B2(new_n541), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n549), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n548), .B(KEYINPUT13), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n550), .B2(new_n551), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n505), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(KEYINPUT95), .A3(new_n551), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n559), .B(new_n504), .C1(new_n550), .C2(new_n551), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT95), .B1(new_n550), .B2(new_n551), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  NAND3_X1  g376(.A1(new_n530), .A2(new_n531), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n575), .B(new_n576), .ZN(new_n581));
  AND2_X1   g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n528), .A2(new_n581), .B1(KEYINPUT41), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n578), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n580), .B1(new_n578), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n582), .A2(KEYINPUT41), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n595), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n600), .B2(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n594), .B(KEYINPUT98), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n581), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n577), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G230gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n376), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n609), .A2(new_n612), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n246), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n541), .B1(new_n608), .B2(KEYINPUT21), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n638), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n216), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n592), .B(new_n632), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n499), .A2(new_n568), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n287), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n367), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(G8gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G8gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT42), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(KEYINPUT42), .B2(new_n656), .ZN(G1325gat));
  INV_X1    g457(.A(G15gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n659), .A3(new_n448), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n650), .A2(new_n467), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n662), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n650), .A2(new_n451), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n443), .A2(new_n450), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n447), .B1(new_n368), .B2(new_n373), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n498), .B1(new_n669), .B2(KEYINPUT104), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n671), .B(new_n447), .C1(new_n368), .C2(new_n373), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  INV_X1    g473(.A(new_n592), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n677), .B(KEYINPUT44), .C1(new_n499), .C2(new_n592), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n458), .A2(new_n498), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n446), .A2(new_n449), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(KEYINPUT35), .B2(new_n442), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n675), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n677), .B1(new_n683), .B2(KEYINPUT44), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n641), .B(new_n646), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(new_n568), .A3(new_n631), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G29gat), .B1(new_n688), .B2(new_n455), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n458), .A2(new_n498), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n592), .B1(new_n668), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n687), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n455), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(G1328gat));
  OAI21_X1  g494(.A(G36gat), .B1(new_n688), .B2(new_n369), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n692), .A2(G36gat), .A3(new_n369), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(new_n467), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n516), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n687), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n516), .B1(new_n692), .B2(new_n405), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT47), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n702), .A2(new_n709), .A3(new_n703), .A4(new_n704), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n708), .A3(new_n710), .ZN(G1330gat));
  OAI211_X1 g510(.A(new_n451), .B(new_n687), .C1(new_n679), .C2(new_n684), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n447), .A2(G50gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n713), .B(KEYINPUT48), .C1(new_n692), .C2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT107), .B1(new_n692), .B2(new_n715), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n691), .A2(new_n718), .A3(new_n687), .A4(new_n714), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n720), .B1(new_n712), .B2(G50gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT48), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n716), .B1(new_n724), .B2(new_n727), .ZN(G1331gat));
  INV_X1    g527(.A(new_n686), .ZN(new_n729));
  INV_X1    g528(.A(new_n568), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n729), .A2(new_n730), .A3(new_n675), .A4(new_n632), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n673), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n287), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n369), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n732), .B2(new_n700), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n405), .A2(G71gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n451), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g546(.A1(new_n673), .A2(new_n675), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n686), .A2(new_n730), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT51), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n632), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n572), .A3(new_n287), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n686), .A2(new_n730), .A3(new_n632), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n685), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n455), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1336gat));
  NOR2_X1   g557(.A1(new_n369), .A2(G92gat), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n631), .B(new_n759), .C1(new_n750), .C2(new_n751), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n367), .B(new_n755), .C1(new_n679), .C2(new_n684), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT110), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1337gat));
  INV_X1    g566(.A(G99gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n768), .A3(new_n448), .ZN(new_n769));
  OAI21_X1  g568(.A(G99gat), .B1(new_n756), .B2(new_n700), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  NOR2_X1   g570(.A1(new_n447), .A2(G106gat), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n631), .B(new_n772), .C1(new_n750), .C2(new_n751), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n451), .B(new_n755), .C1(new_n679), .C2(new_n684), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g576(.A1(new_n649), .A2(new_n730), .ZN(new_n778));
  INV_X1    g577(.A(new_n565), .ZN(new_n779));
  INV_X1    g578(.A(new_n566), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n563), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n503), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(G229gat), .A3(G233gat), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n557), .A2(new_n558), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n781), .A2(new_n787), .A3(KEYINPUT112), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n619), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n617), .B1(new_n613), .B2(new_n614), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n629), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n630), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n792), .B2(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n792), .A2(new_n795), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(KEYINPUT111), .A3(new_n630), .A4(new_n796), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n675), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT112), .B1(new_n781), .B2(new_n787), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n789), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n799), .B(new_n803), .C1(new_n562), .C2(new_n567), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n787), .A3(new_n631), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n675), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n729), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n778), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n455), .A2(new_n367), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n441), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n568), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n803), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n808), .B1(new_n568), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n592), .ZN(new_n817));
  INV_X1    g616(.A(new_n804), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n781), .A2(new_n787), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n821), .A3(new_n788), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n686), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n649), .A2(new_n730), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n287), .B(new_n441), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n367), .B1(new_n825), .B2(KEYINPUT113), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n827), .A3(new_n287), .A4(new_n441), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n730), .A2(new_n240), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n814), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT114), .Z(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n813), .B2(new_n632), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n631), .A2(new_n242), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT115), .Z(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n829), .B2(new_n835), .ZN(G1341gat));
  NOR3_X1   g635(.A1(new_n813), .A2(new_n246), .A3(new_n729), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT116), .Z(new_n838));
  NAND3_X1  g637(.A1(new_n826), .A2(new_n686), .A3(new_n828), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n246), .B2(new_n839), .ZN(G1342gat));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n592), .A2(G134gat), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(new_n828), .A3(new_n369), .A4(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n826), .A2(KEYINPUT117), .A3(new_n828), .A4(new_n842), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n813), .B2(new_n592), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n845), .A2(new_n847), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(KEYINPUT56), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT118), .B(new_n846), .C1(new_n845), .C2(new_n847), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n823), .A2(new_n824), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n455), .ZN(new_n857));
  INV_X1    g656(.A(G141gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n467), .A2(new_n367), .A3(new_n447), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n730), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n447), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n567), .A2(new_n632), .A3(new_n786), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n802), .A2(new_n630), .A3(new_n796), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n781), .B2(new_n561), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n592), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n686), .B1(new_n822), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(new_n824), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT119), .B(new_n862), .C1(new_n867), .C2(new_n824), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n447), .B1(new_n778), .B2(new_n810), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n870), .B(new_n871), .C1(KEYINPUT57), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n700), .A2(new_n812), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n873), .A2(new_n730), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n860), .B1(new_n876), .B2(new_n858), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n879), .B(new_n860), .C1(new_n876), .C2(new_n858), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n631), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n864), .A2(KEYINPUT121), .A3(new_n592), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT121), .B1(new_n864), .B2(new_n592), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n821), .A2(new_n883), .A3(new_n788), .A4(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n866), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n778), .B1(new_n886), .B2(new_n686), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n451), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n811), .A2(new_n862), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n631), .A3(new_n875), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n892), .A2(KEYINPUT59), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n894), .A2(KEYINPUT120), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n857), .A2(new_n892), .A3(new_n631), .A4(new_n859), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1345gat));
  NAND2_X1  g699(.A1(new_n811), .A2(new_n451), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n901), .A2(new_n861), .B1(new_n869), .B2(new_n868), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n874), .B1(new_n902), .B2(new_n871), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n216), .B1(new_n903), .B2(new_n686), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n857), .A2(new_n859), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(G155gat), .A3(new_n729), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n904), .A2(new_n906), .ZN(G1346gat));
  NAND3_X1  g706(.A1(new_n903), .A2(G162gat), .A3(new_n675), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n217), .B1(new_n905), .B2(new_n592), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1347gat));
  NAND2_X1  g713(.A1(new_n455), .A2(new_n367), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n856), .A2(new_n449), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n730), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n631), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT123), .B(G176gat), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n916), .A2(new_n686), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n308), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n297), .B2(new_n922), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g724(.A1(new_n916), .A2(new_n675), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(G190gat), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(G190gat), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1351gat));
  NOR2_X1   g730(.A1(new_n467), .A2(new_n915), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n872), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(G197gat), .A3(new_n568), .ZN(new_n934));
  INV_X1    g733(.A(new_n890), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n730), .B(new_n932), .C1(new_n935), .C2(new_n888), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n936), .B2(G197gat), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT125), .ZN(G1352gat));
  NOR3_X1   g737(.A1(new_n933), .A2(G204gat), .A3(new_n632), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT62), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n467), .B(new_n915), .C1(new_n889), .C2(new_n890), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(new_n631), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(new_n345), .ZN(G1353gat));
  OR3_X1    g742(.A1(new_n933), .A2(G211gat), .A3(new_n729), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n686), .B(new_n932), .C1(new_n935), .C2(new_n888), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  NAND2_X1  g747(.A1(new_n675), .A2(G218gat), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT126), .ZN(new_n950));
  INV_X1    g749(.A(G218gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n872), .A2(new_n675), .A3(new_n932), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n941), .A2(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1355gat));
endmodule


