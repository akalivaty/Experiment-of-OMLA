

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n721), .ZN(n511) );
  NAND2_X2 U549 ( .A1(n678), .A2(n760), .ZN(n721) );
  NOR2_X2 U550 ( .A1(G2105), .A2(n537), .ZN(n868) );
  AND2_X1 U551 ( .A1(G160), .A2(G40), .ZN(n678) );
  OR2_X1 U552 ( .A1(n744), .A2(n754), .ZN(n512) );
  OR2_X1 U553 ( .A1(n758), .A2(n757), .ZN(n513) );
  AND2_X1 U554 ( .A1(n916), .A2(n805), .ZN(n514) );
  INV_X1 U555 ( .A(G168), .ZN(n711) );
  AND2_X1 U556 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U557 ( .A1(n715), .A2(n714), .ZN(n717) );
  NOR2_X1 U558 ( .A1(n754), .A2(G1966), .ZN(n708) );
  NAND2_X1 U559 ( .A1(n921), .A2(n512), .ZN(n745) );
  NOR2_X1 U560 ( .A1(n793), .A2(n514), .ZN(n794) );
  NOR2_X2 U561 ( .A1(G2104), .A2(n536), .ZN(n861) );
  NOR2_X1 U562 ( .A1(G651), .A2(n636), .ZN(n646) );
  AND2_X1 U563 ( .A1(n541), .A2(n540), .ZN(G160) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U565 ( .A1(n642), .A2(G89), .ZN(n515) );
  XNOR2_X1 U566 ( .A(KEYINPUT4), .B(n515), .ZN(n518) );
  XOR2_X1 U567 ( .A(G543), .B(KEYINPUT0), .Z(n636) );
  INV_X1 U568 ( .A(G651), .ZN(n520) );
  NOR2_X1 U569 ( .A1(n636), .A2(n520), .ZN(n643) );
  NAND2_X1 U570 ( .A1(n643), .A2(G76), .ZN(n516) );
  XOR2_X1 U571 ( .A(KEYINPUT69), .B(n516), .Z(n517) );
  NAND2_X1 U572 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U573 ( .A(n519), .B(KEYINPUT5), .ZN(n527) );
  NOR2_X1 U574 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n521), .Z(n647) );
  NAND2_X1 U576 ( .A1(n647), .A2(G63), .ZN(n522) );
  XNOR2_X1 U577 ( .A(n522), .B(KEYINPUT70), .ZN(n524) );
  NAND2_X1 U578 ( .A1(G51), .A2(n646), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n525), .Z(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U582 ( .A(n528), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U584 ( .A(KEYINPUT23), .ZN(n530) );
  INV_X1 U585 ( .A(G2104), .ZN(n537) );
  NAND2_X1 U586 ( .A1(G101), .A2(n868), .ZN(n529) );
  XNOR2_X1 U587 ( .A(n530), .B(n529), .ZN(n533) );
  INV_X1 U588 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G125), .A2(n861), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n531), .B(KEYINPUT64), .ZN(n532) );
  AND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n541) );
  XNOR2_X1 U592 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n535) );
  NOR2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XNOR2_X2 U594 ( .A(n535), .B(n534), .ZN(n865) );
  AND2_X1 U595 ( .A1(G137), .A2(n865), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n860) );
  AND2_X1 U597 ( .A1(G113), .A2(n860), .ZN(n538) );
  NOR2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U599 ( .A1(G102), .A2(n868), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G138), .A2(n865), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G114), .A2(n860), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G126), .A2(n861), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U606 ( .A1(G85), .A2(n642), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G72), .A2(n643), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G47), .A2(n646), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G60), .A2(n647), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U612 ( .A1(n553), .A2(n552), .ZN(G290) );
  XNOR2_X1 U613 ( .A(G2454), .B(G2443), .ZN(n563) );
  XOR2_X1 U614 ( .A(KEYINPUT96), .B(G2430), .Z(n555) );
  XNOR2_X1 U615 ( .A(G2446), .B(KEYINPUT97), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n555), .B(n554), .ZN(n559) );
  XOR2_X1 U617 ( .A(G2451), .B(G2427), .Z(n557) );
  XNOR2_X1 U618 ( .A(G1348), .B(G1341), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U620 ( .A(n559), .B(n558), .Z(n561) );
  XNOR2_X1 U621 ( .A(G2435), .B(G2438), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n563), .B(n562), .ZN(n564) );
  AND2_X1 U624 ( .A1(n564), .A2(G14), .ZN(G401) );
  NAND2_X1 U625 ( .A1(G52), .A2(n646), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G64), .A2(n647), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G90), .A2(n642), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G77), .A2(n643), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U632 ( .A1(n571), .A2(n570), .ZN(G171) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U634 ( .A1(G123), .A2(n861), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT18), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G135), .A2(n865), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G111), .A2(n860), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n868), .A2(G99), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(n575), .Z(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n992) );
  XNOR2_X1 U643 ( .A(G2096), .B(n992), .ZN(n580) );
  OR2_X1 U644 ( .A1(G2100), .A2(n580), .ZN(G156) );
  INV_X1 U645 ( .A(G132), .ZN(G219) );
  INV_X1 U646 ( .A(G82), .ZN(G220) );
  INV_X1 U647 ( .A(G120), .ZN(G236) );
  INV_X1 U648 ( .A(G57), .ZN(G237) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U650 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n811) );
  NAND2_X1 U652 ( .A1(n811), .A2(G567), .ZN(n582) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  XOR2_X1 U654 ( .A(G860), .B(KEYINPUT67), .Z(n612) );
  NAND2_X1 U655 ( .A1(n642), .A2(G81), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G68), .A2(n643), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT13), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G43), .A2(n646), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n647), .A2(G56), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(n589), .Z(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT66), .B(n592), .Z(n881) );
  INV_X1 U666 ( .A(n881), .ZN(n615) );
  NAND2_X1 U667 ( .A1(n612), .A2(n615), .ZN(G153) );
  XOR2_X1 U668 ( .A(G171), .B(KEYINPUT68), .Z(G301) );
  NAND2_X1 U669 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G54), .A2(n646), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G66), .A2(n647), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G92), .A2(n642), .ZN(n596) );
  NAND2_X1 U674 ( .A1(G79), .A2(n643), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n599), .B(KEYINPUT15), .ZN(n910) );
  INV_X1 U678 ( .A(G868), .ZN(n660) );
  NAND2_X1 U679 ( .A1(n910), .A2(n660), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U681 ( .A1(G91), .A2(n642), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G78), .A2(n643), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G53), .A2(n646), .ZN(n605) );
  NAND2_X1 U685 ( .A1(G65), .A2(n647), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n901) );
  NAND2_X1 U688 ( .A1(n901), .A2(n660), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT71), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n660), .A2(G286), .ZN(n609) );
  NOR2_X1 U691 ( .A1(n610), .A2(n609), .ZN(G297) );
  INV_X1 U692 ( .A(n901), .ZN(G299) );
  INV_X1 U693 ( .A(G559), .ZN(n611) );
  NOR2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n910), .A2(n613), .ZN(n614) );
  XOR2_X1 U696 ( .A(KEYINPUT16), .B(n614), .Z(G148) );
  INV_X1 U697 ( .A(n615), .ZN(n900) );
  NOR2_X1 U698 ( .A1(n900), .A2(G868), .ZN(n618) );
  INV_X1 U699 ( .A(n910), .ZN(n640) );
  NAND2_X1 U700 ( .A1(G868), .A2(n640), .ZN(n616) );
  NOR2_X1 U701 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U702 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U703 ( .A1(G86), .A2(n642), .ZN(n620) );
  NAND2_X1 U704 ( .A1(G61), .A2(n647), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U706 ( .A(KEYINPUT76), .B(n621), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n643), .A2(G73), .ZN(n622) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n646), .A2(G48), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U712 ( .A1(G88), .A2(n642), .ZN(n628) );
  NAND2_X1 U713 ( .A1(G75), .A2(n643), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G50), .A2(n646), .ZN(n630) );
  NAND2_X1 U716 ( .A1(G62), .A2(n647), .ZN(n629) );
  NAND2_X1 U717 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n632), .A2(n631), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G49), .A2(n646), .ZN(n634) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U722 ( .A1(n647), .A2(n635), .ZN(n639) );
  NAND2_X1 U723 ( .A1(G87), .A2(n636), .ZN(n637) );
  XOR2_X1 U724 ( .A(KEYINPUT75), .B(n637), .Z(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G559), .A2(n640), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n641), .B(n900), .ZN(n895) );
  NAND2_X1 U728 ( .A1(G93), .A2(n642), .ZN(n645) );
  NAND2_X1 U729 ( .A1(G80), .A2(n643), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G55), .A2(n646), .ZN(n649) );
  NAND2_X1 U732 ( .A1(G67), .A2(n647), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U735 ( .A(KEYINPUT74), .B(n652), .Z(n894) );
  XNOR2_X1 U736 ( .A(n894), .B(G290), .ZN(n653) );
  XNOR2_X1 U737 ( .A(n653), .B(G305), .ZN(n654) );
  XOR2_X1 U738 ( .A(n654), .B(KEYINPUT19), .Z(n656) );
  XNOR2_X1 U739 ( .A(G166), .B(KEYINPUT77), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U741 ( .A(n657), .B(G299), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(G288), .ZN(n884) );
  XNOR2_X1 U743 ( .A(n895), .B(n884), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n659), .A2(G868), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n894), .A2(n660), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n666), .A2(G2072), .ZN(n667) );
  XNOR2_X1 U752 ( .A(KEYINPUT78), .B(n667), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G237), .A2(G236), .ZN(n668) );
  NAND2_X1 U755 ( .A1(G69), .A2(n668), .ZN(n669) );
  XNOR2_X1 U756 ( .A(KEYINPUT79), .B(n669), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n670), .A2(G108), .ZN(n898) );
  NAND2_X1 U758 ( .A1(G567), .A2(n898), .ZN(n675) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U761 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U762 ( .A1(G96), .A2(n673), .ZN(n899) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n899), .ZN(n674) );
  NAND2_X1 U764 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U765 ( .A(KEYINPUT80), .B(n676), .ZN(n888) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n677) );
  NOR2_X1 U767 ( .A1(n888), .A2(n677), .ZN(n817) );
  NAND2_X1 U768 ( .A1(n817), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n760) );
  NAND2_X1 U771 ( .A1(G8), .A2(n721), .ZN(n754) );
  NAND2_X1 U772 ( .A1(G1348), .A2(n721), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G2067), .A2(n511), .ZN(n679) );
  NAND2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n691) );
  AND2_X1 U775 ( .A1(n910), .A2(n691), .ZN(n681) );
  OR2_X1 U776 ( .A1(n881), .A2(n681), .ZN(n687) );
  NAND2_X1 U777 ( .A1(G1996), .A2(n511), .ZN(n682) );
  XNOR2_X1 U778 ( .A(n682), .B(KEYINPUT26), .ZN(n684) );
  NAND2_X1 U779 ( .A1(G1341), .A2(n721), .ZN(n683) );
  NAND2_X1 U780 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U781 ( .A(KEYINPUT88), .B(n685), .ZN(n686) );
  NOR2_X1 U782 ( .A1(n687), .A2(n686), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n511), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U784 ( .A(n688), .B(KEYINPUT27), .ZN(n690) );
  INV_X1 U785 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U786 ( .A1(n949), .A2(n511), .ZN(n689) );
  NOR2_X1 U787 ( .A1(n690), .A2(n689), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n696), .A2(n901), .ZN(n693) );
  OR2_X1 U789 ( .A1(n910), .A2(n691), .ZN(n692) );
  NAND2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n696), .A2(n901), .ZN(n698) );
  INV_X1 U793 ( .A(KEYINPUT28), .ZN(n697) );
  XNOR2_X1 U794 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U796 ( .A(KEYINPUT29), .B(KEYINPUT89), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n702), .B(n701), .ZN(n706) );
  OR2_X1 U798 ( .A1(n511), .A2(G1961), .ZN(n704) );
  XNOR2_X1 U799 ( .A(KEYINPUT25), .B(G2078), .ZN(n928) );
  NAND2_X1 U800 ( .A1(n511), .A2(n928), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n713) );
  NAND2_X1 U802 ( .A1(G171), .A2(n713), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U804 ( .A(n707), .B(KEYINPUT90), .ZN(n719) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n721), .ZN(n730) );
  XNOR2_X1 U806 ( .A(n708), .B(KEYINPUT87), .ZN(n732) );
  NAND2_X1 U807 ( .A1(G8), .A2(n732), .ZN(n709) );
  NOR2_X1 U808 ( .A1(n730), .A2(n709), .ZN(n710) );
  XNOR2_X1 U809 ( .A(n710), .B(KEYINPUT30), .ZN(n712) );
  NOR2_X1 U810 ( .A1(G171), .A2(n713), .ZN(n714) );
  INV_X1 U811 ( .A(KEYINPUT31), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n731) );
  NAND2_X1 U814 ( .A1(n731), .A2(G286), .ZN(n726) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n754), .ZN(n720) );
  XOR2_X1 U816 ( .A(KEYINPUT91), .B(n720), .Z(n723) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n721), .ZN(n722) );
  NOR2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n724), .A2(G303), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U821 ( .A(n727), .B(KEYINPUT92), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n728), .A2(G8), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n729), .B(KEYINPUT32), .ZN(n736) );
  NAND2_X1 U824 ( .A1(G8), .A2(n730), .ZN(n734) );
  AND2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n749) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n743) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n743), .A2(n737), .ZN(n904) );
  NAND2_X1 U831 ( .A1(n749), .A2(n904), .ZN(n738) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n903) );
  NAND2_X1 U833 ( .A1(n738), .A2(n903), .ZN(n739) );
  XNOR2_X1 U834 ( .A(KEYINPUT93), .B(n739), .ZN(n740) );
  INV_X1 U835 ( .A(n740), .ZN(n741) );
  NOR2_X1 U836 ( .A1(n754), .A2(n741), .ZN(n742) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n742), .ZN(n746) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n921) );
  NAND2_X1 U839 ( .A1(n743), .A2(KEYINPUT33), .ZN(n744) );
  NOR2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n758) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n747) );
  XNOR2_X1 U842 ( .A(n747), .B(KEYINPUT94), .ZN(n748) );
  NAND2_X1 U843 ( .A1(n748), .A2(G8), .ZN(n750) );
  NAND2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U845 ( .A1(n751), .A2(n754), .ZN(n756) );
  NOR2_X1 U846 ( .A1(G1981), .A2(G305), .ZN(n752) );
  XOR2_X1 U847 ( .A(n752), .B(KEYINPUT24), .Z(n753) );
  OR2_X1 U848 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U849 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U850 ( .A1(G160), .A2(G40), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n805) );
  XOR2_X1 U852 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n772) );
  NAND2_X1 U853 ( .A1(G104), .A2(n868), .ZN(n762) );
  NAND2_X1 U854 ( .A1(G140), .A2(n865), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U856 ( .A(KEYINPUT34), .B(n763), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G116), .A2(n860), .ZN(n765) );
  NAND2_X1 U858 ( .A1(G128), .A2(n861), .ZN(n764) );
  NAND2_X1 U859 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U860 ( .A(KEYINPUT82), .B(n766), .Z(n767) );
  XNOR2_X1 U861 ( .A(KEYINPUT35), .B(n767), .ZN(n768) );
  NOR2_X1 U862 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U863 ( .A(n770), .B(KEYINPUT36), .ZN(n771) );
  XNOR2_X1 U864 ( .A(n772), .B(n771), .ZN(n877) );
  XOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .Z(n773) );
  XNOR2_X1 U866 ( .A(KEYINPUT81), .B(n773), .ZN(n803) );
  NOR2_X1 U867 ( .A1(n877), .A2(n803), .ZN(n998) );
  NAND2_X1 U868 ( .A1(n805), .A2(n998), .ZN(n801) );
  XOR2_X1 U869 ( .A(KEYINPUT86), .B(KEYINPUT38), .Z(n775) );
  NAND2_X1 U870 ( .A1(G105), .A2(n868), .ZN(n774) );
  XNOR2_X1 U871 ( .A(n775), .B(n774), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G117), .A2(n860), .ZN(n777) );
  NAND2_X1 U873 ( .A1(G129), .A2(n861), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U875 ( .A(KEYINPUT85), .B(n778), .Z(n779) );
  NOR2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U877 ( .A1(n865), .A2(G141), .ZN(n781) );
  NAND2_X1 U878 ( .A1(n782), .A2(n781), .ZN(n846) );
  AND2_X1 U879 ( .A1(n846), .A2(G1996), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G95), .A2(n868), .ZN(n784) );
  NAND2_X1 U881 ( .A1(G131), .A2(n865), .ZN(n783) );
  NAND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G107), .A2(n860), .ZN(n786) );
  NAND2_X1 U884 ( .A1(G119), .A2(n861), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U886 ( .A1(n788), .A2(n787), .ZN(n873) );
  INV_X1 U887 ( .A(G1991), .ZN(n795) );
  NOR2_X1 U888 ( .A1(n873), .A2(n795), .ZN(n789) );
  NOR2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n990) );
  INV_X1 U890 ( .A(n805), .ZN(n791) );
  NOR2_X1 U891 ( .A1(n990), .A2(n791), .ZN(n798) );
  INV_X1 U892 ( .A(n798), .ZN(n792) );
  NAND2_X1 U893 ( .A1(n801), .A2(n792), .ZN(n793) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n916) );
  NAND2_X1 U895 ( .A1(n513), .A2(n794), .ZN(n808) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n846), .ZN(n987) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n796) );
  AND2_X1 U898 ( .A1(n795), .A2(n873), .ZN(n995) );
  NOR2_X1 U899 ( .A1(n796), .A2(n995), .ZN(n797) );
  NOR2_X1 U900 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U901 ( .A1(n987), .A2(n799), .ZN(n800) );
  XNOR2_X1 U902 ( .A(n800), .B(KEYINPUT39), .ZN(n802) );
  NAND2_X1 U903 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U904 ( .A1(n877), .A2(n803), .ZN(n999) );
  NAND2_X1 U905 ( .A1(n804), .A2(n999), .ZN(n806) );
  NAND2_X1 U906 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n810) );
  XOR2_X1 U908 ( .A(KEYINPUT40), .B(KEYINPUT95), .Z(n809) );
  XNOR2_X1 U909 ( .A(n810), .B(n809), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n811), .ZN(G217) );
  INV_X1 U911 ( .A(G661), .ZN(n813) );
  NAND2_X1 U912 ( .A1(G2), .A2(G15), .ZN(n812) );
  NOR2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U914 ( .A(KEYINPUT98), .B(n814), .Z(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n815) );
  XOR2_X1 U916 ( .A(KEYINPUT99), .B(n815), .Z(n816) );
  NAND2_X1 U917 ( .A1(n817), .A2(n816), .ZN(G188) );
  XOR2_X1 U918 ( .A(G69), .B(KEYINPUT100), .Z(G235) );
  XOR2_X1 U919 ( .A(G2100), .B(G2096), .Z(n819) );
  XNOR2_X1 U920 ( .A(KEYINPUT42), .B(G2678), .ZN(n818) );
  XNOR2_X1 U921 ( .A(n819), .B(n818), .ZN(n823) );
  XOR2_X1 U922 ( .A(KEYINPUT43), .B(G2090), .Z(n821) );
  XNOR2_X1 U923 ( .A(G2067), .B(G2072), .ZN(n820) );
  XNOR2_X1 U924 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U925 ( .A(n823), .B(n822), .Z(n825) );
  XNOR2_X1 U926 ( .A(G2084), .B(G2078), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(G227) );
  XOR2_X1 U928 ( .A(KEYINPUT103), .B(G1981), .Z(n827) );
  XNOR2_X1 U929 ( .A(G1996), .B(G1991), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n828), .B(KEYINPUT41), .Z(n830) );
  XNOR2_X1 U932 ( .A(G1971), .B(G1976), .ZN(n829) );
  XNOR2_X1 U933 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U934 ( .A(G1956), .B(G1961), .Z(n832) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1966), .ZN(n831) );
  XNOR2_X1 U936 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U937 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U938 ( .A(KEYINPUT102), .B(G2474), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(G229) );
  NAND2_X1 U940 ( .A1(G124), .A2(n861), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n837), .B(KEYINPUT104), .ZN(n838) );
  XNOR2_X1 U942 ( .A(KEYINPUT44), .B(n838), .ZN(n841) );
  NAND2_X1 U943 ( .A1(G100), .A2(n868), .ZN(n839) );
  XOR2_X1 U944 ( .A(KEYINPUT105), .B(n839), .Z(n840) );
  NAND2_X1 U945 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U946 ( .A1(G136), .A2(n865), .ZN(n843) );
  NAND2_X1 U947 ( .A1(G112), .A2(n860), .ZN(n842) );
  NAND2_X1 U948 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U949 ( .A1(n845), .A2(n844), .ZN(G162) );
  XNOR2_X1 U950 ( .A(n992), .B(G162), .ZN(n848) );
  XOR2_X1 U951 ( .A(G160), .B(n846), .Z(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G118), .A2(n860), .ZN(n850) );
  NAND2_X1 U954 ( .A1(G130), .A2(n861), .ZN(n849) );
  NAND2_X1 U955 ( .A1(n850), .A2(n849), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G106), .A2(n868), .ZN(n852) );
  NAND2_X1 U957 ( .A1(G142), .A2(n865), .ZN(n851) );
  NAND2_X1 U958 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U959 ( .A(n853), .B(KEYINPUT45), .Z(n854) );
  NOR2_X1 U960 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U961 ( .A(n857), .B(n856), .Z(n879) );
  XOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n859) );
  XNOR2_X1 U963 ( .A(KEYINPUT108), .B(KEYINPUT48), .ZN(n858) );
  XNOR2_X1 U964 ( .A(n859), .B(n858), .ZN(n872) );
  NAND2_X1 U965 ( .A1(G115), .A2(n860), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G127), .A2(n861), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n864), .B(KEYINPUT47), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G139), .A2(n865), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n868), .A2(G103), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT106), .B(n869), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n982) );
  XOR2_X1 U974 ( .A(n872), .B(n982), .Z(n875) );
  XNOR2_X1 U975 ( .A(G164), .B(n873), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n877), .B(n876), .Z(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U979 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U980 ( .A(n910), .B(KEYINPUT109), .ZN(n883) );
  XNOR2_X1 U981 ( .A(G171), .B(n881), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n886) );
  XOR2_X1 U983 ( .A(G286), .B(n884), .Z(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U985 ( .A1(G37), .A2(n887), .ZN(G397) );
  XNOR2_X1 U986 ( .A(KEYINPUT101), .B(n888), .ZN(G319) );
  NOR2_X1 U987 ( .A1(G227), .A2(G229), .ZN(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT49), .B(n889), .ZN(n890) );
  NOR2_X1 U989 ( .A1(G401), .A2(n890), .ZN(n892) );
  NOR2_X1 U990 ( .A1(G395), .A2(G397), .ZN(n891) );
  AND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n893), .A2(G319), .ZN(G225) );
  XOR2_X1 U993 ( .A(KEYINPUT110), .B(G225), .Z(G308) );
  XNOR2_X1 U995 ( .A(n894), .B(KEYINPUT73), .ZN(n897) );
  NOR2_X1 U996 ( .A1(n895), .A2(G860), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(G145) );
  INV_X1 U998 ( .A(G108), .ZN(G238) );
  INV_X1 U999 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(G325) );
  INV_X1 U1001 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1002 ( .A(n900), .B(G1341), .Z(n919) );
  NAND2_X1 U1003 ( .A1(G303), .A2(G1971), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n901), .B(KEYINPUT118), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(n902), .B(n949), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1007 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(KEYINPUT119), .ZN(n914) );
  XOR2_X1 U1010 ( .A(G171), .B(G1961), .Z(n912) );
  XNOR2_X1 U1011 ( .A(n910), .B(G1348), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT120), .B(n917), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n925) );
  XOR2_X1 U1017 ( .A(G1966), .B(G168), .Z(n920) );
  XNOR2_X1 U1018 ( .A(KEYINPUT117), .B(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1020 ( .A(KEYINPUT57), .B(n923), .Z(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1022 ( .A(KEYINPUT56), .B(G16), .Z(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n1013) );
  XNOR2_X1 U1024 ( .A(G1991), .B(G25), .ZN(n938) );
  XNOR2_X1 U1025 ( .A(G27), .B(n928), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G32), .B(G1996), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT114), .B(G2072), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G33), .B(n933), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(KEYINPUT115), .B(n936), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(G28), .A2(n939), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT53), .B(n940), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT116), .B(G34), .Z(n942) );
  XNOR2_X1 U1038 ( .A(G2084), .B(KEYINPUT54), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G35), .B(G2090), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n975) );
  NAND2_X1 U1043 ( .A1(KEYINPUT55), .A2(n975), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(G11), .A2(n947), .ZN(n981) );
  XNOR2_X1 U1045 ( .A(KEYINPUT121), .B(G1961), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(G5), .ZN(n961) );
  XNOR2_X1 U1047 ( .A(G20), .B(n949), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G1341), .B(G19), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G1981), .B(G6), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1052 ( .A(KEYINPUT59), .B(G1348), .Z(n954) );
  XNOR2_X1 U1053 ( .A(G4), .B(n954), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1055 ( .A(KEYINPUT60), .B(n957), .Z(n959) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G21), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n970) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n966) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G22), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(G23), .B(G1976), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(n964), .B(KEYINPUT122), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1065 ( .A(KEYINPUT58), .B(n967), .Z(n968) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n968), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1068 ( .A(n971), .B(KEYINPUT124), .Z(n972) );
  XNOR2_X1 U1069 ( .A(KEYINPUT61), .B(n972), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(G16), .A2(n973), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(KEYINPUT125), .B(n974), .ZN(n979) );
  INV_X1 U1072 ( .A(n975), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(G29), .A2(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n1011) );
  XOR2_X1 U1077 ( .A(G2072), .B(n982), .Z(n984) );
  XOR2_X1 U1078 ( .A(G164), .B(G2078), .Z(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1080 ( .A(KEYINPUT50), .B(n985), .Z(n1005) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1083 ( .A(KEYINPUT112), .B(n988), .Z(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT51), .B(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(G160), .B(G2084), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT111), .B(n996), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT113), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT52), .B(n1006), .ZN(n1008) );
  INV_X1 U1096 ( .A(KEYINPUT55), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(G29), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1015), .ZN(G150) );
  INV_X1 U1103 ( .A(G150), .ZN(G311) );
endmodule

