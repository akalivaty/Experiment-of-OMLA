//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n464), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n475), .B(new_n477), .C1(G124), .C2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n484), .A2(new_n486), .A3(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(new_n464), .A3(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n480), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n489), .B2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT68), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n462), .A2(new_n496), .A3(new_n464), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n488), .B1(new_n494), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT69), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n505), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n509), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n506), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n514), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n507), .A2(new_n531), .B1(new_n509), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AND2_X1   g109(.A1(new_n505), .A2(G56), .ZN(new_n535));
  AND2_X1   g110(.A1(G68), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT70), .ZN(new_n538));
  INV_X1    g113(.A(new_n507), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT71), .B(G81), .Z(new_n540));
  INV_X1    g115(.A(new_n509), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(G43), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n537), .A2(KEYINPUT70), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND3_X1  g125(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n507), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n558), .A2(new_n529), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  OAI21_X1  g140(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n566));
  INV_X1    g141(.A(G49), .ZN(new_n567));
  INV_X1    g142(.A(G87), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n566), .B1(new_n509), .B2(new_n567), .C1(new_n568), .C2(new_n507), .ZN(G288));
  NAND3_X1  g144(.A1(new_n505), .A2(new_n506), .A3(G86), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n541), .A2(G48), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n505), .A2(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n529), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n539), .A2(KEYINPUT75), .A3(G86), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n514), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n529), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n583), .B2(new_n582), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n539), .A2(G85), .B1(new_n541), .B2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n505), .A2(new_n506), .A3(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT77), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n509), .B2(KEYINPUT78), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n514), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n594), .A2(new_n596), .B1(new_n599), .B2(G651), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n592), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n592), .A2(new_n593), .A3(new_n600), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n589), .B1(new_n606), .B2(new_n588), .ZN(G284));
  AOI21_X1  g182(.A(new_n589), .B1(new_n606), .B2(new_n588), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n562), .ZN(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G860), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g189(.A1(new_n543), .A2(new_n544), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n588), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n602), .A2(new_n612), .A3(new_n605), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n588), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n462), .A2(new_n469), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n481), .A2(G123), .B1(G135), .B2(new_n468), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n628), .A2(KEYINPUT83), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(KEYINPUT83), .B2(new_n628), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT84), .Z(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(G401));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n444), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT17), .Z(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  INV_X1    g235(.A(new_n653), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n656), .C1(new_n661), .C2(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n655), .A3(new_n657), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT32), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(G288), .A2(KEYINPUT91), .ZN(new_n690));
  NAND2_X1  g265(.A1(G288), .A2(KEYINPUT91), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G23), .B(new_n692), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT92), .Z(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G1971), .Z(new_n700));
  NAND3_X1  g275(.A1(new_n689), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n481), .A2(G119), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n468), .A2(G131), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n464), .A2(G107), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n709), .S(G29), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT87), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT88), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n710), .B(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G24), .B(G290), .S(G16), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n716), .B2(KEYINPUT89), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(KEYINPUT89), .B2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n703), .A2(new_n704), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT36), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n696), .A2(G20), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT23), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n562), .B2(new_n696), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1956), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT96), .B(G1966), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n696), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n696), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT95), .Z(new_n729));
  AOI21_X1  g304(.A(new_n724), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G1341), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n545), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G16), .B2(G19), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n730), .B1(new_n731), .B2(new_n733), .C1(new_n726), .C2(new_n729), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT30), .B(G28), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n632), .B2(new_n736), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n468), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n742), .B(new_n744), .C1(G129), .C2(new_n481), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n736), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n736), .B2(G32), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n736), .A2(G33), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n751));
  NAND2_X1  g326(.A1(G103), .A2(G2104), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(G2105), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n468), .A2(G139), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n464), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n442), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n481), .A2(G128), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n468), .A2(G140), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n464), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n736), .A2(G26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT93), .B(G2067), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n749), .A2(new_n760), .A3(new_n761), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n696), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n696), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n778), .B2(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT24), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n471), .B2(new_n736), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G2084), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n777), .B(new_n783), .C1(new_n747), .C2(new_n748), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n736), .A2(G27), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n736), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n758), .A2(new_n442), .B1(new_n787), .B2(G2078), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n788), .B1(G2078), .B2(new_n787), .C1(new_n782), .C2(G2084), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n734), .A2(new_n773), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n736), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n736), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT29), .Z(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n733), .A2(new_n731), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n790), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n696), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n606), .B2(new_n696), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n720), .A2(new_n798), .A3(new_n801), .ZN(G311));
  INV_X1    g377(.A(G311), .ZN(G150));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  INV_X1    g379(.A(G55), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n507), .A2(new_n804), .B1(new_n509), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n529), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT99), .B(G860), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n606), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n545), .B(new_n809), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT39), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(new_n810), .ZN(G145));
  XNOR2_X1  g394(.A(new_n745), .B(new_n757), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n709), .B(new_n622), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n494), .A2(new_n499), .ZN(new_n823));
  INV_X1    g398(.A(new_n488), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n766), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n481), .A2(G130), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n464), .A2(G118), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G142), .B2(new_n468), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n822), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(G162), .B(new_n471), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n632), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT101), .B(G37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g414(.A(G303), .B(G305), .Z(new_n840));
  XOR2_X1   g415(.A(new_n692), .B(G290), .Z(new_n841));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n809), .B(new_n615), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n617), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n603), .B(G299), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n603), .B(new_n562), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT41), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n847), .A2(new_n850), .A3(new_n848), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n858), .B1(new_n857), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n845), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT42), .ZN(new_n865));
  INV_X1    g440(.A(new_n845), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n588), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n809), .A2(new_n588), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT103), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n861), .A2(new_n845), .A3(new_n862), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n866), .B1(new_n865), .B2(new_n860), .ZN(new_n873));
  OAI21_X1  g448(.A(G868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n876), .ZN(G295));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n869), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n879));
  XNOR2_X1  g454(.A(G171), .B(G168), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n816), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n846), .A2(new_n880), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n846), .A2(KEYINPUT105), .A3(new_n880), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n850), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(KEYINPUT104), .A3(new_n884), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n846), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n855), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n845), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n891), .A2(new_n845), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n879), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n837), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n891), .B2(new_n845), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n855), .A2(new_n886), .A3(new_n885), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n888), .A2(new_n889), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n853), .ZN(new_n901));
  AOI211_X1 g476(.A(KEYINPUT106), .B(new_n845), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n899), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n866), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n898), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n896), .B1(new_n879), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n894), .B2(new_n895), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(KEYINPUT43), .B2(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(G397));
  XNOR2_X1  g488(.A(KEYINPUT107), .B(G1384), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n825), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n465), .A2(G40), .A3(new_n470), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n766), .B(G2067), .Z(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n745), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT124), .Z(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT46), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT47), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n919), .A2(new_n924), .A3(new_n745), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT108), .Z(new_n930));
  OAI21_X1  g505(.A(new_n921), .B1(new_n924), .B2(new_n745), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n919), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n709), .B(new_n712), .Z(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n920), .A2(G1986), .A3(G290), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT126), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n928), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n709), .A2(new_n712), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G2067), .B2(new_n766), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n920), .B1(new_n942), .B2(KEYINPUT123), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT122), .ZN(new_n946));
  INV_X1    g521(.A(G48), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n570), .B1(new_n947), .B2(new_n509), .ZN(new_n948));
  OAI21_X1  g523(.A(G1981), .B1(new_n948), .B2(new_n576), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n572), .A2(new_n577), .A3(new_n688), .A4(new_n578), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(G1981), .C1(new_n948), .C2(new_n576), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n950), .A2(KEYINPUT49), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n465), .A2(G40), .A3(new_n470), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(G164), .B2(G1384), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n495), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n462), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n490), .A2(new_n498), .A3(G138), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n491), .A2(new_n960), .B1(new_n961), .B2(new_n468), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n957), .B(new_n958), .C1(new_n962), .C2(new_n488), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n956), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT49), .B1(new_n967), .B2(KEYINPUT112), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n950), .A2(new_n970), .A3(new_n951), .A4(new_n953), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n954), .B(new_n966), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(G288), .A2(G1976), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT114), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n951), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n966), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n690), .A2(G1976), .A3(new_n691), .ZN(new_n980));
  INV_X1    g555(.A(G1976), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(G288), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n966), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(G8), .A3(new_n964), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT52), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n825), .A2(new_n958), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n918), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n956), .A2(new_n963), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n992), .B(new_n794), .C1(new_n993), .C2(KEYINPUT50), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n916), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n825), .A2(KEYINPUT45), .A3(new_n914), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n955), .A3(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(KEYINPUT109), .B(G1971), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n990), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n974), .A2(new_n986), .A3(new_n989), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n979), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n989), .A2(new_n1000), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT63), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n989), .B2(new_n1000), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n974), .A3(new_n1005), .A4(new_n986), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n991), .A2(new_n916), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n918), .B1(new_n993), .B2(new_n916), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n956), .B2(new_n963), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n1011), .B2(new_n918), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n726), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n992), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(G2084), .ZN(new_n1015));
  OAI211_X1 g590(.A(G8), .B(G168), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n987), .B(KEYINPUT55), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n955), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n956), .B2(new_n963), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1022), .A2(new_n794), .B1(new_n998), .B2(new_n997), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1018), .B1(new_n1023), .B2(new_n990), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n989), .A2(new_n1000), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n974), .A2(new_n1024), .A3(new_n986), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1004), .B1(new_n1026), .B2(new_n1016), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1017), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT116), .B(new_n1004), .C1(new_n1026), .C2(new_n1016), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1002), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1010), .A2(new_n1012), .A3(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n995), .A2(new_n955), .A3(new_n996), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n443), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1036), .A2(new_n1032), .B1(new_n776), .B2(new_n1014), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G171), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G168), .A2(new_n990), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(KEYINPUT120), .B2(KEYINPUT51), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n957), .B1(new_n825), .B2(new_n958), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT110), .B(G1384), .C1(new_n823), .C2(new_n824), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n916), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n1009), .A3(new_n955), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1007), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1012), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1015), .B1(new_n1048), .B2(new_n725), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1042), .B1(new_n1049), .B2(new_n990), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1016), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n725), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1015), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n990), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1040), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1051), .B1(new_n1056), .B2(KEYINPUT51), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1039), .B1(new_n1057), .B2(KEYINPUT62), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1051), .C1(new_n1056), .C2(KEYINPUT51), .ZN(new_n1060));
  XNOR2_X1  g635(.A(G171), .B(KEYINPUT54), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1038), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n917), .A2(new_n1064), .A3(new_n955), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n917), .B2(new_n955), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n996), .B(new_n1033), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1037), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  AOI22_X1  g646(.A1(new_n1035), .A2(new_n924), .B1(new_n964), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n1072), .A2(new_n615), .B1(KEYINPUT119), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1014), .A2(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n964), .A2(G2067), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n603), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n964), .A2(new_n1071), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n997), .B2(G1996), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1073), .A2(KEYINPUT119), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n545), .A3(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1074), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n562), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1035), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1095), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1093), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1077), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n601), .A3(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1083), .A2(new_n1096), .A3(new_n1099), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n603), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1095), .B1(new_n1106), .B2(new_n1093), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(new_n1095), .C1(new_n1106), .C2(new_n1093), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1070), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1058), .A2(new_n1060), .B1(new_n1057), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1031), .B1(new_n1113), .B2(new_n1026), .ZN(new_n1114));
  XNOR2_X1  g689(.A(G290), .B(G1986), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n934), .B1(new_n919), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n946), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1050), .A2(new_n1016), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1055), .B(G8), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT51), .B1(new_n1119), .B2(new_n1041), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1039), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1060), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1112), .A2(new_n1057), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1026), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1017), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1030), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1002), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n946), .B(new_n1116), .C1(new_n1125), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n945), .B1(new_n1117), .B2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g708(.A(G319), .ZN(new_n1135));
  NOR3_X1   g709(.A1(G227), .A2(new_n650), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g710(.A1(new_n684), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g711(.A(new_n1137), .B(KEYINPUT127), .ZN(new_n1138));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n838), .A3(new_n1138), .ZN(G225));
  INV_X1    g713(.A(G225), .ZN(G308));
endmodule


