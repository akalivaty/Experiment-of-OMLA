//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1287, new_n1288,
    new_n1289;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT68), .B1(new_n469), .B2(G101), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI22_X1  g048(.A1(new_n467), .A2(new_n468), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n476), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G138), .B(new_n466), .C1(new_n475), .C2(new_n476), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n492), .A3(G138), .A4(new_n466), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n466), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n498), .A2(new_n502), .B1(new_n484), .B2(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  AND2_X1   g081(.A1(G75), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n507), .B1(new_n514), .B2(G62), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n518), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .A3(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(new_n521), .B1(KEYINPUT6), .B2(new_n516), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(new_n514), .A3(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G50), .A3(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  AOI211_X1 g101(.A(new_n526), .B(new_n509), .C1(new_n511), .C2(new_n513), .ZN(new_n527));
  OAI211_X1 g102(.A(KEYINPUT72), .B(G651), .C1(new_n527), .C2(new_n507), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n517), .A2(new_n525), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n522), .A2(new_n514), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n522), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n514), .A2(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n522), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n531), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n516), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n531), .A2(new_n550), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n516), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n514), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g137(.A(KEYINPUT73), .B(new_n509), .C1(new_n511), .C2(new_n513), .ZN(new_n563));
  OAI21_X1  g138(.A(G65), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n516), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n519), .A2(new_n521), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n567), .A2(G53), .A3(G543), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n522), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n532), .A2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  NAND3_X1  g153(.A1(new_n522), .A2(new_n514), .A3(G87), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n522), .A2(G49), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g159(.A(KEYINPUT74), .B(G651), .C1(new_n514), .C2(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  INV_X1    g162(.A(new_n509), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n512), .B1(KEYINPUT5), .B2(new_n508), .ZN(new_n589));
  NOR3_X1   g164(.A1(new_n510), .A2(KEYINPUT71), .A3(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(G61), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n514), .A2(KEYINPUT75), .A3(G61), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  INV_X1    g173(.A(G48), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n531), .A2(new_n598), .B1(new_n544), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n531), .A2(new_n603), .B1(new_n544), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n516), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G171), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT76), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n522), .A2(new_n514), .A3(G92), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n534), .A2(G54), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT73), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n514), .A2(new_n561), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G66), .ZN(new_n624));
  NAND2_X1  g199(.A1(G79), .A2(G543), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n516), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n612), .B1(G868), .B2(new_n627), .ZN(G284));
  OAI21_X1  g203(.A(new_n612), .B1(G868), .B2(new_n627), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n576), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n576), .B2(G868), .ZN(G280));
  XNOR2_X1  g207(.A(KEYINPUT78), .B(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n627), .B1(G860), .B2(new_n633), .ZN(G148));
  OAI21_X1  g209(.A(KEYINPUT80), .B1(new_n555), .B2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n624), .A2(new_n625), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G651), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n615), .A2(new_n616), .B1(G54), .B2(new_n534), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(new_n638), .A3(new_n633), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G868), .ZN(new_n644));
  MUX2_X1   g219(.A(KEYINPUT80), .B(new_n635), .S(new_n644), .Z(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n465), .A2(new_n469), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT13), .Z(new_n649));
  INV_X1    g224(.A(G2100), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n484), .A2(G123), .ZN(new_n653));
  OR2_X1    g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n655));
  INV_X1    g230(.A(G135), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n655), .C1(new_n656), .C2(new_n467), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(G2096), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n652), .A3(new_n658), .ZN(G156));
  INV_X1    g234(.A(G14), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n660), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n673), .B(KEYINPUT81), .C1(new_n672), .C2(new_n671), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n675));
  INV_X1    g250(.A(new_n669), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n668), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n666), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n672), .ZN(new_n679));
  OAI21_X1  g254(.A(G14), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n671), .A2(new_n672), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n674), .A2(new_n682), .ZN(G401));
  XOR2_X1   g258(.A(G2067), .B(G2678), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT82), .ZN(new_n685));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  XNOR2_X1  g261(.A(G2084), .B(G2090), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT18), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(KEYINPUT17), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n687), .C1(new_n685), .C2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n687), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n691), .A2(new_n685), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G2096), .B(G2100), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n689), .A2(new_n692), .A3(new_n694), .A4(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(G227));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1956), .B(G2474), .Z(new_n706));
  XOR2_X1   g281(.A(G1961), .B(G1966), .Z(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT20), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  OR3_X1    g287(.A1(new_n705), .A2(new_n708), .A3(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n709), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n713), .A2(new_n712), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(new_n715), .ZN(new_n722));
  XOR2_X1   g297(.A(G1991), .B(G1996), .Z(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AND3_X1   g299(.A1(new_n717), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n717), .B2(new_n722), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n702), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n714), .A2(new_n716), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n721), .A2(new_n715), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n717), .A2(new_n722), .A3(new_n724), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n730), .A2(new_n701), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(G229));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G25), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G131), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT83), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n740));
  INV_X1    g315(.A(G107), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G2105), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G119), .B2(new_n484), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n737), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n608), .B2(new_n751), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G1986), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(G1986), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n749), .A2(new_n750), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n586), .A2(new_n751), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n751), .B2(G23), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT33), .B(G1976), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G166), .A2(G16), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G1971), .C1(G16), .C2(G22), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(G16), .B2(G22), .ZN(new_n763));
  INV_X1    g338(.A(G1971), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n758), .A2(new_n759), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n760), .A2(new_n762), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n597), .A2(new_n601), .A3(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G6), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT32), .B(G1981), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n768), .B(new_n770), .C1(G6), .C2(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT85), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n767), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT34), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n756), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n760), .A2(new_n765), .A3(new_n766), .ZN(new_n784));
  INV_X1    g359(.A(new_n778), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n784), .A2(new_n785), .A3(new_n776), .A4(new_n762), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n786), .A2(KEYINPUT86), .A3(KEYINPUT34), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n781), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n488), .A2(G29), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n735), .A2(G35), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2090), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n798), .A2(KEYINPUT97), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT97), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n751), .A2(G20), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT23), .Z(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G299), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT98), .B(G1956), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(G164), .A2(G29), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G27), .B2(G29), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT96), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT96), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n443), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(G2078), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n802), .B(new_n807), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n735), .A2(G32), .ZN(new_n816));
  NAND3_X1  g391(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT26), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G129), .B2(new_n484), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n816), .B1(new_n822), .B2(new_n735), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT27), .B(G1996), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n735), .A2(G33), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n465), .A2(G127), .ZN(new_n827));
  AND2_X1   g402(.A1(G115), .A2(G2104), .ZN(new_n828));
  OAI21_X1  g403(.A(G2105), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n830));
  NAND2_X1  g405(.A1(G103), .A2(G2104), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G2105), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n482), .A2(G139), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n826), .B1(new_n835), .B2(new_n735), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n442), .ZN(new_n837));
  INV_X1    g412(.A(G34), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT24), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(KEYINPUT24), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n735), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G160), .B2(new_n735), .ZN(new_n842));
  INV_X1    g417(.A(G2084), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n825), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n751), .A2(G19), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n555), .B2(new_n751), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(G1341), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n798), .A2(new_n799), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n484), .A2(G128), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT89), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(G116), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(G2105), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n482), .B2(G140), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G29), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n735), .A2(G26), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT28), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G2067), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(G2067), .A3(new_n859), .ZN(new_n863));
  NOR2_X1   g438(.A1(G5), .A2(G16), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT93), .Z(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(G301), .B2(new_n751), .ZN(new_n866));
  INV_X1    g441(.A(G1961), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n862), .A2(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n845), .A2(new_n848), .A3(new_n849), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n627), .A2(G16), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(G4), .B2(G16), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT88), .B(G1348), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n815), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n751), .A2(G21), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G168), .B2(new_n751), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT90), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G1966), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n866), .A2(new_n880), .A3(new_n867), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n866), .B2(new_n867), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT31), .B(G11), .ZN(new_n884));
  XOR2_X1   g459(.A(KEYINPUT30), .B(G28), .Z(new_n885));
  NOR2_X1   g460(.A1(new_n657), .A2(new_n735), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n884), .B1(G29), .B2(new_n885), .C1(new_n886), .C2(KEYINPUT91), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(KEYINPUT91), .B2(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT90), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n877), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G1966), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT92), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT92), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n878), .A2(new_n895), .A3(G1966), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n890), .B(KEYINPUT95), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n889), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n875), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n781), .A2(new_n783), .A3(new_n787), .A4(new_n790), .ZN(new_n903));
  AND4_X1   g478(.A1(KEYINPUT99), .A2(new_n793), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n788), .B2(new_n792), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT99), .B1(new_n905), .B2(new_n903), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(G311));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n903), .ZN(G150));
  INV_X1    g483(.A(G93), .ZN(new_n909));
  INV_X1    g484(.A(G55), .ZN(new_n910));
  OAI22_X1  g485(.A1(new_n531), .A2(new_n909), .B1(new_n544), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n516), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G860), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT37), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n627), .A2(G559), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT38), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n552), .A2(new_n554), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n914), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n911), .A2(new_n913), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n555), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n918), .B(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT39), .ZN(new_n925));
  AOI21_X1  g500(.A(G860), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n916), .B1(new_n929), .B2(new_n930), .ZN(G145));
  XNOR2_X1  g506(.A(KEYINPUT102), .B(G37), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n744), .A2(new_n648), .ZN(new_n933));
  INV_X1    g508(.A(new_n648), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n739), .A3(new_n743), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n835), .B(new_n821), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n822), .B(new_n835), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n933), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n856), .A2(new_n504), .ZN(new_n942));
  NAND3_X1  g517(.A1(G164), .A2(new_n851), .A3(new_n855), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n484), .A2(G130), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT101), .Z(new_n946));
  OAI21_X1  g521(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n947));
  INV_X1    g522(.A(G118), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(G2105), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n482), .A2(G142), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n944), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n952), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n488), .B(new_n657), .Z(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(G160), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n953), .A2(new_n938), .A3(new_n940), .A4(new_n954), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n956), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n932), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT103), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n932), .C1(new_n962), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g544(.A(G305), .B(new_n608), .ZN(new_n970));
  XNOR2_X1  g545(.A(G303), .B(new_n586), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n970), .B(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n637), .A2(new_n638), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(G299), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n627), .A2(new_n576), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n920), .A2(new_n922), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n641), .A2(new_n642), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n641), .B2(new_n642), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n981), .A2(KEYINPUT41), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n979), .B2(new_n980), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n643), .A2(new_n923), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n983), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n976), .B1(new_n977), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n974), .A2(new_n986), .A3(new_n992), .A4(new_n975), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G868), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n921), .A2(G868), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(G295));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1001), .A3(new_n999), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n610), .B1(new_n994), .B2(new_n995), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT106), .B1(new_n1003), .B2(new_n998), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(G331));
  NAND2_X1  g580(.A1(new_n982), .A2(G301), .ZN(new_n1006));
  AOI21_X1  g581(.A(G301), .B1(new_n920), .B2(new_n922), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(G168), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n923), .A2(G171), .ZN(new_n1010));
  OAI21_X1  g585(.A(G286), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT41), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n981), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n981), .B2(new_n988), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n972), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1009), .B(new_n1011), .C1(new_n987), .C2(new_n989), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n972), .A3(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n932), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G37), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n972), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT43), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1020), .A2(new_n932), .A3(new_n1023), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1021), .ZN(new_n1032));
  MUX2_X1   g607(.A(new_n1029), .B(new_n1032), .S(KEYINPUT44), .Z(G397));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n504), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n471), .A2(new_n472), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n469), .A2(KEYINPUT68), .A3(G101), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n482), .A2(G137), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n479), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(G40), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT108), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n856), .B(new_n861), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n821), .B2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1037), .A2(G1996), .A3(new_n1042), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT107), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1047), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT47), .ZN(new_n1054));
  INV_X1    g629(.A(G1996), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1045), .B1(new_n1055), .B2(new_n822), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1049), .A2(new_n822), .B1(new_n1044), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n746), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n748), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n856), .A2(G2067), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1044), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR4_X1   g636(.A1(G290), .A2(new_n1037), .A3(G1986), .A4(new_n1042), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n1062), .B(KEYINPUT48), .Z(new_n1063));
  XOR2_X1   g638(.A(new_n744), .B(new_n748), .Z(new_n1064));
  NAND2_X1  g639(.A1(new_n1044), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1054), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT45), .B1(new_n504), .B2(new_n1034), .ZN(new_n1068));
  AOI211_X1 g643(.A(new_n1036), .B(G1384), .C1(new_n494), .C2(new_n503), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G40), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n474), .A2(new_n1071), .A3(new_n479), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(new_n442), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1384), .B1(new_n494), .B2(new_n503), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n504), .A2(new_n1077), .A3(new_n1034), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(KEYINPUT114), .A3(new_n1077), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1075), .B1(new_n1083), .B2(G1956), .ZN(new_n1084));
  INV_X1    g659(.A(G65), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n621), .B2(new_n622), .ZN(new_n1086));
  INV_X1    g661(.A(new_n565), .ZN(new_n1087));
  OAI21_X1  g662(.A(G651), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n570), .A2(new_n572), .B1(new_n532), .B2(G91), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT115), .B1(new_n570), .B2(new_n572), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1088), .B(new_n1089), .C1(KEYINPUT57), .C2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(KEYINPUT57), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n566), .B2(new_n575), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1094), .B(new_n1075), .C1(G1956), .C2(new_n1083), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT61), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n623), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n638), .B(KEYINPUT60), .C1(new_n1099), .C2(new_n516), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT121), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n637), .A2(new_n1102), .A3(KEYINPUT60), .A4(new_n638), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n619), .B2(new_n626), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n861), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1079), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1078), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1106), .B(new_n1109), .C1(G1348), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1042), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1079), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1115), .A2(new_n1116), .B1(new_n861), .B2(new_n1108), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(new_n1103), .A3(new_n1101), .A4(new_n1106), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1098), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1097), .B2(KEYINPUT120), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1082), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT114), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1114), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1956), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1068), .A2(new_n1069), .A3(new_n1042), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1125), .A2(new_n1126), .B1(new_n1127), .B2(new_n1074), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT117), .B1(new_n1128), .B2(new_n1094), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1084), .A2(new_n1130), .A3(new_n1095), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1132), .A3(new_n1094), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1122), .A2(new_n1129), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1076), .A2(KEYINPUT45), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1042), .A2(G1996), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1037), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1107), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1137), .A2(KEYINPUT118), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT118), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n555), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT119), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n555), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT59), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(KEYINPUT119), .A3(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1120), .A2(new_n1134), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1129), .B(new_n1131), .C1(new_n978), .C2(new_n1117), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1097), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1037), .A2(new_n1072), .A3(new_n1135), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n893), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(new_n843), .A3(new_n1072), .A4(new_n1079), .ZN(new_n1157));
  NAND2_X1  g732(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT51), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1161));
  OAI211_X1 g736(.A(G8), .B(new_n1160), .C1(new_n1161), .C2(G286), .ZN(new_n1162));
  OAI211_X1 g737(.A(G168), .B(new_n1157), .C1(new_n1127), .C2(G1966), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(G8), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1159), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT110), .B(G2090), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1114), .A2(new_n1079), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1127), .B2(G1971), .ZN(new_n1169));
  NAND2_X1  g744(.A1(G303), .A2(G8), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT55), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1169), .A2(G8), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT111), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G8), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1154), .A2(new_n764), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1178), .B1(new_n1179), .B2(new_n1168), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(KEYINPUT111), .A3(new_n1174), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1178), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n584), .A2(new_n585), .ZN(new_n1184));
  INV_X1    g759(.A(new_n581), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(G1976), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT112), .B1(new_n1187), .B2(KEYINPUT52), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT112), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT52), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1189), .B(new_n1190), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n586), .B2(G1976), .ZN(new_n1192));
  OAI22_X1  g767(.A1(new_n1188), .A2(new_n1191), .B1(new_n1187), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(G1981), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n597), .A2(new_n601), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n595), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1196), .B1(new_n591), .B2(new_n592), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n516), .B1(new_n1197), .B2(new_n594), .ZN(new_n1198));
  OAI21_X1  g773(.A(G1981), .B1(new_n1198), .B2(new_n600), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1195), .A2(new_n1199), .A3(KEYINPUT49), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT113), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT113), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1195), .A2(new_n1199), .A3(new_n1202), .A4(KEYINPUT49), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT49), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1183), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1193), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g783(.A1(new_n1083), .A2(new_n1167), .B1(new_n1154), .B2(new_n764), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1172), .B(new_n1173), .C1(new_n1209), .C2(new_n1178), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1166), .A2(new_n1182), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1037), .A2(new_n443), .A3(new_n1072), .A4(new_n1135), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT53), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1070), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1072), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n867), .B1(new_n1078), .B2(new_n1110), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1217), .A2(G171), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT54), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1214), .A2(new_n1215), .A3(G301), .A4(new_n1216), .ZN(new_n1220));
  AND3_X1   g795(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1219), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1153), .B1(new_n1211), .B2(new_n1223), .ZN(new_n1224));
  AND4_X1   g799(.A1(KEYINPUT111), .A2(new_n1169), .A3(G8), .A4(new_n1174), .ZN(new_n1225));
  AOI21_X1  g800(.A(KEYINPUT111), .B1(new_n1180), .B2(new_n1174), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1187), .A2(KEYINPUT52), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1189), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1187), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1229), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1210), .A2(new_n1228), .A3(new_n1233), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g810(.A1(new_n867), .A2(new_n1115), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1236));
  AOI21_X1  g811(.A(G301), .B1(new_n1236), .B2(new_n1215), .ZN(new_n1237));
  INV_X1    g812(.A(new_n1220), .ZN(new_n1238));
  OAI21_X1  g813(.A(KEYINPUT54), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g816(.A1(new_n1235), .A2(KEYINPUT123), .A3(new_n1241), .A4(new_n1166), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1152), .A2(new_n1224), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1228), .A2(new_n1233), .ZN(new_n1244));
  NAND2_X1  g819(.A1(G168), .A2(G8), .ZN(new_n1245));
  AOI21_X1  g820(.A(new_n1245), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1246), .B1(new_n1180), .B2(new_n1174), .ZN(new_n1247));
  OAI21_X1  g822(.A(KEYINPUT63), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  OR2_X1    g823(.A1(G288), .A2(G1976), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1249), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1250));
  INV_X1    g825(.A(new_n1195), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1183), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  AOI211_X1 g827(.A(KEYINPUT63), .B(new_n1245), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1253));
  AOI22_X1  g828(.A1(new_n1177), .A2(new_n1181), .B1(new_n1210), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g829(.A(new_n1248), .B(new_n1252), .C1(new_n1254), .C2(new_n1244), .ZN(new_n1255));
  INV_X1    g830(.A(KEYINPUT124), .ZN(new_n1256));
  AOI21_X1  g831(.A(new_n1256), .B1(new_n1166), .B2(KEYINPUT62), .ZN(new_n1257));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1258));
  NAND3_X1  g833(.A1(new_n1162), .A2(new_n1258), .A3(new_n1165), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1259), .A2(new_n1237), .ZN(new_n1260));
  NOR2_X1   g835(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g836(.A(KEYINPUT124), .B(new_n1258), .C1(new_n1162), .C2(new_n1165), .ZN(new_n1262));
  NAND3_X1  g837(.A1(new_n1182), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1263));
  NOR2_X1   g838(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g839(.A(new_n1255), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1243), .A2(new_n1265), .ZN(new_n1266));
  XOR2_X1   g841(.A(new_n608), .B(G1986), .Z(new_n1267));
  NAND2_X1  g842(.A1(new_n1267), .A2(new_n1043), .ZN(new_n1268));
  NAND3_X1  g843(.A1(new_n1057), .A2(new_n1268), .A3(new_n1065), .ZN(new_n1269));
  XNOR2_X1  g844(.A(new_n1269), .B(KEYINPUT109), .ZN(new_n1270));
  INV_X1    g845(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g846(.A(KEYINPUT125), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g847(.A(KEYINPUT125), .ZN(new_n1273));
  AOI211_X1 g848(.A(new_n1273), .B(new_n1270), .C1(new_n1243), .C2(new_n1265), .ZN(new_n1274));
  OAI21_X1  g849(.A(new_n1067), .B1(new_n1272), .B2(new_n1274), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g850(.A1(new_n698), .A2(G319), .A3(new_n699), .ZN(new_n1277));
  AOI21_X1  g851(.A(new_n1277), .B1(new_n674), .B2(new_n682), .ZN(new_n1278));
  AND3_X1   g852(.A1(new_n733), .A2(new_n1278), .A3(KEYINPUT126), .ZN(new_n1279));
  AOI21_X1  g853(.A(KEYINPUT126), .B1(new_n733), .B2(new_n1278), .ZN(new_n1280));
  NOR2_X1   g854(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g855(.A(new_n1281), .B1(new_n965), .B2(new_n967), .ZN(new_n1282));
  INV_X1    g856(.A(KEYINPUT127), .ZN(new_n1283));
  AND3_X1   g857(.A1(new_n1029), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g858(.A(new_n1283), .B1(new_n1029), .B2(new_n1282), .ZN(new_n1285));
  NOR2_X1   g859(.A1(new_n1284), .A2(new_n1285), .ZN(G308));
  NAND2_X1  g860(.A1(new_n1029), .A2(new_n1282), .ZN(new_n1287));
  NAND2_X1  g861(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1288));
  NAND3_X1  g862(.A1(new_n1029), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1289));
  NAND2_X1  g863(.A1(new_n1288), .A2(new_n1289), .ZN(G225));
endmodule


