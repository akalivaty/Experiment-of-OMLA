

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n366, n367, n368, n369, n370, n371, n372,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748;

  BUF_X1 U372 ( .A(n677), .Z(n350) );
  AND2_X1 U373 ( .A1(n658), .A2(n428), .ZN(n551) );
  NOR2_X1 U374 ( .A1(n535), .A2(n572), .ZN(n525) );
  XNOR2_X1 U375 ( .A(n351), .B(KEYINPUT19), .ZN(n584) );
  NAND2_X1 U376 ( .A1(n427), .A2(n631), .ZN(n351) );
  XNOR2_X1 U377 ( .A(n353), .B(G122), .ZN(n491) );
  INV_X2 U378 ( .A(G107), .ZN(n353) );
  NOR2_X1 U379 ( .A1(n352), .A2(n673), .ZN(n530) );
  NOR2_X1 U380 ( .A1(n528), .A2(n527), .ZN(n352) );
  XNOR2_X2 U381 ( .A(n730), .B(n499), .ZN(n655) );
  XNOR2_X2 U382 ( .A(n435), .B(n492), .ZN(n730) );
  XNOR2_X1 U383 ( .A(G113), .B(G122), .ZN(n465) );
  INV_X2 U384 ( .A(G104), .ZN(n382) );
  AND2_X2 U385 ( .A1(n632), .A2(n631), .ZN(n568) );
  XNOR2_X2 U386 ( .A(n578), .B(KEYINPUT38), .ZN(n632) );
  XNOR2_X2 U387 ( .A(n510), .B(KEYINPUT0), .ZN(n535) );
  NOR2_X2 U388 ( .A1(n748), .A2(n747), .ZN(n577) );
  NOR2_X1 U389 ( .A1(n374), .A2(n570), .ZN(n677) );
  AND2_X2 U390 ( .A1(n404), .A2(n664), .ZN(n716) );
  NAND2_X1 U391 ( .A1(n663), .A2(n662), .ZN(n404) );
  AND2_X1 U392 ( .A1(n590), .A2(n589), .ZN(n603) );
  XNOR2_X1 U393 ( .A(n540), .B(n539), .ZN(n744) );
  NOR2_X1 U394 ( .A1(n677), .A2(n695), .ZN(n385) );
  XNOR2_X1 U395 ( .A(n377), .B(n376), .ZN(n650) );
  XNOR2_X1 U396 ( .A(n571), .B(n383), .ZN(n424) );
  INV_X1 U397 ( .A(n570), .ZN(n620) );
  INV_X1 U398 ( .A(n450), .ZN(n570) );
  XNOR2_X1 U399 ( .A(n426), .B(n425), .ZN(n552) );
  OR2_X1 U400 ( .A1(n718), .A2(G902), .ZN(n426) );
  XNOR2_X1 U401 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U402 ( .A(n461), .B(n460), .ZN(n718) );
  XNOR2_X1 U403 ( .A(n381), .B(n490), .ZN(n514) );
  XNOR2_X1 U404 ( .A(n382), .B(G110), .ZN(n381) );
  XNOR2_X1 U405 ( .A(n392), .B(G143), .ZN(n494) );
  INV_X1 U406 ( .A(KEYINPUT93), .ZN(n384) );
  XNOR2_X1 U407 ( .A(n494), .B(n439), .ZN(n482) );
  INV_X1 U408 ( .A(G134), .ZN(n439) );
  NAND2_X1 U409 ( .A1(n744), .A2(n549), .ZN(n400) );
  NOR2_X1 U410 ( .A1(n746), .A2(n390), .ZN(n549) );
  XNOR2_X1 U411 ( .A(n380), .B(n482), .ZN(n734) );
  XNOR2_X1 U412 ( .A(n524), .B(KEYINPUT1), .ZN(n621) );
  NOR2_X1 U413 ( .A1(n522), .A2(n552), .ZN(n622) );
  XNOR2_X1 U414 ( .A(KEYINPUT6), .B(KEYINPUT99), .ZN(n451) );
  XNOR2_X1 U415 ( .A(n447), .B(n446), .ZN(n492) );
  INV_X1 U416 ( .A(G119), .ZN(n446) );
  NAND2_X1 U417 ( .A1(n613), .A2(n614), .ZN(n664) );
  XNOR2_X1 U418 ( .A(n415), .B(n414), .ZN(n733) );
  INV_X1 U419 ( .A(KEYINPUT10), .ZN(n414) );
  XNOR2_X1 U420 ( .A(G140), .B(G125), .ZN(n415) );
  XOR2_X1 U421 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n456) );
  NAND2_X1 U422 ( .A1(n621), .A2(n622), .ZN(n532) );
  XNOR2_X1 U423 ( .A(n400), .B(n399), .ZN(n398) );
  XOR2_X1 U424 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n453) );
  XNOR2_X1 U425 ( .A(G110), .B(G128), .ZN(n452) );
  XNOR2_X1 U426 ( .A(G119), .B(G137), .ZN(n457) );
  XNOR2_X1 U427 ( .A(n733), .B(n413), .ZN(n474) );
  INV_X1 U428 ( .A(G146), .ZN(n413) );
  XNOR2_X1 U429 ( .A(n514), .B(n372), .ZN(n517) );
  XNOR2_X1 U430 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U431 ( .A(n494), .B(n393), .ZN(n498) );
  NAND2_X1 U432 ( .A1(n572), .A2(n422), .ZN(n421) );
  AND2_X1 U433 ( .A1(n421), .A2(n419), .ZN(n378) );
  NAND2_X1 U434 ( .A1(n354), .A2(n369), .ZN(n418) );
  AND2_X1 U435 ( .A1(n370), .A2(n424), .ZN(n369) );
  INV_X1 U436 ( .A(n572), .ZN(n370) );
  BUF_X1 U437 ( .A(n621), .Z(n386) );
  NOR2_X1 U438 ( .A1(n560), .A2(n559), .ZN(n594) );
  INV_X1 U439 ( .A(n621), .ZN(n543) );
  XNOR2_X1 U440 ( .A(n366), .B(KEYINPUT22), .ZN(n547) );
  XNOR2_X1 U441 ( .A(n464), .B(KEYINPUT25), .ZN(n425) );
  XNOR2_X1 U442 ( .A(n412), .B(n669), .ZN(n411) );
  INV_X1 U443 ( .A(G953), .ZN(n737) );
  XNOR2_X1 U444 ( .A(n396), .B(G146), .ZN(n493) );
  INV_X1 U445 ( .A(KEYINPUT4), .ZN(n396) );
  INV_X1 U446 ( .A(KEYINPUT48), .ZN(n604) );
  XNOR2_X1 U447 ( .A(KEYINPUT67), .B(G469), .ZN(n519) );
  XNOR2_X1 U448 ( .A(KEYINPUT3), .B(G116), .ZN(n443) );
  INV_X1 U449 ( .A(KEYINPUT44), .ZN(n399) );
  INV_X1 U450 ( .A(KEYINPUT101), .ZN(n402) );
  XNOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  XNOR2_X1 U452 ( .A(G131), .B(KEYINPUT11), .ZN(n467) );
  XOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT94), .Z(n468) );
  XOR2_X1 U454 ( .A(G143), .B(G104), .Z(n466) );
  XNOR2_X1 U455 ( .A(n513), .B(n515), .ZN(n372) );
  INV_X1 U456 ( .A(G140), .ZN(n515) );
  XOR2_X1 U457 ( .A(G101), .B(G107), .Z(n513) );
  XNOR2_X1 U458 ( .A(n493), .B(n394), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n395), .B(G125), .ZN(n394) );
  INV_X1 U460 ( .A(KEYINPUT18), .ZN(n395) );
  XNOR2_X1 U461 ( .A(G128), .B(KEYINPUT64), .ZN(n392) );
  INV_X1 U462 ( .A(KEYINPUT17), .ZN(n495) );
  XNOR2_X1 U463 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n607) );
  INV_X1 U464 ( .A(KEYINPUT30), .ZN(n383) );
  NAND2_X1 U465 ( .A1(n570), .A2(n631), .ZN(n571) );
  XNOR2_X1 U466 ( .A(n438), .B(n734), .ZN(n668) );
  XNOR2_X1 U467 ( .A(n492), .B(n375), .ZN(n438) );
  XNOR2_X1 U468 ( .A(n442), .B(n448), .ZN(n375) );
  NOR2_X1 U469 ( .A1(n660), .A2(n658), .ZN(n659) );
  XNOR2_X1 U470 ( .A(n482), .B(n379), .ZN(n483) );
  XNOR2_X1 U471 ( .A(n491), .B(KEYINPUT97), .ZN(n379) );
  XNOR2_X1 U472 ( .A(n534), .B(n533), .ZN(n641) );
  NOR2_X1 U473 ( .A1(n532), .A2(n531), .ZN(n534) );
  INV_X1 U474 ( .A(KEYINPUT41), .ZN(n376) );
  NOR2_X1 U475 ( .A1(n532), .A2(n620), .ZN(n627) );
  XNOR2_X1 U476 ( .A(G478), .B(n487), .ZN(n536) );
  NOR2_X1 U477 ( .A1(n547), .A2(n386), .ZN(n542) );
  XNOR2_X1 U478 ( .A(n436), .B(n514), .ZN(n435) );
  INV_X1 U479 ( .A(KEYINPUT16), .ZN(n437) );
  NAND2_X1 U480 ( .A1(n429), .A2(n737), .ZN(n727) );
  XNOR2_X1 U481 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U482 ( .A(n708), .B(n707), .ZN(n709) );
  INV_X1 U483 ( .A(n418), .ZN(n417) );
  AND2_X1 U484 ( .A1(n594), .A2(n356), .ZN(n595) );
  AND2_X1 U485 ( .A1(n405), .A2(n355), .ZN(n540) );
  XNOR2_X1 U486 ( .A(n391), .B(KEYINPUT32), .ZN(n746) );
  NOR2_X1 U487 ( .A1(n547), .A2(n548), .ZN(n391) );
  AND2_X1 U488 ( .A1(n411), .A2(n410), .ZN(n672) );
  XNOR2_X1 U489 ( .A(n387), .B(KEYINPUT119), .ZN(G54) );
  NAND2_X1 U490 ( .A1(n388), .A2(n410), .ZN(n387) );
  XNOR2_X1 U491 ( .A(n704), .B(n361), .ZN(n388) );
  INV_X1 U492 ( .A(KEYINPUT53), .ZN(n430) );
  AND2_X1 U493 ( .A1(n574), .A2(KEYINPUT39), .ZN(n354) );
  XOR2_X1 U494 ( .A(n580), .B(KEYINPUT71), .Z(n355) );
  NOR2_X1 U495 ( .A1(n593), .A2(n592), .ZN(n356) );
  AND2_X1 U496 ( .A1(n654), .A2(n653), .ZN(n357) );
  NOR2_X1 U497 ( .A1(n564), .A2(n427), .ZN(n358) );
  NOR2_X1 U498 ( .A1(n572), .A2(n573), .ZN(n359) );
  AND2_X1 U499 ( .A1(n421), .A2(n420), .ZN(n360) );
  INV_X1 U500 ( .A(KEYINPUT39), .ZN(n422) );
  XOR2_X1 U501 ( .A(n703), .B(n702), .Z(n361) );
  XOR2_X1 U502 ( .A(n657), .B(n656), .Z(n362) );
  XOR2_X1 U503 ( .A(n604), .B(KEYINPUT83), .Z(n363) );
  XNOR2_X1 U504 ( .A(n403), .B(n362), .ZN(n665) );
  XNOR2_X1 U505 ( .A(n568), .B(KEYINPUT105), .ZN(n635) );
  NOR2_X1 U506 ( .A1(n722), .A2(n665), .ZN(n667) );
  INV_X1 U507 ( .A(n722), .ZN(n410) );
  NOR2_X1 U508 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U509 ( .A1(n709), .A2(n722), .ZN(n371) );
  XNOR2_X1 U510 ( .A(n491), .B(n437), .ZN(n436) );
  BUF_X1 U511 ( .A(n650), .Z(n364) );
  XNOR2_X1 U512 ( .A(n409), .B(n363), .ZN(n367) );
  NAND2_X1 U513 ( .A1(n367), .A2(n408), .ZN(n368) );
  INV_X1 U514 ( .A(n535), .ZN(n389) );
  NAND2_X1 U515 ( .A1(n511), .A2(n512), .ZN(n366) );
  NOR2_X1 U516 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X2 U517 ( .A(n368), .B(KEYINPUT81), .ZN(n613) );
  XNOR2_X1 U518 ( .A(n440), .B(G137), .ZN(n380) );
  NAND2_X1 U519 ( .A1(n420), .A2(n378), .ZN(n416) );
  NOR2_X1 U520 ( .A1(n417), .A2(n416), .ZN(n576) );
  XNOR2_X1 U521 ( .A(n371), .B(n711), .ZN(G60) );
  XNOR2_X1 U522 ( .A(n520), .B(n519), .ZN(n524) );
  XNOR2_X1 U523 ( .A(n385), .B(n384), .ZN(n528) );
  NAND2_X1 U524 ( .A1(n389), .A2(n627), .ZN(n523) );
  XNOR2_X1 U525 ( .A(n525), .B(KEYINPUT91), .ZN(n374) );
  NOR2_X1 U526 ( .A1(n535), .A2(n522), .ZN(n511) );
  NAND2_X1 U527 ( .A1(n655), .A2(n660), .ZN(n502) );
  OR2_X2 U528 ( .A1(n635), .A2(n634), .ZN(n377) );
  XNOR2_X2 U529 ( .A(n502), .B(n501), .ZN(n578) );
  NOR2_X1 U530 ( .A1(n736), .A2(n607), .ZN(n608) );
  AND2_X2 U531 ( .A1(n613), .A2(n700), .ZN(n736) );
  NOR2_X1 U532 ( .A1(n650), .A2(n583), .ZN(n569) );
  INV_X1 U533 ( .A(n424), .ZN(n573) );
  NAND2_X1 U534 ( .A1(n424), .A2(n574), .ZN(n423) );
  NAND2_X1 U535 ( .A1(n603), .A2(n602), .ZN(n409) );
  INV_X1 U536 ( .A(n683), .ZN(n390) );
  XNOR2_X2 U537 ( .A(n397), .B(n550), .ZN(n658) );
  NAND2_X1 U538 ( .A1(n401), .A2(n398), .ZN(n397) );
  XNOR2_X1 U539 ( .A(n530), .B(n402), .ZN(n401) );
  NAND2_X1 U540 ( .A1(n716), .A2(G210), .ZN(n403) );
  INV_X1 U541 ( .A(n641), .ZN(n651) );
  XNOR2_X1 U542 ( .A(n407), .B(n406), .ZN(n405) );
  INV_X1 U543 ( .A(KEYINPUT34), .ZN(n406) );
  NAND2_X1 U544 ( .A1(n641), .A2(n389), .ZN(n407) );
  INV_X1 U545 ( .A(n358), .ZN(n408) );
  NAND2_X1 U546 ( .A1(n716), .A2(G472), .ZN(n412) );
  NAND2_X1 U547 ( .A1(n360), .A2(n418), .ZN(n605) );
  INV_X1 U548 ( .A(n575), .ZN(n419) );
  NAND2_X1 U549 ( .A1(n423), .A2(n422), .ZN(n420) );
  INV_X1 U550 ( .A(n578), .ZN(n427) );
  INV_X1 U551 ( .A(n607), .ZN(n428) );
  INV_X1 U552 ( .A(n658), .ZN(n429) );
  XNOR2_X1 U553 ( .A(n431), .B(n430), .ZN(G75) );
  NAND2_X1 U554 ( .A1(n432), .A2(n357), .ZN(n431) );
  XNOR2_X1 U555 ( .A(n434), .B(n433), .ZN(n432) );
  INV_X1 U556 ( .A(KEYINPUT79), .ZN(n433) );
  NAND2_X1 U557 ( .A1(n615), .A2(n664), .ZN(n434) );
  INV_X1 U558 ( .A(n364), .ZN(n629) );
  XNOR2_X1 U559 ( .A(n441), .B(KEYINPUT68), .ZN(n442) );
  INV_X1 U560 ( .A(KEYINPUT45), .ZN(n550) );
  XNOR2_X1 U561 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n734), .B(n518), .ZN(n701) );
  XNOR2_X1 U564 ( .A(n620), .B(n451), .ZN(n531) );
  XNOR2_X1 U565 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U566 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U567 ( .A1(G952), .A2(n737), .ZN(n722) );
  XOR2_X1 U568 ( .A(n493), .B(G131), .Z(n440) );
  XOR2_X1 U569 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n441) );
  INV_X1 U570 ( .A(n443), .ZN(n445) );
  XNOR2_X1 U571 ( .A(G113), .B(G101), .ZN(n444) );
  XNOR2_X1 U572 ( .A(n445), .B(n444), .ZN(n447) );
  NOR2_X1 U573 ( .A1(G953), .A2(G237), .ZN(n471) );
  NAND2_X1 U574 ( .A1(n471), .A2(G210), .ZN(n448) );
  NOR2_X1 U575 ( .A1(G902), .A2(n668), .ZN(n449) );
  XNOR2_X1 U576 ( .A(G472), .B(n449), .ZN(n450) );
  INV_X1 U577 ( .A(n531), .ZN(n558) );
  XNOR2_X1 U578 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U579 ( .A(n474), .B(n454), .ZN(n461) );
  NAND2_X1 U580 ( .A1(G234), .A2(n737), .ZN(n455) );
  XNOR2_X1 U581 ( .A(n456), .B(n455), .ZN(n481) );
  NAND2_X1 U582 ( .A1(G221), .A2(n481), .ZN(n459) );
  XNOR2_X1 U583 ( .A(n457), .B(KEYINPUT24), .ZN(n458) );
  NAND2_X1 U584 ( .A1(n660), .A2(G234), .ZN(n463) );
  XNOR2_X1 U585 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n462) );
  XNOR2_X1 U586 ( .A(n463), .B(n462), .ZN(n488) );
  NAND2_X1 U587 ( .A1(G217), .A2(n488), .ZN(n464) );
  XOR2_X1 U588 ( .A(KEYINPUT100), .B(n552), .Z(n617) );
  XNOR2_X1 U589 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n477) );
  XNOR2_X1 U590 ( .A(n466), .B(n465), .ZN(n470) );
  XNOR2_X1 U591 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U592 ( .A(n470), .B(n469), .Z(n473) );
  NAND2_X1 U593 ( .A1(n471), .A2(G214), .ZN(n472) );
  XNOR2_X1 U594 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n475), .B(n474), .ZN(n706) );
  NOR2_X1 U596 ( .A1(G902), .A2(n706), .ZN(n476) );
  XNOR2_X1 U597 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U598 ( .A(G475), .B(n478), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n480) );
  XNOR2_X1 U600 ( .A(G116), .B(KEYINPUT96), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n480), .B(n479), .ZN(n486) );
  NAND2_X1 U602 ( .A1(G217), .A2(n481), .ZN(n484) );
  XNOR2_X1 U603 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U604 ( .A(n486), .B(n485), .ZN(n712) );
  NOR2_X1 U605 ( .A1(G902), .A2(n712), .ZN(n487) );
  NAND2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n634) );
  INV_X1 U607 ( .A(n634), .ZN(n512) );
  NAND2_X1 U608 ( .A1(n488), .A2(G221), .ZN(n489) );
  XOR2_X1 U609 ( .A(n489), .B(KEYINPUT21), .Z(n616) );
  INV_X1 U610 ( .A(n616), .ZN(n522) );
  OR2_X1 U611 ( .A1(G237), .A2(G902), .ZN(n500) );
  NAND2_X1 U612 ( .A1(G214), .A2(n500), .ZN(n631) );
  XNOR2_X1 U613 ( .A(KEYINPUT69), .B(KEYINPUT86), .ZN(n490) );
  NAND2_X1 U614 ( .A1(G224), .A2(n737), .ZN(n496) );
  NAND2_X1 U615 ( .A1(G210), .A2(n500), .ZN(n501) );
  NOR2_X1 U616 ( .A1(G898), .A2(n737), .ZN(n729) );
  NAND2_X1 U617 ( .A1(G234), .A2(G237), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n503), .B(KEYINPUT87), .ZN(n504) );
  XOR2_X1 U619 ( .A(KEYINPUT14), .B(n504), .Z(n506) );
  NAND2_X1 U620 ( .A1(G902), .A2(n506), .ZN(n553) );
  INV_X1 U621 ( .A(n553), .ZN(n505) );
  NAND2_X1 U622 ( .A1(n729), .A2(n505), .ZN(n508) );
  NAND2_X1 U623 ( .A1(n506), .A2(G952), .ZN(n647) );
  NOR2_X1 U624 ( .A1(G953), .A2(n647), .ZN(n507) );
  XOR2_X1 U625 ( .A(KEYINPUT88), .B(n507), .Z(n556) );
  NAND2_X1 U626 ( .A1(n508), .A2(n556), .ZN(n509) );
  NAND2_X1 U627 ( .A1(n584), .A2(n509), .ZN(n510) );
  NAND2_X1 U628 ( .A1(G227), .A2(n737), .ZN(n516) );
  NOR2_X1 U629 ( .A1(G902), .A2(n701), .ZN(n520) );
  NAND2_X1 U630 ( .A1(n617), .A2(n542), .ZN(n521) );
  NOR2_X1 U631 ( .A1(n558), .A2(n521), .ZN(n673) );
  XNOR2_X1 U632 ( .A(n523), .B(KEYINPUT31), .ZN(n695) );
  NAND2_X1 U633 ( .A1(n524), .A2(n622), .ZN(n572) );
  INV_X1 U634 ( .A(n537), .ZN(n526) );
  NAND2_X1 U635 ( .A1(n536), .A2(n526), .ZN(n575) );
  NOR2_X1 U636 ( .A1(n526), .A2(n536), .ZN(n694) );
  XOR2_X1 U637 ( .A(KEYINPUT98), .B(n694), .Z(n606) );
  NAND2_X1 U638 ( .A1(n575), .A2(n606), .ZN(n586) );
  XNOR2_X1 U639 ( .A(n586), .B(KEYINPUT77), .ZN(n527) );
  INV_X1 U640 ( .A(KEYINPUT33), .ZN(n533) );
  OR2_X1 U641 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U642 ( .A(KEYINPUT103), .B(n538), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT35), .B(KEYINPUT70), .ZN(n539) );
  AND2_X1 U644 ( .A1(n620), .A2(n552), .ZN(n541) );
  NAND2_X1 U645 ( .A1(n542), .A2(n541), .ZN(n683) );
  NOR2_X1 U646 ( .A1(n543), .A2(n617), .ZN(n544) );
  XNOR2_X1 U647 ( .A(n544), .B(KEYINPUT102), .ZN(n546) );
  XOR2_X1 U648 ( .A(n558), .B(KEYINPUT72), .Z(n545) );
  NAND2_X1 U649 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U650 ( .A(n551), .B(KEYINPUT78), .ZN(n609) );
  NAND2_X1 U651 ( .A1(n616), .A2(n552), .ZN(n593) );
  INV_X1 U652 ( .A(n593), .ZN(n561) );
  NOR2_X1 U653 ( .A1(G900), .A2(n553), .ZN(n554) );
  NAND2_X1 U654 ( .A1(G953), .A2(n554), .ZN(n555) );
  XNOR2_X1 U655 ( .A(KEYINPUT104), .B(n555), .ZN(n557) );
  NAND2_X1 U656 ( .A1(n557), .A2(n556), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n631), .A2(n579), .ZN(n560) );
  NAND2_X1 U658 ( .A1(n419), .A2(n558), .ZN(n559) );
  NAND2_X1 U659 ( .A1(n561), .A2(n594), .ZN(n562) );
  NOR2_X1 U660 ( .A1(n386), .A2(n562), .ZN(n563) );
  XNOR2_X1 U661 ( .A(n563), .B(KEYINPUT43), .ZN(n564) );
  NAND2_X1 U662 ( .A1(n570), .A2(n579), .ZN(n565) );
  NOR2_X1 U663 ( .A1(n593), .A2(n565), .ZN(n566) );
  XNOR2_X1 U664 ( .A(KEYINPUT28), .B(n566), .ZN(n567) );
  NAND2_X1 U665 ( .A1(n567), .A2(n524), .ZN(n583) );
  XNOR2_X1 U666 ( .A(n569), .B(KEYINPUT42), .ZN(n748) );
  AND2_X1 U667 ( .A1(n632), .A2(n579), .ZN(n574) );
  XNOR2_X1 U668 ( .A(KEYINPUT40), .B(n576), .ZN(n747) );
  XNOR2_X1 U669 ( .A(n577), .B(KEYINPUT46), .ZN(n590) );
  BUF_X1 U670 ( .A(n578), .Z(n592) );
  AND2_X1 U671 ( .A1(n359), .A2(n579), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U673 ( .A1(n592), .A2(n582), .ZN(n688) );
  INV_X1 U674 ( .A(n583), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n585), .A2(n584), .ZN(n684) );
  INV_X1 U676 ( .A(n586), .ZN(n636) );
  NAND2_X1 U677 ( .A1(n636), .A2(KEYINPUT77), .ZN(n587) );
  NOR2_X1 U678 ( .A1(n684), .A2(n587), .ZN(n588) );
  NOR2_X1 U679 ( .A1(n688), .A2(n588), .ZN(n589) );
  NOR2_X1 U680 ( .A1(n684), .A2(n636), .ZN(n598) );
  INV_X1 U681 ( .A(n598), .ZN(n591) );
  NAND2_X1 U682 ( .A1(n591), .A2(KEYINPUT47), .ZN(n601) );
  XNOR2_X1 U683 ( .A(n595), .B(KEYINPUT36), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n596), .A2(n386), .ZN(n697) );
  NOR2_X1 U685 ( .A1(KEYINPUT77), .A2(KEYINPUT47), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U687 ( .A1(n697), .A2(n599), .ZN(n600) );
  AND2_X1 U688 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n700) );
  XNOR2_X1 U690 ( .A(n610), .B(KEYINPUT74), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n700), .A2(KEYINPUT2), .ZN(n611) );
  XOR2_X1 U692 ( .A(KEYINPUT73), .B(n611), .Z(n612) );
  NOR2_X1 U693 ( .A1(n658), .A2(n612), .ZN(n614) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n618), .B(KEYINPUT49), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n625) );
  NOR2_X1 U697 ( .A1(n622), .A2(n386), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT50), .ZN(n624) );
  NOR2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n628), .B(KEYINPUT51), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n644) );
  NOR2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT114), .ZN(n638) );
  NOR2_X1 U707 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U708 ( .A(KEYINPUT115), .B(n640), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n644), .A2(n643), .ZN(n646) );
  XOR2_X1 U711 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n645) );
  XNOR2_X1 U712 ( .A(n646), .B(n645), .ZN(n648) );
  NOR2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U714 ( .A1(G953), .A2(n649), .ZN(n654) );
  NOR2_X1 U715 ( .A1(n651), .A2(n364), .ZN(n652) );
  XNOR2_X1 U716 ( .A(n652), .B(KEYINPUT117), .ZN(n653) );
  XNOR2_X1 U717 ( .A(KEYINPUT55), .B(KEYINPUT75), .ZN(n657) );
  XNOR2_X1 U718 ( .A(n655), .B(KEYINPUT54), .ZN(n656) );
  NAND2_X1 U719 ( .A1(n659), .A2(n736), .ZN(n663) );
  XOR2_X1 U720 ( .A(KEYINPUT80), .B(n660), .Z(n661) );
  NAND2_X1 U721 ( .A1(KEYINPUT2), .A2(n661), .ZN(n662) );
  XNOR2_X1 U722 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n666) );
  XNOR2_X1 U723 ( .A(n667), .B(n666), .ZN(G51) );
  XOR2_X1 U724 ( .A(KEYINPUT62), .B(n668), .Z(n669) );
  XNOR2_X1 U725 ( .A(KEYINPUT63), .B(KEYINPUT84), .ZN(n670) );
  XNOR2_X1 U726 ( .A(n670), .B(KEYINPUT85), .ZN(n671) );
  XNOR2_X1 U727 ( .A(n672), .B(n671), .ZN(G57) );
  XOR2_X1 U728 ( .A(G101), .B(n673), .Z(n674) );
  XNOR2_X1 U729 ( .A(KEYINPUT106), .B(n674), .ZN(G3) );
  XOR2_X1 U730 ( .A(G104), .B(KEYINPUT107), .Z(n676) );
  NAND2_X1 U731 ( .A1(n350), .A2(n419), .ZN(n675) );
  XNOR2_X1 U732 ( .A(n676), .B(n675), .ZN(G6) );
  XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT26), .ZN(n681) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT108), .Z(n679) );
  NAND2_X1 U735 ( .A1(n350), .A2(n694), .ZN(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n681), .B(n680), .ZN(G9) );
  XOR2_X1 U738 ( .A(G110), .B(KEYINPUT109), .Z(n682) );
  XNOR2_X1 U739 ( .A(n683), .B(n682), .ZN(G12) );
  XOR2_X1 U740 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n686) );
  INV_X1 U741 ( .A(n684), .ZN(n689) );
  NAND2_X1 U742 ( .A1(n694), .A2(n689), .ZN(n685) );
  XNOR2_X1 U743 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U744 ( .A(G128), .B(n687), .ZN(G30) );
  XOR2_X1 U745 ( .A(G143), .B(n688), .Z(G45) );
  XOR2_X1 U746 ( .A(G146), .B(KEYINPUT111), .Z(n691) );
  NAND2_X1 U747 ( .A1(n689), .A2(n419), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n691), .B(n690), .ZN(G48) );
  NAND2_X1 U749 ( .A1(n695), .A2(n419), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n692), .B(KEYINPUT112), .ZN(n693) );
  XNOR2_X1 U751 ( .A(G113), .B(n693), .ZN(G15) );
  NAND2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n696), .B(G116), .ZN(G18) );
  XNOR2_X1 U754 ( .A(KEYINPUT37), .B(KEYINPUT113), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U756 ( .A(G125), .B(n699), .ZN(G27) );
  XNOR2_X1 U757 ( .A(G134), .B(n700), .ZN(G36) );
  XOR2_X1 U758 ( .A(G140), .B(n358), .Z(G42) );
  XOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U760 ( .A(n701), .B(KEYINPUT118), .ZN(n702) );
  NAND2_X1 U761 ( .A1(n716), .A2(G469), .ZN(n704) );
  NAND2_X1 U762 ( .A1(n716), .A2(G475), .ZN(n708) );
  XOR2_X1 U763 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n705) );
  XNOR2_X1 U764 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n710), .B(KEYINPUT65), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT122), .ZN(n714) );
  NAND2_X1 U767 ( .A1(G478), .A2(n716), .ZN(n713) );
  XNOR2_X1 U768 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n722), .A2(n715), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n716), .A2(G217), .ZN(n720) );
  INV_X1 U771 ( .A(KEYINPUT123), .ZN(n717) );
  XNOR2_X1 U772 ( .A(KEYINPUT124), .B(n723), .ZN(G66) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n724) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n724), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n728), .B(KEYINPUT125), .ZN(n732) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U779 ( .A(n732), .B(n731), .Z(G69) );
  XNOR2_X1 U780 ( .A(n734), .B(n733), .ZN(n739) );
  INV_X1 U781 ( .A(n739), .ZN(n735) );
  XOR2_X1 U782 ( .A(n736), .B(n735), .Z(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(n737), .ZN(n743) );
  XOR2_X1 U784 ( .A(G227), .B(n739), .Z(n740) );
  NAND2_X1 U785 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U786 ( .A1(n741), .A2(G953), .ZN(n742) );
  NAND2_X1 U787 ( .A1(n743), .A2(n742), .ZN(G72) );
  XNOR2_X1 U788 ( .A(G122), .B(n744), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n745), .B(KEYINPUT126), .ZN(G24) );
  XOR2_X1 U790 ( .A(G119), .B(n746), .Z(G21) );
  XOR2_X1 U791 ( .A(n747), .B(G131), .Z(G33) );
  XOR2_X1 U792 ( .A(n748), .B(G137), .Z(G39) );
endmodule

