

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(G651), .A2(n627), .ZN(n637) );
  XNOR2_X1 U547 ( .A(n574), .B(KEYINPUT81), .ZN(n511) );
  NOR2_X1 U548 ( .A1(n698), .A2(n987), .ZN(n700) );
  INV_X1 U549 ( .A(KEYINPUT29), .ZN(n718) );
  NOR2_X1 U550 ( .A1(G1384), .A2(G164), .ZN(n676) );
  AND2_X1 U551 ( .A1(n575), .A2(n511), .ZN(n576) );
  NOR2_X2 U552 ( .A1(G2104), .A2(n517), .ZN(n883) );
  XOR2_X1 U553 ( .A(KEYINPUT1), .B(n537), .Z(n638) );
  NOR2_X1 U554 ( .A1(n523), .A2(n522), .ZN(G160) );
  INV_X1 U555 ( .A(G2105), .ZN(n517) );
  INV_X1 U556 ( .A(G2104), .ZN(n515) );
  NOR2_X1 U557 ( .A1(n517), .A2(n515), .ZN(n884) );
  NAND2_X1 U558 ( .A1(n884), .A2(G113), .ZN(n514) );
  NOR2_X2 U559 ( .A1(G2105), .A2(G2104), .ZN(n512) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n512), .Z(n888) );
  NAND2_X1 U561 ( .A1(n888), .A2(G137), .ZN(n513) );
  NAND2_X1 U562 ( .A1(n514), .A2(n513), .ZN(n523) );
  NOR2_X2 U563 ( .A1(G2105), .A2(n515), .ZN(n887) );
  NAND2_X1 U564 ( .A1(n887), .A2(G101), .ZN(n516) );
  XNOR2_X1 U565 ( .A(KEYINPUT23), .B(n516), .ZN(n520) );
  NAND2_X1 U566 ( .A1(n883), .A2(G125), .ZN(n518) );
  XOR2_X1 U567 ( .A(KEYINPUT66), .B(n518), .Z(n519) );
  NOR2_X1 U568 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U569 ( .A(n521), .B(KEYINPUT67), .ZN(n522) );
  NAND2_X1 U570 ( .A1(G138), .A2(n888), .ZN(n525) );
  NAND2_X1 U571 ( .A1(G126), .A2(n883), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U573 ( .A1(G102), .A2(n887), .ZN(n527) );
  NAND2_X1 U574 ( .A1(G114), .A2(n884), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U576 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U577 ( .A(n530), .B(KEYINPUT93), .Z(G164) );
  XOR2_X1 U578 ( .A(KEYINPUT68), .B(G651), .Z(n536) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  NOR2_X1 U580 ( .A1(n536), .A2(n627), .ZN(n641) );
  NAND2_X1 U581 ( .A1(n641), .A2(G77), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n531), .B(KEYINPUT70), .ZN(n534) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT65), .B(n532), .Z(n642) );
  NAND2_X1 U585 ( .A1(G90), .A2(n642), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U587 ( .A(KEYINPUT9), .B(n535), .ZN(n541) );
  NAND2_X1 U588 ( .A1(G52), .A2(n637), .ZN(n539) );
  NOR2_X1 U589 ( .A1(n536), .A2(G543), .ZN(n537) );
  NAND2_X1 U590 ( .A1(G64), .A2(n638), .ZN(n538) );
  AND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(G301) );
  INV_X1 U593 ( .A(G301), .ZN(G171) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U595 ( .A(G132), .ZN(G219) );
  INV_X1 U596 ( .A(G82), .ZN(G220) );
  INV_X1 U597 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U598 ( .A(KEYINPUT84), .B(KEYINPUT6), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G51), .A2(n637), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G63), .A2(n638), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n545), .B(n544), .ZN(n552) );
  NAND2_X1 U603 ( .A1(n642), .A2(G89), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G76), .A2(n641), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U607 ( .A(KEYINPUT83), .B(n549), .ZN(n550) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n550), .ZN(n551) );
  NOR2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(n553), .Z(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n554), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U614 ( .A(G223), .ZN(n825) );
  NAND2_X1 U615 ( .A1(n825), .A2(G567), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT75), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT11), .B(n556), .ZN(G234) );
  XOR2_X1 U618 ( .A(G860), .B(KEYINPUT78), .Z(n591) );
  NAND2_X1 U619 ( .A1(n641), .A2(G68), .ZN(n557) );
  XNOR2_X1 U620 ( .A(KEYINPUT76), .B(n557), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n642), .A2(G81), .ZN(n558) );
  XNOR2_X1 U622 ( .A(KEYINPUT12), .B(n558), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U624 ( .A(n561), .B(KEYINPUT13), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G43), .A2(n637), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n638), .A2(G56), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT77), .B(n567), .ZN(n987) );
  OR2_X1 U631 ( .A1(n591), .A2(n987), .ZN(G153) );
  NAND2_X1 U632 ( .A1(G92), .A2(n642), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G66), .A2(n638), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT79), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n637), .A2(G54), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT80), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G79), .A2(n641), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT15), .B(n576), .Z(n577) );
  XNOR2_X2 U641 ( .A(KEYINPUT82), .B(n577), .ZN(n1002) );
  INV_X1 U642 ( .A(n1002), .ZN(n595) );
  NOR2_X1 U643 ( .A1(n595), .A2(G868), .ZN(n579) );
  INV_X1 U644 ( .A(G868), .ZN(n658) );
  NOR2_X1 U645 ( .A1(n658), .A2(G301), .ZN(n578) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(G284) );
  NAND2_X1 U647 ( .A1(n638), .A2(G65), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT72), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G53), .A2(n637), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U651 ( .A(n583), .B(KEYINPUT73), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G78), .A2(n641), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G91), .A2(n642), .ZN(n586) );
  XNOR2_X1 U655 ( .A(KEYINPUT71), .B(n586), .ZN(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n988) );
  XOR2_X1 U657 ( .A(n988), .B(KEYINPUT74), .Z(G299) );
  NOR2_X1 U658 ( .A1(G299), .A2(G868), .ZN(n590) );
  NOR2_X1 U659 ( .A1(G286), .A2(n658), .ZN(n589) );
  NOR2_X1 U660 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U661 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n592), .A2(n1002), .ZN(n593) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT85), .ZN(n594) );
  XOR2_X1 U664 ( .A(KEYINPUT16), .B(n594), .Z(G148) );
  OR2_X1 U665 ( .A1(G559), .A2(n595), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n596), .A2(G868), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n987), .A2(n658), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U669 ( .A1(n883), .A2(G123), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G111), .A2(n884), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G99), .A2(n887), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G135), .A2(n888), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n959) );
  XNOR2_X1 U677 ( .A(G2096), .B(n959), .ZN(n607) );
  INV_X1 U678 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U680 ( .A1(n1002), .A2(G559), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(n987), .ZN(n654) );
  NOR2_X1 U682 ( .A1(n654), .A2(G860), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G80), .A2(n641), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G93), .A2(n642), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G55), .A2(n637), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G67), .A2(n638), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n613) );
  OR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n657) );
  XOR2_X1 U690 ( .A(n615), .B(n657), .Z(G145) );
  NAND2_X1 U691 ( .A1(G61), .A2(n638), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT86), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G86), .A2(n642), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G48), .A2(n637), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n641), .A2(G73), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT2), .B(n619), .Z(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(G305) );
  NAND2_X1 U700 ( .A1(G49), .A2(n637), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n638), .A2(n626), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G85), .A2(n642), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G47), .A2(n637), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G72), .A2(n641), .ZN(n632) );
  XNOR2_X1 U710 ( .A(KEYINPUT69), .B(n632), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n638), .A2(G60), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G50), .A2(n637), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G62), .A2(n638), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n647) );
  NAND2_X1 U717 ( .A1(G75), .A2(n641), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G88), .A2(n642), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U720 ( .A(KEYINPUT87), .B(n645), .Z(n646) );
  NOR2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U722 ( .A(KEYINPUT88), .B(n648), .Z(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U724 ( .A(KEYINPUT19), .B(G305), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(G288), .ZN(n650) );
  XOR2_X1 U726 ( .A(n657), .B(n650), .Z(n652) );
  XNOR2_X1 U727 ( .A(G290), .B(G299), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(G166), .ZN(n850) );
  XNOR2_X1 U730 ( .A(KEYINPUT89), .B(n654), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n850), .B(n655), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U739 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(KEYINPUT90), .B(G44), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U742 ( .A1(G120), .A2(G108), .ZN(n666) );
  NOR2_X1 U743 ( .A1(G235), .A2(n666), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n667), .A2(G57), .ZN(n668) );
  XOR2_X1 U745 ( .A(KEYINPUT91), .B(n668), .Z(n829) );
  NAND2_X1 U746 ( .A1(n829), .A2(G567), .ZN(n673) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U749 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(G96), .A2(n671), .ZN(n830) );
  NAND2_X1 U751 ( .A1(n830), .A2(G2106), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n855) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n674) );
  XNOR2_X1 U754 ( .A(KEYINPUT92), .B(n674), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n855), .A2(n675), .ZN(n828) );
  NAND2_X1 U756 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U758 ( .A(n768), .ZN(n677) );
  XNOR2_X1 U759 ( .A(n676), .B(KEYINPUT64), .ZN(n767) );
  NAND2_X1 U760 ( .A1(n677), .A2(n767), .ZN(n694) );
  NAND2_X1 U761 ( .A1(G8), .A2(n694), .ZN(n759) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n678) );
  XNOR2_X1 U763 ( .A(n678), .B(KEYINPUT95), .ZN(n679) );
  XNOR2_X1 U764 ( .A(KEYINPUT24), .B(n679), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n759), .A2(n680), .ZN(n749) );
  NOR2_X1 U766 ( .A1(G303), .A2(G2090), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G8), .A2(n681), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n682), .B(KEYINPUT102), .ZN(n746) );
  NOR2_X1 U769 ( .A1(G1966), .A2(n759), .ZN(n724) );
  BUF_X2 U770 ( .A(n694), .Z(n730) );
  NOR2_X1 U771 ( .A1(G2084), .A2(n730), .ZN(n726) );
  NOR2_X1 U772 ( .A1(n724), .A2(n726), .ZN(n683) );
  NAND2_X1 U773 ( .A1(G8), .A2(n683), .ZN(n684) );
  XNOR2_X1 U774 ( .A(KEYINPUT99), .B(n684), .ZN(n685) );
  XOR2_X1 U775 ( .A(KEYINPUT30), .B(n685), .Z(n686) );
  NOR2_X1 U776 ( .A1(G168), .A2(n686), .ZN(n691) );
  INV_X1 U777 ( .A(n730), .ZN(n708) );
  NOR2_X1 U778 ( .A1(n708), .A2(G1961), .ZN(n687) );
  XOR2_X1 U779 ( .A(KEYINPUT96), .B(n687), .Z(n689) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .ZN(n947) );
  NAND2_X1 U781 ( .A1(n708), .A2(n947), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n720) );
  NOR2_X1 U783 ( .A1(G171), .A2(n720), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U785 ( .A(KEYINPUT31), .B(n692), .Z(n734) );
  INV_X1 U786 ( .A(G1996), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U788 ( .A(KEYINPUT26), .B(n695), .Z(n697) );
  NAND2_X1 U789 ( .A1(n730), .A2(G1341), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n700), .A2(n1002), .ZN(n699) );
  XNOR2_X1 U792 ( .A(n699), .B(KEYINPUT97), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n700), .A2(n1002), .ZN(n704) );
  NOR2_X1 U794 ( .A1(n708), .A2(G1348), .ZN(n702) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n730), .ZN(n701) );
  NOR2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n712) );
  NAND2_X1 U799 ( .A1(n708), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U801 ( .A(G1956), .ZN(n923) );
  NOR2_X1 U802 ( .A1(n923), .A2(n708), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n988), .A2(n713), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n988), .A2(n713), .ZN(n714) );
  XNOR2_X1 U807 ( .A(n714), .B(KEYINPUT28), .ZN(n715) );
  INV_X1 U808 ( .A(n715), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U810 ( .A(n719), .B(n718), .ZN(n722) );
  NAND2_X1 U811 ( .A1(G171), .A2(n720), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U813 ( .A(n723), .B(KEYINPUT98), .ZN(n736) );
  AND2_X1 U814 ( .A1(n734), .A2(n736), .ZN(n725) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U816 ( .A1(G8), .A2(n726), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U818 ( .A(KEYINPUT100), .B(n729), .ZN(n745) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n759), .ZN(n732) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U822 ( .A1(G303), .A2(n733), .ZN(n737) );
  AND2_X1 U823 ( .A1(n734), .A2(n737), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n740) );
  INV_X1 U825 ( .A(n737), .ZN(n738) );
  OR2_X1 U826 ( .A1(n738), .A2(G286), .ZN(n739) );
  AND2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U828 ( .A1(G8), .A2(n741), .ZN(n743) );
  XOR2_X1 U829 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n742) );
  XNOR2_X1 U830 ( .A(n743), .B(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n753) );
  NAND2_X1 U832 ( .A1(n746), .A2(n753), .ZN(n747) );
  AND2_X1 U833 ( .A1(n747), .A2(n759), .ZN(n748) );
  NOR2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n766) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n758) );
  NOR2_X1 U836 ( .A1(G303), .A2(G1971), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n758), .A2(n750), .ZN(n1001) );
  INV_X1 U838 ( .A(KEYINPUT33), .ZN(n751) );
  AND2_X1 U839 ( .A1(n1001), .A2(n751), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n757) );
  INV_X1 U841 ( .A(n759), .ZN(n754) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n994) );
  AND2_X1 U843 ( .A1(n754), .A2(n994), .ZN(n755) );
  OR2_X1 U844 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  AND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n764) );
  NAND2_X1 U846 ( .A1(n758), .A2(KEYINPUT33), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n762) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n991) );
  INV_X1 U849 ( .A(n991), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  AND2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n796) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n809) );
  NAND2_X1 U854 ( .A1(G104), .A2(n887), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G140), .A2(n888), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U857 ( .A(KEYINPUT34), .B(n771), .ZN(n776) );
  NAND2_X1 U858 ( .A1(G128), .A2(n883), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G116), .A2(n884), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U861 ( .A(KEYINPUT35), .B(n774), .Z(n775) );
  NOR2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U863 ( .A(KEYINPUT36), .B(n777), .ZN(n897) );
  XNOR2_X1 U864 ( .A(KEYINPUT37), .B(G2067), .ZN(n807) );
  NOR2_X1 U865 ( .A1(n897), .A2(n807), .ZN(n974) );
  NAND2_X1 U866 ( .A1(n809), .A2(n974), .ZN(n805) );
  NAND2_X1 U867 ( .A1(G119), .A2(n883), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G131), .A2(n888), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n887), .A2(G95), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT94), .B(n780), .Z(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n884), .A2(G107), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n872) );
  AND2_X1 U875 ( .A1(n872), .A2(G1991), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G129), .A2(n883), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G141), .A2(n888), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n887), .A2(G105), .ZN(n787) );
  XOR2_X1 U880 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n884), .A2(G117), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n873) );
  AND2_X1 U884 ( .A1(n873), .A2(G1996), .ZN(n792) );
  NOR2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n965) );
  INV_X1 U886 ( .A(n809), .ZN(n797) );
  NOR2_X1 U887 ( .A1(n965), .A2(n797), .ZN(n802) );
  INV_X1 U888 ( .A(n802), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n805), .A2(n794), .ZN(n795) );
  NOR2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n799) );
  XOR2_X1 U891 ( .A(G1986), .B(G290), .Z(n995) );
  OR2_X1 U892 ( .A1(n995), .A2(n797), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n812) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n873), .ZN(n971) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n872), .ZN(n960) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n960), .A2(n800), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n971), .A2(n803), .ZN(n804) );
  XNOR2_X1 U900 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n897), .A2(n807), .ZN(n964) );
  NAND2_X1 U903 ( .A1(n808), .A2(n964), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U906 ( .A(n813), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U907 ( .A(G2427), .B(G2451), .ZN(n823) );
  XOR2_X1 U908 ( .A(G2430), .B(G2443), .Z(n815) );
  XNOR2_X1 U909 ( .A(G2435), .B(KEYINPUT103), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(n819) );
  XOR2_X1 U911 ( .A(G2438), .B(G2454), .Z(n817) );
  XNOR2_X1 U912 ( .A(G1348), .B(G1341), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n817), .B(n816), .ZN(n818) );
  XOR2_X1 U914 ( .A(n819), .B(n818), .Z(n821) );
  XNOR2_X1 U915 ( .A(KEYINPUT104), .B(G2446), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(G14), .ZN(n903) );
  XNOR2_X1 U919 ( .A(KEYINPUT105), .B(n903), .ZN(G401) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U922 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U925 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  XNOR2_X1 U926 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U931 ( .A(G1956), .B(G2474), .ZN(n840) );
  XOR2_X1 U932 ( .A(G1976), .B(G1981), .Z(n832) );
  XNOR2_X1 U933 ( .A(G1966), .B(G1961), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U935 ( .A(G1971), .B(G1986), .Z(n834) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U937 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U938 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U939 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U942 ( .A(KEYINPUT107), .B(G2084), .Z(n842) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n843), .B(G2096), .Z(n845) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n847) );
  XNOR2_X1 U949 ( .A(G2678), .B(G2100), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(G227) );
  XNOR2_X1 U952 ( .A(n987), .B(n850), .ZN(n852) );
  XNOR2_X1 U953 ( .A(G286), .B(G171), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(n1002), .ZN(n854) );
  NOR2_X1 U956 ( .A1(G37), .A2(n854), .ZN(G397) );
  INV_X1 U957 ( .A(n855), .ZN(G319) );
  NAND2_X1 U958 ( .A1(G112), .A2(n884), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n856), .B(KEYINPUT110), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n858) );
  NAND2_X1 U961 ( .A1(G124), .A2(n883), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G100), .A2(n887), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G136), .A2(n888), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G103), .A2(n887), .ZN(n866) );
  NAND2_X1 U969 ( .A1(G139), .A2(n888), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G127), .A2(n883), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G115), .A2(n884), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n966) );
  XOR2_X1 U976 ( .A(G162), .B(n966), .Z(n875) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n882) );
  XOR2_X1 U979 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n877) );
  XNOR2_X1 U980 ( .A(KEYINPUT114), .B(KEYINPUT113), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(n878), .B(n959), .Z(n880) );
  XNOR2_X1 U983 ( .A(G164), .B(G160), .ZN(n879) );
  XNOR2_X1 U984 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U985 ( .A(n882), .B(n881), .ZN(n899) );
  NAND2_X1 U986 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n895) );
  XNOR2_X1 U989 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n887), .A2(G106), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n888), .A2(G142), .ZN(n889) );
  XOR2_X1 U992 ( .A(KEYINPUT111), .B(n889), .Z(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U999 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n903), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G397), .A2(n904), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n907), .A2(G395), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1007 ( .A(G308), .ZN(G225) );
  INV_X1 U1008 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1009 ( .A(G1986), .B(G24), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G1971), .B(G22), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(G23), .B(G1976), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n913) );
  XNOR2_X1 U1015 ( .A(n914), .B(n913), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G1966), .B(G21), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(G5), .B(G1961), .ZN(n915) );
  NOR2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n931) );
  XOR2_X1 U1020 ( .A(G1341), .B(G19), .Z(n919) );
  XNOR2_X1 U1021 ( .A(KEYINPUT125), .B(n919), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G6), .B(G1981), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(KEYINPUT126), .B(n922), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n923), .B(G20), .ZN(n924) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1027 ( .A(KEYINPUT59), .B(G1348), .Z(n926) );
  XNOR2_X1 U1028 ( .A(G4), .B(n926), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1030 ( .A(KEYINPUT60), .B(n929), .Z(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(KEYINPUT61), .B(n932), .ZN(n934) );
  INV_X1 U1033 ( .A(G16), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n935), .A2(G11), .ZN(n986) );
  XOR2_X1 U1036 ( .A(KEYINPUT122), .B(G34), .Z(n937) );
  XNOR2_X1 U1037 ( .A(G2084), .B(KEYINPUT54), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(n937), .B(n936), .ZN(n954) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(G2072), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n938), .B(G33), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(G1991), .B(G25), .ZN(n939) );
  NOR2_X1 U1044 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1045 ( .A1(G28), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(KEYINPUT120), .B(G2067), .ZN(n942) );
  XNOR2_X1 U1047 ( .A(G26), .B(n942), .ZN(n943) );
  NOR2_X1 U1048 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1050 ( .A(G27), .B(n947), .Z(n948) );
  NOR2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n950), .ZN(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(KEYINPUT123), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(G29), .A2(n956), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(n957), .B(KEYINPUT55), .ZN(n984) );
  XNOR2_X1 U1058 ( .A(G160), .B(G2084), .ZN(n958) );
  XNOR2_X1 U1059 ( .A(n958), .B(KEYINPUT118), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1062 ( .A(KEYINPUT119), .B(n963), .ZN(n980) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n978) );
  XOR2_X1 U1064 ( .A(G2072), .B(n966), .Z(n968) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n969), .ZN(n976) );
  XOR2_X1 U1068 ( .A(G2090), .B(G162), .Z(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(n972), .B(KEYINPUT51), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT52), .B(n981), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(G29), .A2(n982), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n1013) );
  XOR2_X1 U1079 ( .A(n987), .B(G1341), .Z(n990) );
  XNOR2_X1 U1080 ( .A(n988), .B(G1956), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1008) );
  XNOR2_X1 U1082 ( .A(G168), .B(G1966), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT57), .ZN(n1006) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1961), .B(G171), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(G1348), .B(n1002), .Z(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(KEYINPUT124), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1096 ( .A(G16), .B(KEYINPUT56), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1014), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

