

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725;

  NOR2_X1 U364 ( .A1(n392), .A2(n387), .ZN(n611) );
  NOR2_X1 U365 ( .A1(n579), .A2(n367), .ZN(n584) );
  NOR2_X1 U366 ( .A1(n574), .A2(n667), .ZN(n575) );
  XNOR2_X1 U367 ( .A(n383), .B(KEYINPUT19), .ZN(n565) );
  XNOR2_X1 U368 ( .A(n433), .B(n432), .ZN(n475) );
  XNOR2_X2 U369 ( .A(n362), .B(n409), .ZN(n675) );
  INV_X1 U370 ( .A(G953), .ZN(n714) );
  XNOR2_X2 U371 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n432) );
  XNOR2_X2 U372 ( .A(n459), .B(KEYINPUT4), .ZN(n710) );
  NOR2_X2 U373 ( .A1(G902), .A2(n604), .ZN(n482) );
  XNOR2_X1 U374 ( .A(n601), .B(n600), .ZN(n713) );
  NOR2_X2 U375 ( .A1(n725), .A2(n724), .ZN(n544) );
  XNOR2_X1 U376 ( .A(n425), .B(n408), .ZN(n481) );
  INV_X2 U377 ( .A(G143), .ZN(n416) );
  OR2_X1 U378 ( .A1(n599), .A2(n697), .ZN(n636) );
  XNOR2_X1 U379 ( .A(n370), .B(n537), .ZN(n657) );
  XNOR2_X1 U380 ( .A(n526), .B(KEYINPUT69), .ZN(n541) );
  XNOR2_X1 U381 ( .A(n522), .B(KEYINPUT1), .ZN(n638) );
  NOR2_X2 U382 ( .A1(G902), .A2(n677), .ZN(n424) );
  XNOR2_X1 U383 ( .A(n710), .B(G101), .ZN(n425) );
  NAND2_X1 U384 ( .A1(n372), .A2(n371), .ZN(n635) );
  NAND2_X1 U385 ( .A1(n697), .A2(n373), .ZN(n371) );
  NAND2_X1 U386 ( .A1(n713), .A2(n373), .ZN(n372) );
  XNOR2_X1 U387 ( .A(n540), .B(KEYINPUT42), .ZN(n725) );
  NOR2_X1 U388 ( .A1(n657), .A2(n656), .ZN(n369) );
  NOR2_X1 U389 ( .A1(n568), .A2(n511), .ZN(n631) );
  OR2_X1 U390 ( .A1(n536), .A2(n361), .ZN(n383) );
  XNOR2_X1 U391 ( .A(n587), .B(n405), .ZN(n586) );
  XNOR2_X1 U392 ( .A(n578), .B(n414), .ZN(n723) );
  XOR2_X1 U393 ( .A(G146), .B(G125), .Z(n444) );
  XNOR2_X1 U394 ( .A(n709), .B(G146), .ZN(n408) );
  XNOR2_X1 U395 ( .A(n473), .B(n472), .ZN(n528) );
  XNOR2_X1 U396 ( .A(KEYINPUT103), .B(G478), .ZN(n472) );
  XNOR2_X1 U397 ( .A(n394), .B(n542), .ZN(n555) );
  XOR2_X1 U398 ( .A(KEYINPUT18), .B(KEYINPUT70), .Z(n435) );
  NAND2_X1 U399 ( .A1(n431), .A2(n430), .ZN(n433) );
  XNOR2_X1 U400 ( .A(n476), .B(G116), .ZN(n366) );
  XOR2_X1 U401 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n476) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n477) );
  XNOR2_X1 U403 ( .A(n377), .B(n379), .ZN(n437) );
  XNOR2_X1 U404 ( .A(n448), .B(n380), .ZN(n379) );
  XNOR2_X1 U405 ( .A(n475), .B(n378), .ZN(n377) );
  INV_X1 U406 ( .A(KEYINPUT16), .ZN(n380) );
  NOR2_X1 U407 ( .A1(n723), .A2(n582), .ZN(n413) );
  XOR2_X1 U408 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n488) );
  XNOR2_X1 U409 ( .A(G128), .B(G110), .ZN(n487) );
  XOR2_X1 U410 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n491) );
  XOR2_X1 U411 ( .A(KEYINPUT8), .B(KEYINPUT64), .Z(n465) );
  XNOR2_X1 U412 ( .A(n444), .B(n439), .ZN(n411) );
  INV_X1 U413 ( .A(n586), .ZN(n572) );
  XNOR2_X1 U414 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n460) );
  XNOR2_X1 U415 ( .A(n441), .B(n440), .ZN(n442) );
  AND2_X1 U416 ( .A1(n407), .A2(n586), .ZN(n510) );
  XNOR2_X1 U417 ( .A(n567), .B(KEYINPUT22), .ZN(n579) );
  NAND2_X1 U418 ( .A1(n474), .A2(n535), .ZN(n546) );
  XNOR2_X1 U419 ( .A(n401), .B(n637), .ZN(n400) );
  XNOR2_X1 U420 ( .A(n635), .B(n403), .ZN(n402) );
  INV_X1 U421 ( .A(n469), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n381), .B(G104), .ZN(n448) );
  INV_X1 U423 ( .A(G122), .ZN(n381) );
  INV_X1 U424 ( .A(KEYINPUT48), .ZN(n374) );
  OR2_X1 U425 ( .A1(G237), .A2(G902), .ZN(n509) );
  XNOR2_X1 U426 ( .A(G137), .B(G134), .ZN(n417) );
  XNOR2_X1 U427 ( .A(G122), .B(KEYINPUT7), .ZN(n458) );
  XOR2_X1 U428 ( .A(KEYINPUT102), .B(KEYINPUT100), .Z(n461) );
  XOR2_X1 U429 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n450) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n445) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(G131), .Z(n446) );
  NAND2_X1 U432 ( .A1(G234), .A2(G237), .ZN(n503) );
  XOR2_X1 U433 ( .A(KEYINPUT67), .B(KEYINPUT14), .Z(n504) );
  XOR2_X1 U434 ( .A(G902), .B(KEYINPUT15), .Z(n602) );
  NOR2_X1 U435 ( .A1(n580), .A2(n344), .ZN(n512) );
  XNOR2_X1 U436 ( .A(n571), .B(KEYINPUT68), .ZN(n588) );
  INV_X1 U437 ( .A(KEYINPUT30), .ZN(n519) );
  XNOR2_X1 U438 ( .A(n480), .B(n481), .ZN(n604) );
  XNOR2_X1 U439 ( .A(n475), .B(n366), .ZN(n479) );
  BUF_X1 U440 ( .A(n638), .Z(n367) );
  XNOR2_X1 U441 ( .A(n489), .B(n492), .ZN(n399) );
  XNOR2_X1 U442 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U443 ( .A(n444), .B(n398), .ZN(n708) );
  XNOR2_X1 U444 ( .A(KEYINPUT10), .B(G140), .ZN(n398) );
  XNOR2_X1 U445 ( .A(n481), .B(n422), .ZN(n677) );
  XNOR2_X1 U446 ( .A(G107), .B(G104), .ZN(n421) );
  XNOR2_X1 U447 ( .A(n425), .B(n410), .ZN(n409) );
  XNOR2_X1 U448 ( .A(n411), .B(n427), .ZN(n410) );
  BUF_X1 U449 ( .A(n668), .Z(n363) );
  XNOR2_X1 U450 ( .A(n365), .B(n364), .ZN(n599) );
  INV_X1 U451 ( .A(KEYINPUT79), .ZN(n364) );
  INV_X1 U452 ( .A(n642), .ZN(n396) );
  INV_X1 U453 ( .A(KEYINPUT0), .ZN(n368) );
  INV_X1 U454 ( .A(KEYINPUT6), .ZN(n405) );
  NAND2_X1 U455 ( .A1(n391), .A2(n388), .ZN(n387) );
  AND2_X1 U456 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n683), .A2(n347), .ZN(n391) );
  NAND2_X1 U458 ( .A1(n607), .A2(n406), .ZN(n390) );
  NOR2_X1 U459 ( .A1(n683), .A2(n393), .ZN(n392) );
  INV_X1 U460 ( .A(n607), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n497), .B(n496), .ZN(n690) );
  XNOR2_X1 U462 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U463 ( .A(n399), .B(n708), .ZN(n497) );
  XNOR2_X1 U464 ( .A(G119), .B(G137), .ZN(n494) );
  XNOR2_X1 U465 ( .A(n471), .B(n470), .ZN(n687) );
  INV_X1 U466 ( .A(G134), .ZN(n468) );
  NOR2_X1 U467 ( .A1(n555), .A2(n546), .ZN(n543) );
  INV_X1 U468 ( .A(KEYINPUT36), .ZN(n359) );
  XNOR2_X1 U469 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n384), .B(n349), .ZN(n722) );
  OR2_X1 U471 ( .A1(n579), .A2(n385), .ZN(n384) );
  NAND2_X1 U472 ( .A1(n343), .A2(n570), .ZN(n385) );
  INV_X1 U473 ( .A(KEYINPUT60), .ZN(n352) );
  NAND2_X1 U474 ( .A1(n400), .A2(n357), .ZN(n672) );
  AND2_X1 U475 ( .A1(n671), .A2(n714), .ZN(n357) );
  XNOR2_X1 U476 ( .A(KEYINPUT107), .B(n569), .ZN(n343) );
  OR2_X1 U477 ( .A1(n523), .A2(n642), .ZN(n344) );
  XNOR2_X1 U478 ( .A(n536), .B(KEYINPUT38), .ZN(n653) );
  XNOR2_X1 U479 ( .A(n502), .B(n501), .ZN(n521) );
  OR2_X1 U480 ( .A1(KEYINPUT47), .A2(n548), .ZN(n345) );
  NOR2_X1 U481 ( .A1(n367), .A2(n397), .ZN(n346) );
  XNOR2_X1 U482 ( .A(n543), .B(KEYINPUT40), .ZN(n724) );
  NOR2_X1 U483 ( .A1(n607), .A2(n406), .ZN(n347) );
  XOR2_X1 U484 ( .A(n675), .B(n674), .Z(n348) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n349) );
  XOR2_X1 U486 ( .A(n684), .B(n415), .Z(n350) );
  NOR2_X1 U487 ( .A1(G952), .A2(n714), .ZN(n692) );
  INV_X1 U488 ( .A(n692), .ZN(n389) );
  XNOR2_X1 U489 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n351) );
  INV_X1 U490 ( .A(G472), .ZN(n406) );
  AND2_X1 U491 ( .A1(n512), .A2(n654), .ZN(n407) );
  INV_X1 U492 ( .A(n654), .ZN(n361) );
  XNOR2_X1 U493 ( .A(n353), .B(n352), .ZN(G60) );
  NAND2_X1 U494 ( .A1(n355), .A2(n389), .ZN(n353) );
  XNOR2_X1 U495 ( .A(n354), .B(n351), .ZN(G51) );
  NAND2_X1 U496 ( .A1(n358), .A2(n389), .ZN(n354) );
  XNOR2_X1 U497 ( .A(n685), .B(n350), .ZN(n355) );
  XNOR2_X1 U498 ( .A(n356), .B(n374), .ZN(n404) );
  NAND2_X1 U499 ( .A1(n375), .A2(n376), .ZN(n356) );
  NAND2_X1 U500 ( .A1(n601), .A2(KEYINPUT2), .ZN(n365) );
  XNOR2_X1 U501 ( .A(n369), .B(KEYINPUT41), .ZN(n668) );
  NAND2_X1 U502 ( .A1(n653), .A2(n654), .ZN(n370) );
  XNOR2_X1 U503 ( .A(n676), .B(n348), .ZN(n358) );
  XNOR2_X1 U504 ( .A(n544), .B(KEYINPUT46), .ZN(n375) );
  XNOR2_X1 U505 ( .A(n360), .B(n359), .ZN(n511) );
  NOR2_X1 U506 ( .A1(n549), .A2(n536), .ZN(n360) );
  NAND2_X1 U507 ( .A1(n541), .A2(n653), .ZN(n394) );
  XNOR2_X1 U508 ( .A(n520), .B(n519), .ZN(n525) );
  NAND2_X1 U509 ( .A1(n413), .A2(n722), .ZN(n583) );
  NAND2_X1 U510 ( .A1(n580), .A2(n395), .ZN(n592) );
  NAND2_X1 U511 ( .A1(n412), .A2(n386), .ZN(n362) );
  AND2_X1 U512 ( .A1(n545), .A2(n345), .ZN(n376) );
  INV_X1 U513 ( .A(n590), .ZN(n574) );
  NAND2_X1 U514 ( .A1(n590), .A2(n566), .ZN(n567) );
  XNOR2_X2 U515 ( .A(n382), .B(n368), .ZN(n590) );
  NOR2_X1 U516 ( .A1(n612), .A2(n594), .ZN(n595) );
  NOR2_X2 U517 ( .A1(n585), .A2(n586), .ZN(n612) );
  NAND2_X1 U518 ( .A1(n700), .A2(n438), .ZN(n412) );
  XNOR2_X2 U519 ( .A(n598), .B(KEYINPUT45), .ZN(n697) );
  INV_X1 U520 ( .A(KEYINPUT2), .ZN(n373) );
  INV_X1 U521 ( .A(n437), .ZN(n700) );
  NAND2_X1 U522 ( .A1(n565), .A2(n564), .ZN(n382) );
  NOR2_X2 U523 ( .A1(n675), .A2(n602), .ZN(n443) );
  NAND2_X1 U524 ( .A1(n437), .A2(n436), .ZN(n386) );
  AND2_X2 U525 ( .A1(n603), .A2(n636), .ZN(n683) );
  AND2_X1 U526 ( .A1(n522), .A2(n396), .ZN(n395) );
  NOR2_X1 U527 ( .A1(n521), .A2(n642), .ZN(n397) );
  NAND2_X1 U528 ( .A1(n397), .A2(n638), .ZN(n571) );
  NAND2_X1 U529 ( .A1(n402), .A2(n636), .ZN(n401) );
  INV_X1 U530 ( .A(KEYINPUT74), .ZN(n403) );
  AND2_X2 U531 ( .A1(n404), .A2(n558), .ZN(n601) );
  XNOR2_X2 U532 ( .A(n482), .B(n406), .ZN(n587) );
  NAND2_X1 U533 ( .A1(n683), .A2(G475), .ZN(n685) );
  NOR2_X1 U534 ( .A1(n635), .A2(n483), .ZN(n603) );
  NOR2_X2 U535 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U536 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n415) );
  INV_X1 U537 ( .A(n634), .ZN(n557) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  AND2_X1 U539 ( .A1(n721), .A2(n557), .ZN(n558) );
  INV_X1 U540 ( .A(KEYINPUT93), .ZN(n490) );
  XNOR2_X1 U541 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n513) );
  INV_X1 U542 ( .A(KEYINPUT78), .ZN(n600) );
  INV_X1 U543 ( .A(KEYINPUT77), .ZN(n637) );
  XNOR2_X1 U544 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U545 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X2 U546 ( .A(n416), .B(G128), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n417), .B(G131), .ZN(n709) );
  XOR2_X1 U548 ( .A(KEYINPUT66), .B(G110), .Z(n426) );
  XOR2_X1 U549 ( .A(G140), .B(n426), .Z(n419) );
  NAND2_X1 U550 ( .A1(G227), .A2(n714), .ZN(n418) );
  XNOR2_X1 U551 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U552 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U553 ( .A(KEYINPUT65), .B(G469), .ZN(n423) );
  XNOR2_X2 U554 ( .A(n424), .B(n423), .ZN(n522) );
  XNOR2_X1 U555 ( .A(KEYINPUT85), .B(n638), .ZN(n568) );
  INV_X1 U556 ( .A(n426), .ZN(n427) );
  INV_X1 U557 ( .A(G119), .ZN(n428) );
  NAND2_X1 U558 ( .A1(n428), .A2(G113), .ZN(n431) );
  INV_X1 U559 ( .A(G113), .ZN(n429) );
  NAND2_X1 U560 ( .A1(n429), .A2(G119), .ZN(n430) );
  XOR2_X1 U561 ( .A(G116), .B(G107), .Z(n469) );
  NAND2_X1 U562 ( .A1(G224), .A2(n714), .ZN(n434) );
  XOR2_X1 U563 ( .A(n435), .B(n434), .Z(n438) );
  INV_X1 U564 ( .A(n438), .ZN(n436) );
  XNOR2_X1 U565 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n439) );
  NAND2_X1 U566 ( .A1(G210), .A2(n509), .ZN(n441) );
  INV_X1 U567 ( .A(KEYINPUT88), .ZN(n440) );
  XNOR2_X2 U568 ( .A(n443), .B(n442), .ZN(n536) );
  XNOR2_X1 U569 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n456) );
  XNOR2_X1 U570 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U571 ( .A(n708), .B(n447), .ZN(n454) );
  XNOR2_X1 U572 ( .A(n448), .B(KEYINPUT11), .ZN(n452) );
  NAND2_X1 U573 ( .A1(G214), .A2(n477), .ZN(n449) );
  XNOR2_X1 U574 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U575 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U576 ( .A(n454), .B(n453), .ZN(n684) );
  NOR2_X1 U577 ( .A1(G902), .A2(n684), .ZN(n455) );
  XNOR2_X1 U578 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U579 ( .A(G475), .B(n457), .ZN(n534) );
  INV_X1 U580 ( .A(n534), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n459), .B(n458), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U583 ( .A(n463), .B(n462), .Z(n467) );
  NAND2_X1 U584 ( .A1(G234), .A2(n714), .ZN(n464) );
  XNOR2_X1 U585 ( .A(n465), .B(n464), .ZN(n493) );
  NAND2_X1 U586 ( .A1(n493), .A2(G217), .ZN(n466) );
  XNOR2_X1 U587 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U589 ( .A1(n687), .A2(G902), .ZN(n473) );
  INV_X1 U590 ( .A(n528), .ZN(n535) );
  INV_X1 U591 ( .A(n546), .ZN(n626) );
  NAND2_X1 U592 ( .A1(n477), .A2(G210), .ZN(n478) );
  XOR2_X1 U593 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n486) );
  INV_X1 U594 ( .A(n602), .ZN(n483) );
  NAND2_X1 U595 ( .A1(G234), .A2(n483), .ZN(n484) );
  XNOR2_X1 U596 ( .A(KEYINPUT20), .B(n484), .ZN(n498) );
  NAND2_X1 U597 ( .A1(n498), .A2(G221), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n486), .B(n485), .ZN(n642) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U600 ( .A1(G221), .A2(n493), .ZN(n495) );
  NOR2_X1 U601 ( .A1(n690), .A2(G902), .ZN(n502) );
  XOR2_X1 U602 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n500) );
  NAND2_X1 U603 ( .A1(n498), .A2(G217), .ZN(n499) );
  XNOR2_X1 U604 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U605 ( .A(n521), .ZN(n580) );
  XNOR2_X1 U606 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U607 ( .A1(G952), .A2(n505), .ZN(n666) );
  NOR2_X1 U608 ( .A1(G953), .A2(n666), .ZN(n562) );
  NAND2_X1 U609 ( .A1(G902), .A2(n505), .ZN(n560) );
  OR2_X1 U610 ( .A1(n714), .A2(n560), .ZN(n506) );
  NOR2_X1 U611 ( .A1(G900), .A2(n506), .ZN(n507) );
  NOR2_X1 U612 ( .A1(n562), .A2(n507), .ZN(n508) );
  XOR2_X1 U613 ( .A(KEYINPUT73), .B(n508), .Z(n523) );
  NAND2_X1 U614 ( .A1(G214), .A2(n509), .ZN(n654) );
  NAND2_X1 U615 ( .A1(n626), .A2(n510), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n631), .B(KEYINPUT81), .ZN(n518) );
  INV_X1 U617 ( .A(n536), .ZN(n553) );
  INV_X1 U618 ( .A(n522), .ZN(n516) );
  NAND2_X1 U619 ( .A1(n512), .A2(n587), .ZN(n514) );
  NOR2_X1 U620 ( .A1(n516), .A2(n515), .ZN(n538) );
  NAND2_X1 U621 ( .A1(n565), .A2(n538), .ZN(n547) );
  NAND2_X1 U622 ( .A1(KEYINPUT47), .A2(n547), .ZN(n517) );
  NAND2_X1 U623 ( .A1(n518), .A2(n517), .ZN(n533) );
  NAND2_X1 U624 ( .A1(n587), .A2(n654), .ZN(n520) );
  NOR2_X1 U625 ( .A1(n592), .A2(n523), .ZN(n524) );
  NAND2_X1 U626 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U627 ( .A1(n535), .A2(n534), .ZN(n576) );
  AND2_X1 U628 ( .A1(n553), .A2(n576), .ZN(n527) );
  NAND2_X1 U629 ( .A1(n541), .A2(n527), .ZN(n624) );
  XNOR2_X1 U630 ( .A(n624), .B(KEYINPUT76), .ZN(n530) );
  NAND2_X1 U631 ( .A1(n528), .A2(n534), .ZN(n556) );
  INV_X1 U632 ( .A(n556), .ZN(n628) );
  NOR2_X1 U633 ( .A1(n626), .A2(n628), .ZN(n658) );
  NAND2_X1 U634 ( .A1(KEYINPUT47), .A2(n658), .ZN(n529) );
  NAND2_X1 U635 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U636 ( .A(KEYINPUT75), .B(n531), .Z(n532) );
  NOR2_X1 U637 ( .A1(n533), .A2(n532), .ZN(n545) );
  NAND2_X1 U638 ( .A1(n535), .A2(n534), .ZN(n656) );
  INV_X1 U639 ( .A(KEYINPUT111), .ZN(n537) );
  INV_X1 U640 ( .A(n538), .ZN(n539) );
  NOR2_X1 U641 ( .A1(n668), .A2(n539), .ZN(n540) );
  INV_X1 U642 ( .A(KEYINPUT39), .ZN(n542) );
  NOR2_X1 U643 ( .A1(n546), .A2(n547), .ZN(n625) );
  NOR2_X1 U644 ( .A1(n556), .A2(n547), .ZN(n622) );
  NOR2_X1 U645 ( .A1(n625), .A2(n622), .ZN(n548) );
  NOR2_X1 U646 ( .A1(n367), .A2(n549), .ZN(n551) );
  XNOR2_X1 U647 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n550) );
  XNOR2_X1 U648 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U649 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U650 ( .A(n554), .B(KEYINPUT109), .ZN(n721) );
  NOR2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n634) );
  XNOR2_X1 U652 ( .A(n572), .B(KEYINPUT72), .ZN(n570) );
  NOR2_X1 U653 ( .A1(n642), .A2(n656), .ZN(n559) );
  XNOR2_X1 U654 ( .A(KEYINPUT104), .B(n559), .ZN(n566) );
  XNOR2_X1 U655 ( .A(G898), .B(KEYINPUT89), .ZN(n695) );
  NAND2_X1 U656 ( .A1(G953), .A2(n695), .ZN(n703) );
  NOR2_X1 U657 ( .A1(n703), .A2(n560), .ZN(n561) );
  NOR2_X1 U658 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U659 ( .A(KEYINPUT90), .B(n563), .Z(n564) );
  XOR2_X1 U660 ( .A(n580), .B(KEYINPUT105), .Z(n640) );
  OR2_X1 U661 ( .A1(n568), .A2(n640), .ZN(n569) );
  NOR2_X1 U662 ( .A1(n588), .A2(n572), .ZN(n573) );
  XNOR2_X1 U663 ( .A(n573), .B(KEYINPUT33), .ZN(n667) );
  XNOR2_X1 U664 ( .A(n575), .B(KEYINPUT34), .ZN(n577) );
  NAND2_X1 U665 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U666 ( .A1(n587), .A2(n580), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n584), .A2(n581), .ZN(n621) );
  INV_X1 U668 ( .A(n621), .ZN(n582) );
  XNOR2_X1 U669 ( .A(n583), .B(KEYINPUT44), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n640), .A2(n584), .ZN(n585) );
  INV_X1 U671 ( .A(n587), .ZN(n645) );
  NOR2_X1 U672 ( .A1(n588), .A2(n645), .ZN(n649) );
  NAND2_X1 U673 ( .A1(n590), .A2(n649), .ZN(n589) );
  XNOR2_X1 U674 ( .A(n589), .B(KEYINPUT31), .ZN(n629) );
  NAND2_X1 U675 ( .A1(n590), .A2(n645), .ZN(n591) );
  NOR2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n618) );
  NOR2_X1 U677 ( .A1(n629), .A2(n618), .ZN(n593) );
  NOR2_X1 U678 ( .A1(n658), .A2(n593), .ZN(n594) );
  XOR2_X1 U679 ( .A(KEYINPUT106), .B(n595), .Z(n596) );
  XOR2_X1 U680 ( .A(n604), .B(KEYINPUT62), .Z(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT84), .B(KEYINPUT112), .Z(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT82), .B(KEYINPUT113), .Z(n609) );
  XNOR2_X1 U683 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n609), .B(n608), .ZN(n610) );
  XOR2_X1 U685 ( .A(n611), .B(n610), .Z(G57) );
  XOR2_X1 U686 ( .A(n612), .B(G101), .Z(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT114), .B(n613), .ZN(G3) );
  NAND2_X1 U688 ( .A1(n618), .A2(n626), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(G104), .ZN(G6) );
  XOR2_X1 U690 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n616) );
  XNOR2_X1 U691 ( .A(G107), .B(KEYINPUT26), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n616), .B(n615), .ZN(n617) );
  XOR2_X1 U693 ( .A(KEYINPUT115), .B(n617), .Z(n620) );
  NAND2_X1 U694 ( .A1(n618), .A2(n628), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n620), .B(n619), .ZN(G9) );
  XNOR2_X1 U696 ( .A(G110), .B(n621), .ZN(G12) );
  XNOR2_X1 U697 ( .A(G128), .B(n622), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT29), .ZN(G30) );
  XNOR2_X1 U699 ( .A(G143), .B(n624), .ZN(G45) );
  XOR2_X1 U700 ( .A(G146), .B(n625), .Z(G48) );
  NAND2_X1 U701 ( .A1(n629), .A2(n626), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(G113), .ZN(G15) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(G116), .ZN(G18) );
  XOR2_X1 U705 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n633) );
  XNOR2_X1 U706 ( .A(n631), .B(G125), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n633), .B(n632), .ZN(G27) );
  XOR2_X1 U708 ( .A(G134), .B(n634), .Z(G36) );
  XOR2_X1 U709 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n673) );
  XNOR2_X1 U710 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n346), .B(n639), .ZN(n647) );
  INV_X1 U712 ( .A(n640), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U714 ( .A(KEYINPUT49), .B(n643), .Z(n644) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT119), .ZN(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT51), .B(n651), .ZN(n652) );
  NOR2_X1 U720 ( .A1(n363), .A2(n652), .ZN(n663) );
  NOR2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U722 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n661), .A2(n667), .ZN(n662) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U727 ( .A(n664), .B(KEYINPUT52), .ZN(n665) );
  NOR2_X1 U728 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U729 ( .A1(n363), .A2(n667), .ZN(n669) );
  NOR2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n673), .B(n672), .ZN(G75) );
  NAND2_X1 U732 ( .A1(n683), .A2(G210), .ZN(n676) );
  XOR2_X1 U733 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n674) );
  XNOR2_X1 U734 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n677), .B(KEYINPUT57), .ZN(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U737 ( .A1(n683), .A2(G469), .ZN(n680) );
  XOR2_X1 U738 ( .A(n681), .B(n680), .Z(n682) );
  NOR2_X1 U739 ( .A1(n692), .A2(n682), .ZN(G54) );
  NAND2_X1 U740 ( .A1(G478), .A2(n683), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U742 ( .A1(n692), .A2(n688), .ZN(G63) );
  NAND2_X1 U743 ( .A1(G217), .A2(n683), .ZN(n689) );
  XNOR2_X1 U744 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n692), .A2(n691), .ZN(G66) );
  XNOR2_X1 U746 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n707) );
  XOR2_X1 U747 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n694) );
  NAND2_X1 U748 ( .A1(G224), .A2(G953), .ZN(n693) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U751 ( .A1(G953), .A2(n697), .ZN(n698) );
  NOR2_X1 U752 ( .A1(n699), .A2(n698), .ZN(n705) );
  XNOR2_X1 U753 ( .A(n700), .B(G101), .ZN(n701) );
  XNOR2_X1 U754 ( .A(n701), .B(G110), .ZN(n702) );
  NAND2_X1 U755 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U756 ( .A(n705), .B(n704), .Z(n706) );
  XNOR2_X1 U757 ( .A(n707), .B(n706), .ZN(G69) );
  XNOR2_X1 U758 ( .A(n708), .B(KEYINPUT127), .ZN(n712) );
  XNOR2_X1 U759 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U760 ( .A(n712), .B(n711), .ZN(n716) );
  XNOR2_X1 U761 ( .A(n716), .B(n713), .ZN(n715) );
  NAND2_X1 U762 ( .A1(n715), .A2(n714), .ZN(n720) );
  XNOR2_X1 U763 ( .A(G227), .B(n716), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(G900), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n718), .A2(G953), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n720), .A2(n719), .ZN(G72) );
  XNOR2_X1 U767 ( .A(G140), .B(n721), .ZN(G42) );
  XNOR2_X1 U768 ( .A(G119), .B(n722), .ZN(G21) );
  XOR2_X1 U769 ( .A(n723), .B(G122), .Z(G24) );
  XOR2_X1 U770 ( .A(G131), .B(n724), .Z(G33) );
  XOR2_X1 U771 ( .A(n725), .B(G137), .Z(G39) );
endmodule

