//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT73), .B(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G113gat), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G127gat), .ZN(new_n209));
  INV_X1    g008(.A(G127gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n207), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  OR3_X1    g014(.A1(new_n215), .A2(KEYINPUT84), .A3(G148gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT84), .B1(new_n215), .B2(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(G148gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n223), .B2(KEYINPUT2), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  INV_X1    g024(.A(G148gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G141gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n218), .B2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n223), .A2(new_n220), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n219), .A2(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT71), .B1(new_n210), .B2(G134gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n208), .A3(G127gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(G134gat), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT1), .B1(new_n203), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n230), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT4), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n214), .A2(new_n230), .A3(new_n243), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n230), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n243), .B1(new_n206), .B2(new_n213), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n245), .A2(KEYINPUT85), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n247), .A2(KEYINPUT86), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n206), .A2(new_n213), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n241), .B1(new_n237), .B2(new_n234), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n246), .A4(new_n230), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n267), .A3(KEYINPUT4), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n260), .A2(new_n261), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n255), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n244), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n264), .A2(new_n230), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n256), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n259), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT0), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT87), .ZN(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G85gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT89), .B(KEYINPUT6), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  INV_X1    g086(.A(new_n284), .ZN(new_n288));
  INV_X1    g087(.A(new_n268), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n267), .B1(new_n244), .B2(KEYINPUT4), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n261), .A2(new_n266), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n270), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n288), .B(new_n258), .C1(new_n293), .C2(new_n276), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n278), .A2(KEYINPUT88), .A3(new_n288), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n278), .A2(new_n288), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G226gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT69), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT26), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n305), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n309), .A2(new_n310), .B1(new_n304), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n306), .A2(new_n308), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT70), .B1(new_n314), .B2(new_n304), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n313), .A2(new_n315), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n324));
  INV_X1    g123(.A(G183gat), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n325), .A2(KEYINPUT27), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(KEYINPUT27), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n322), .A2(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n319), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(G183gat), .B2(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(KEYINPUT24), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT23), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n340), .A2(new_n342), .A3(new_n311), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT25), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n342), .A3(new_n311), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(new_n325), .A3(new_n319), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n337), .B(KEYINPUT24), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n351), .B2(KEYINPUT25), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n333), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n301), .B1(new_n353), .B2(KEYINPUT29), .ZN(new_n354));
  INV_X1    g153(.A(G204gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G197gat), .ZN(new_n356));
  INV_X1    g155(.A(G197gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G204gat), .ZN(new_n358));
  INV_X1    g157(.A(G211gat), .ZN(new_n359));
  INV_X1    g158(.A(G218gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n356), .B(new_n358), .C1(new_n361), .C2(KEYINPUT22), .ZN(new_n362));
  XOR2_X1   g161(.A(G211gat), .B(G218gat), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n348), .B(new_n347), .C1(new_n336), .C2(new_n338), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT25), .B1(new_n366), .B2(new_n343), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT25), .A4(new_n311), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n350), .B2(new_n334), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n344), .B(KEYINPUT66), .C1(new_n351), .C2(KEYINPUT25), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n333), .ZN(new_n373));
  INV_X1    g172(.A(new_n301), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT82), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n370), .A2(new_n371), .B1(new_n316), .B2(new_n332), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n301), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n354), .A2(new_n364), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n333), .A2(new_n352), .A3(new_n374), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n364), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n301), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n384), .B(new_n386), .C1(new_n377), .C2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n379), .B(new_n383), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT30), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n389), .B(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n379), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n382), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT90), .B1(new_n300), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n404));
  INV_X1    g203(.A(new_n286), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT88), .B1(new_n278), .B2(new_n288), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n276), .B1(new_n269), .B2(new_n271), .ZN(new_n407));
  NOR4_X1   g206(.A1(new_n407), .A2(new_n295), .A3(new_n284), .A4(new_n259), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n285), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n299), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT31), .B(G50gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n364), .A2(new_n387), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n230), .B1(new_n417), .B2(new_n251), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G228gat), .ZN(new_n420));
  INV_X1    g219(.A(G233gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT29), .B1(new_n230), .B2(new_n251), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n364), .B(KEYINPUT80), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n419), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n364), .ZN(new_n426));
  OAI22_X1  g225(.A1(new_n418), .A2(new_n426), .B1(new_n420), .B2(new_n421), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n416), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n425), .A2(new_n416), .A3(new_n427), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n415), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  INV_X1    g231(.A(new_n415), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n432), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n414), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n432), .B2(new_n428), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n430), .A3(new_n415), .ZN(new_n437));
  INV_X1    g236(.A(new_n414), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n403), .A2(new_n413), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n373), .A2(new_n264), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n377), .A2(new_n253), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n443), .A2(KEYINPUT77), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT77), .B1(new_n443), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n442), .B(KEYINPUT64), .Z(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n447), .A2(KEYINPUT34), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(G15gat), .B(G43gat), .Z(new_n453));
  XNOR2_X1  g252(.A(G71gat), .B(G99gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n443), .A2(new_n444), .A3(new_n449), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(KEYINPUT32), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n458), .A2(KEYINPUT75), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT75), .B1(new_n458), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n457), .B(KEYINPUT32), .C1(new_n459), .C2(new_n456), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT76), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n452), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n460), .A2(new_n468), .A3(new_n455), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT75), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n458), .A2(KEYINPUT75), .A3(new_n460), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n464), .B(KEYINPUT76), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n451), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n467), .A2(KEYINPUT36), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT78), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT78), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n467), .A2(new_n478), .A3(KEYINPUT36), .A4(new_n475), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n451), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(new_n475), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n441), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n255), .B1(new_n248), .B2(new_n254), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n273), .A2(new_n274), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n490), .B(KEYINPUT39), .C1(new_n256), .C2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n288), .C1(KEYINPUT39), .C2(new_n490), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT40), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n410), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n440), .B1(new_n497), .B2(new_n402), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n399), .A2(new_n499), .A3(new_n379), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n382), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(KEYINPUT38), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n354), .A2(new_n378), .A3(new_n375), .ZN(new_n503));
  INV_X1    g302(.A(new_n364), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT91), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n384), .B1(new_n377), .B2(new_n388), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n424), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n505), .A2(KEYINPUT91), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n499), .B1(new_n399), .B2(new_n379), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT38), .B1(new_n501), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n512), .A2(new_n300), .A3(new_n514), .A4(new_n393), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT92), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n498), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n488), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n403), .A2(new_n413), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n473), .A2(new_n474), .A3(new_n451), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n440), .A2(new_n523), .A3(new_n482), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n485), .A2(new_n440), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n300), .A2(new_n402), .A3(KEYINPUT35), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G43gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT15), .B1(new_n532), .B2(G50gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n532), .B2(G50gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(G29gat), .B2(G36gat), .ZN(new_n535));
  OR3_X1    g334(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT95), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(KEYINPUT95), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT94), .B(G43gat), .ZN(new_n542));
  INV_X1    g341(.A(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n532), .A2(G50gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT15), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  OAI22_X1  g348(.A1(new_n538), .A2(KEYINPUT93), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n538), .A2(KEYINPUT93), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n534), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(G1gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n557), .B(new_n558), .C1(G1gat), .C2(new_n555), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n553), .B(KEYINPUT17), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(KEYINPUT18), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n553), .A2(KEYINPUT17), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n553), .A2(KEYINPUT17), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n562), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n553), .B(new_n561), .Z(new_n574));
  XOR2_X1   g373(.A(new_n565), .B(KEYINPUT13), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n566), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT11), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n302), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G197gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT12), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n566), .A2(new_n573), .A3(new_n576), .A4(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n531), .A2(KEYINPUT97), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n488), .A2(new_n520), .B1(new_n526), .B2(new_n529), .ZN(new_n589));
  INV_X1    g388(.A(new_n586), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G57gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT100), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT99), .B(G57gat), .Z(new_n596));
  OAI21_X1  g395(.A(new_n595), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n600), .A2(new_n601), .B1(new_n602), .B2(new_n599), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n597), .B(new_n603), .C1(new_n601), .C2(new_n600), .ZN(new_n604));
  XNOR2_X1  g403(.A(G57gat), .B(G64gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n599), .B(new_n598), .C1(new_n605), .C2(new_n602), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT21), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT102), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT21), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n561), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT103), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n621), .A2(new_n622), .A3(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT104), .ZN(new_n635));
  NAND2_X1  g434(.A1(G85gat), .A2(G92gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT7), .ZN(new_n637));
  INV_X1    g436(.A(G99gat), .ZN(new_n638));
  INV_X1    g437(.A(G106gat), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT8), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n637), .B(new_n640), .C1(G85gat), .C2(G92gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n635), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n563), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n563), .A2(KEYINPUT105), .A3(new_n642), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n554), .B2(new_n642), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n633), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n645), .B2(new_n646), .ZN(new_n652));
  INV_X1    g451(.A(new_n633), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n656));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n651), .B(new_n654), .C1(new_n655), .C2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n655), .B1(new_n652), .B2(new_n653), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n652), .A2(new_n653), .ZN(new_n662));
  AOI211_X1 g461(.A(new_n650), .B(new_n633), .C1(new_n645), .C2(new_n646), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n661), .B(new_n658), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n624), .A2(new_n642), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n624), .A2(new_n642), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n624), .A2(new_n642), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n674), .A2(KEYINPUT10), .B1(new_n624), .B2(new_n642), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n666), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G120gat), .B(G148gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n671), .A2(new_n684), .A3(new_n678), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n632), .A2(new_n665), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n592), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n300), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G1gat), .ZN(new_n690));
  INV_X1    g489(.A(G1gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n691), .A3(new_n300), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1324gat));
  NAND3_X1  g492(.A1(new_n592), .A2(new_n402), .A3(new_n687), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n688), .A2(new_n402), .A3(new_n695), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n694), .B2(G8gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(new_n485), .ZN(new_n702));
  AOI21_X1  g501(.A(G15gat), .B1(new_n688), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n523), .B1(new_n483), .B2(new_n482), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT36), .B1(new_n705), .B2(new_n481), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n477), .A2(new_n479), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n487), .A2(KEYINPUT109), .A3(new_n477), .A4(new_n479), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G15gat), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT110), .Z(new_n712));
  AOI21_X1  g511(.A(new_n703), .B1(new_n688), .B2(new_n712), .ZN(G1326gat));
  NAND3_X1  g512(.A1(new_n592), .A2(new_n440), .A3(new_n687), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NOR2_X1   g515(.A1(new_n631), .A2(new_n686), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n665), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n587), .B2(new_n591), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n411), .A2(G29gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n719), .A2(KEYINPUT45), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n717), .A2(new_n586), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n403), .A2(new_n413), .A3(new_n440), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT111), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n403), .A2(new_n413), .A3(new_n728), .A4(new_n440), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n498), .A2(new_n515), .A3(new_n518), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n518), .B1(new_n498), .B2(new_n515), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n727), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n530), .B1(new_n710), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n665), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n660), .A2(new_n664), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n589), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n411), .B(new_n725), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n723), .B(new_n724), .C1(new_n738), .C2(new_n548), .ZN(G1328gat));
  NOR2_X1   g538(.A1(new_n404), .A2(G36gat), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n719), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT46), .B1(new_n719), .B2(new_n740), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n404), .B(new_n725), .C1(new_n735), .C2(new_n737), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n741), .A2(new_n742), .B1(new_n549), .B2(new_n743), .ZN(G1329gat));
  NAND2_X1  g543(.A1(new_n710), .A2(new_n542), .ZN(new_n745));
  AOI211_X1 g544(.A(new_n725), .B(new_n745), .C1(new_n735), .C2(new_n737), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  INV_X1    g547(.A(new_n718), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n592), .A2(new_n702), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n747), .B(new_n748), .C1(new_n751), .C2(new_n542), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n542), .B1(new_n719), .B2(new_n702), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT47), .B1(new_n753), .B2(new_n746), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1330gat));
  NAND2_X1  g554(.A1(new_n719), .A2(new_n440), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n543), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  INV_X1    g557(.A(new_n440), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n543), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n725), .B(new_n761), .C1(new_n735), .C2(new_n737), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(G50gat), .B1(new_n719), .B2(new_n440), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT48), .B1(new_n765), .B2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1331gat));
  INV_X1    g566(.A(new_n686), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n632), .A2(new_n586), .A3(new_n665), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n733), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n300), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(new_n596), .ZN(G1332gat));
  AOI21_X1  g571(.A(new_n404), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT113), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n774), .B(new_n776), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n770), .A2(new_n778), .A3(new_n702), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n733), .A2(new_n710), .A3(new_n769), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n770), .A2(new_n440), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  AOI22_X1  g584(.A1(new_n517), .A2(new_n519), .B1(new_n441), .B2(new_n728), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(new_n708), .A3(new_n709), .A4(new_n727), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n736), .B1(new_n787), .B2(new_n530), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n631), .B2(new_n586), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n629), .A2(KEYINPUT115), .A3(new_n590), .A4(new_n630), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT51), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n665), .A4(new_n792), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n300), .B(new_n686), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(G85gat), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT116), .B1(new_n792), .B2(new_n686), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n799), .B(new_n768), .C1(new_n790), .C2(new_n791), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n735), .B2(new_n737), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n411), .A2(new_n797), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n796), .A2(new_n797), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NOR2_X1   g603(.A1(new_n404), .A2(G92gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n733), .A2(new_n665), .A3(new_n792), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n768), .B(new_n806), .C1(new_n809), .C2(new_n794), .ZN(new_n810));
  INV_X1    g609(.A(G92gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n802), .B2(new_n402), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n735), .A2(new_n737), .ZN(new_n814));
  INV_X1    g613(.A(new_n801), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n402), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n686), .B(new_n805), .C1(new_n793), .C2(new_n795), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n820), .ZN(G1337gat));
  OAI211_X1 g620(.A(new_n702), .B(new_n686), .C1(new_n793), .C2(new_n795), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n638), .B1(new_n708), .B2(new_n709), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n822), .A2(new_n638), .B1(new_n802), .B2(new_n823), .ZN(G1338gat));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n440), .A2(new_n639), .A3(new_n686), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT117), .Z(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n793), .B2(new_n795), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n802), .A2(new_n440), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n825), .B(new_n828), .C1(new_n829), .C2(new_n639), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n639), .B1(new_n802), .B2(new_n440), .ZN(new_n831));
  INV_X1    g630(.A(new_n827), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n809), .B2(new_n794), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT53), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n834), .ZN(G1339gat));
  NAND4_X1  g634(.A1(new_n631), .A2(new_n736), .A3(new_n590), .A4(new_n768), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n564), .A2(new_n565), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n574), .A2(new_n575), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n581), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n585), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n686), .ZN(new_n841));
  INV_X1    g640(.A(new_n685), .ZN(new_n842));
  XOR2_X1   g641(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n843));
  NAND4_X1  g642(.A1(new_n675), .A2(new_n677), .A3(new_n666), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n678), .A2(KEYINPUT54), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n666), .B1(new_n675), .B2(new_n677), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n682), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n844), .A2(new_n682), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(KEYINPUT55), .C1(new_n846), .C2(new_n845), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n841), .B1(new_n590), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n585), .A2(new_n839), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n660), .B2(new_n664), .ZN(new_n855));
  INV_X1    g654(.A(new_n852), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n736), .A2(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n836), .B1(new_n857), .B2(new_n631), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n858), .A2(new_n300), .A3(new_n404), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n524), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n586), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n527), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n202), .A3(new_n590), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n863), .ZN(G1340gat));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n205), .A3(new_n686), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n862), .B2(new_n768), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  NAND4_X1  g666(.A1(new_n860), .A2(new_n235), .A3(new_n236), .A4(new_n631), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n235), .A2(new_n236), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n862), .B2(new_n632), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1342gat));
  NAND4_X1  g670(.A1(new_n859), .A2(new_n208), .A3(new_n524), .A4(new_n665), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT56), .Z(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n862), .B2(new_n736), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n849), .A2(new_n877), .A3(new_n851), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n849), .B2(new_n851), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n586), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n665), .B1(new_n880), .B2(new_n841), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n665), .A2(new_n856), .A3(new_n840), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n632), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n836), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n876), .B1(new_n885), .B2(new_n440), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n858), .A2(new_n876), .A3(new_n440), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n710), .A2(new_n411), .A3(new_n402), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(G141gat), .A3(new_n586), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n710), .A2(new_n759), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n859), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n215), .B1(new_n893), .B2(new_n590), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n891), .A2(KEYINPUT58), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n853), .A2(new_n736), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n631), .B1(new_n901), .B2(new_n882), .ZN(new_n902));
  AND4_X1   g701(.A1(new_n590), .A2(new_n631), .A3(new_n736), .A4(new_n768), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT57), .B(new_n440), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n858), .A2(new_n906), .A3(KEYINPUT57), .A4(new_n440), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n759), .B1(new_n884), .B2(new_n836), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n905), .B(new_n907), .C1(new_n908), .C2(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n686), .A3(new_n888), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n900), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT59), .B(new_n226), .C1(new_n890), .C2(new_n686), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n686), .A2(new_n226), .ZN(new_n913));
  OAI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n893), .B2(new_n913), .ZN(G1345gat));
  NOR2_X1   g713(.A1(new_n893), .A2(new_n632), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n916));
  AOI21_X1  g715(.A(G155gat), .B1(new_n915), .B2(KEYINPUT121), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n632), .A2(new_n221), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n916), .A2(new_n917), .B1(new_n890), .B2(new_n918), .ZN(G1346gat));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n886), .A2(new_n889), .A3(new_n736), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n222), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n665), .A2(new_n222), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n893), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI221_X1 g724(.A(KEYINPUT122), .B1(new_n893), .B2(new_n923), .C1(new_n921), .C2(new_n222), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n404), .A2(new_n300), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n858), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n524), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n302), .B1(new_n930), .B2(new_n590), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n858), .A2(new_n527), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(G169gat), .A3(new_n586), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT123), .ZN(G1348gat));
  NAND3_X1  g734(.A1(new_n932), .A2(G176gat), .A3(new_n686), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  INV_X1    g736(.A(new_n930), .ZN(new_n938));
  AOI21_X1  g737(.A(G176gat), .B1(new_n938), .B2(new_n686), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(G1349gat));
  NOR2_X1   g739(.A1(new_n632), .A2(new_n330), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n929), .A2(new_n524), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n932), .A2(new_n631), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G183gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n942), .A2(new_n943), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n944), .A2(new_n946), .A3(new_n950), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  AOI21_X1  g751(.A(new_n319), .B1(new_n932), .B2(new_n665), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT61), .Z(new_n954));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n319), .A3(new_n665), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n710), .A2(new_n300), .A3(new_n404), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n909), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n958), .A2(new_n357), .A3(new_n590), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n929), .A2(new_n892), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n586), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n959), .A2(new_n962), .ZN(G1352gat));
  NAND3_X1  g762(.A1(new_n909), .A2(new_n686), .A3(new_n957), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n686), .A2(new_n355), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT62), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n960), .A2(KEYINPUT62), .A3(new_n966), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n965), .B(new_n967), .C1(new_n969), .C2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n909), .A2(new_n631), .A3(new_n957), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G211gat), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT63), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n975), .A3(G211gat), .ZN(new_n976));
  AND4_X1   g775(.A1(new_n359), .A2(new_n929), .A3(new_n631), .A4(new_n892), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n974), .A2(new_n976), .A3(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n958), .B2(new_n736), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n360), .A3(new_n665), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


