

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n641), .A2(n640), .ZN(n644) );
  OR2_X1 U553 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U554 ( .A1(G651), .A2(n598), .ZN(n791) );
  NOR2_X1 U555 ( .A1(n562), .A2(n561), .ZN(G160) );
  AND2_X1 U556 ( .A1(G54), .A2(n791), .ZN(n518) );
  AND2_X1 U557 ( .A1(n944), .A2(n704), .ZN(n519) );
  NOR2_X1 U558 ( .A1(n701), .A2(n698), .ZN(n520) );
  OR2_X1 U559 ( .A1(n701), .A2(n691), .ZN(n521) );
  AND2_X1 U560 ( .A1(n707), .A2(n706), .ZN(n522) );
  OR2_X1 U561 ( .A1(n681), .A2(n657), .ZN(n658) );
  INV_X1 U562 ( .A(n670), .ZN(n651) );
  INV_X1 U563 ( .A(KEYINPUT102), .ZN(n660) );
  AND2_X1 U564 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U565 ( .A(n650), .B(KEYINPUT29), .ZN(n655) );
  INV_X1 U566 ( .A(KEYINPUT103), .ZN(n668) );
  NAND2_X1 U567 ( .A1(G8), .A2(n670), .ZN(n701) );
  NOR2_X1 U568 ( .A1(n632), .A2(n518), .ZN(n633) );
  AND2_X1 U569 ( .A1(n692), .A2(n521), .ZN(n707) );
  NOR2_X1 U570 ( .A1(G1384), .A2(n608), .ZN(n609) );
  BUF_X1 U571 ( .A(n555), .Z(n877) );
  NOR2_X1 U572 ( .A1(n534), .A2(n533), .ZN(n608) );
  BUF_X1 U573 ( .A(n608), .Z(G164) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U575 ( .A1(G114), .A2(n882), .ZN(n523) );
  XNOR2_X1 U576 ( .A(n523), .B(KEYINPUT92), .ZN(n526) );
  AND2_X1 U577 ( .A1(n528), .A2(G2105), .ZN(n881) );
  NAND2_X1 U578 ( .A1(G126), .A2(n881), .ZN(n524) );
  XOR2_X1 U579 ( .A(KEYINPUT91), .B(n524), .Z(n525) );
  NAND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n534) );
  NOR2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XOR2_X1 U582 ( .A(KEYINPUT17), .B(n527), .Z(n551) );
  NAND2_X1 U583 ( .A1(G138), .A2(n551), .ZN(n530) );
  INV_X1 U584 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U585 ( .A1(G2105), .A2(n528), .ZN(n555) );
  NAND2_X1 U586 ( .A1(G102), .A2(n877), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U588 ( .A(KEYINPUT93), .ZN(n531) );
  XNOR2_X1 U589 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .ZN(n535) );
  XOR2_X1 U591 ( .A(n535), .B(KEYINPUT66), .Z(n598) );
  NAND2_X1 U592 ( .A1(n791), .A2(G51), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n536), .B(KEYINPUT80), .ZN(n539) );
  INV_X1 U594 ( .A(G651), .ZN(n542) );
  NOR2_X1 U595 ( .A1(G543), .A2(n542), .ZN(n537) );
  XOR2_X2 U596 ( .A(KEYINPUT1), .B(n537), .Z(n790) );
  NAND2_X1 U597 ( .A1(G63), .A2(n790), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U599 ( .A(KEYINPUT6), .B(n540), .ZN(n549) );
  NOR2_X1 U600 ( .A1(G543), .A2(G651), .ZN(n794) );
  NAND2_X1 U601 ( .A1(n794), .A2(G89), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n541), .B(KEYINPUT4), .ZN(n545) );
  OR2_X1 U603 ( .A1(n598), .A2(n542), .ZN(n543) );
  XNOR2_X2 U604 ( .A(KEYINPUT67), .B(n543), .ZN(n795) );
  NAND2_X1 U605 ( .A1(G76), .A2(n795), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(KEYINPUT79), .B(n546), .ZN(n547) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n547), .ZN(n548) );
  NOR2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(n550), .Z(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(n882), .A2(G113), .ZN(n554) );
  INV_X1 U613 ( .A(n551), .ZN(n552) );
  INV_X2 U614 ( .A(n552), .ZN(n878) );
  NAND2_X1 U615 ( .A1(n878), .A2(G137), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n562) );
  INV_X1 U617 ( .A(KEYINPUT65), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n555), .A2(G101), .ZN(n556) );
  XOR2_X1 U619 ( .A(n556), .B(KEYINPUT23), .Z(n558) );
  NAND2_X1 U620 ( .A1(n881), .A2(G125), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G91), .A2(n794), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G65), .A2(n790), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n791), .A2(G53), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT72), .B(n565), .Z(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n795), .A2(G78), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(G299) );
  NAND2_X1 U631 ( .A1(G64), .A2(n790), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G52), .A2(n791), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n572), .B(KEYINPUT69), .ZN(n578) );
  XNOR2_X1 U635 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G90), .A2(n794), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G77), .A2(n795), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n576), .B(n575), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U641 ( .A(KEYINPUT71), .B(n579), .ZN(G171) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G88), .A2(n794), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G62), .A2(n790), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G75), .A2(n795), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT87), .B(n582), .Z(n584) );
  NAND2_X1 U648 ( .A1(n791), .A2(G50), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(G166) );
  INV_X1 U651 ( .A(G166), .ZN(G303) );
  NAND2_X1 U652 ( .A1(G86), .A2(n794), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G61), .A2(n790), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n795), .A2(G73), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT2), .B(n589), .Z(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n791), .A2(G48), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(G305) );
  NAND2_X1 U660 ( .A1(G49), .A2(n791), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G74), .A2(G651), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U663 ( .A1(n790), .A2(n596), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n597), .B(KEYINPUT86), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G87), .A2(n598), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n600), .A2(n599), .ZN(G288) );
  NAND2_X1 U667 ( .A1(n795), .A2(G72), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n794), .A2(G85), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U670 ( .A(KEYINPUT68), .B(n603), .Z(n607) );
  NAND2_X1 U671 ( .A1(G60), .A2(n790), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G47), .A2(n791), .ZN(n604) );
  AND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n607), .A2(n606), .ZN(G290) );
  INV_X1 U675 ( .A(G299), .ZN(n952) );
  XNOR2_X1 U676 ( .A(n609), .B(KEYINPUT64), .ZN(n708) );
  NAND2_X1 U677 ( .A1(G160), .A2(G40), .ZN(n709) );
  XOR2_X1 U678 ( .A(n709), .B(KEYINPUT100), .Z(n610) );
  NAND2_X2 U679 ( .A1(n708), .A2(n610), .ZN(n670) );
  NAND2_X1 U680 ( .A1(n651), .A2(G2072), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n611), .B(KEYINPUT27), .ZN(n613) );
  XNOR2_X1 U682 ( .A(G1956), .B(KEYINPUT101), .ZN(n979) );
  NOR2_X1 U683 ( .A1(n979), .A2(n651), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n645) );
  NOR2_X1 U685 ( .A1(n952), .A2(n645), .ZN(n614) );
  XOR2_X1 U686 ( .A(n614), .B(KEYINPUT28), .Z(n649) );
  XOR2_X1 U687 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n616) );
  NAND2_X1 U688 ( .A1(G56), .A2(n790), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n794), .A2(G81), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT12), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G68), .A2(n795), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U694 ( .A(KEYINPUT13), .B(n620), .Z(n621) );
  NOR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n791), .A2(G43), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n962) );
  INV_X1 U698 ( .A(G1996), .ZN(n923) );
  NOR2_X1 U699 ( .A1(n670), .A2(n923), .ZN(n625) );
  XOR2_X1 U700 ( .A(n625), .B(KEYINPUT26), .Z(n627) );
  NAND2_X1 U701 ( .A1(n670), .A2(G1341), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n962), .A2(n628), .ZN(n641) );
  NAND2_X1 U704 ( .A1(G92), .A2(n794), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G79), .A2(n795), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n790), .A2(G66), .ZN(n631) );
  XOR2_X1 U708 ( .A(KEYINPUT76), .B(n631), .Z(n632) );
  INV_X1 U709 ( .A(n633), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT15), .ZN(n637) );
  XNOR2_X2 U711 ( .A(KEYINPUT77), .B(n637), .ZN(n949) );
  NAND2_X1 U712 ( .A1(G1348), .A2(n670), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G2067), .A2(n651), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n949), .A2(n642), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n949), .A2(n642), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n952), .A2(n645), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n651), .A2(G1961), .ZN(n653) );
  XOR2_X1 U721 ( .A(G2078), .B(KEYINPUT25), .Z(n924) );
  NOR2_X1 U722 ( .A1(n670), .A2(n924), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n662) );
  OR2_X1 U724 ( .A1(n662), .A2(G301), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n667) );
  NOR2_X1 U726 ( .A1(G1966), .A2(n701), .ZN(n681) );
  NOR2_X1 U727 ( .A1(G2084), .A2(n670), .ZN(n678) );
  INV_X1 U728 ( .A(n678), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n656), .A2(G8), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT30), .B(n658), .ZN(n659) );
  NOR2_X1 U731 ( .A1(G168), .A2(n659), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n662), .A2(G301), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT31), .B(n665), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n679) );
  NAND2_X1 U737 ( .A1(n679), .A2(G286), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n675) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n701), .ZN(n672) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n670), .ZN(n671) );
  NOR2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U742 ( .A1(G303), .A2(n673), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n676), .A2(G8), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(KEYINPUT32), .ZN(n685) );
  NAND2_X1 U746 ( .A1(G8), .A2(n678), .ZN(n683) );
  INV_X1 U747 ( .A(n679), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(KEYINPUT104), .ZN(n696) );
  NOR2_X1 U752 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U753 ( .A1(G8), .A2(n687), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n696), .A2(n688), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n689), .A2(n701), .ZN(n692) );
  NOR2_X1 U756 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U757 ( .A(n690), .B(KEYINPUT24), .Z(n691) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n699) );
  NOR2_X1 U759 ( .A1(G1971), .A2(G303), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n699), .A2(n693), .ZN(n953) );
  INV_X1 U761 ( .A(KEYINPUT33), .ZN(n694) );
  AND2_X1 U762 ( .A1(n953), .A2(n694), .ZN(n695) );
  AND2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  INV_X1 U764 ( .A(n697), .ZN(n705) );
  XOR2_X1 U765 ( .A(G1981), .B(G305), .Z(n944) );
  NAND2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n948) );
  INV_X1 U767 ( .A(n948), .ZN(n698) );
  OR2_X1 U768 ( .A1(KEYINPUT33), .A2(n520), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n699), .A2(KEYINPUT33), .ZN(n700) );
  OR2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n702) );
  AND2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n519), .ZN(n706) );
  XNOR2_X1 U773 ( .A(n522), .B(KEYINPUT105), .ZN(n745) );
  XNOR2_X1 U774 ( .A(G1986), .B(G290), .ZN(n960) );
  NOR2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n756) );
  NAND2_X1 U776 ( .A1(n960), .A2(n756), .ZN(n743) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n754) );
  XNOR2_X1 U778 ( .A(KEYINPUT95), .B(KEYINPUT36), .ZN(n720) );
  NAND2_X1 U779 ( .A1(G128), .A2(n881), .ZN(n711) );
  NAND2_X1 U780 ( .A1(G116), .A2(n882), .ZN(n710) );
  NAND2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U782 ( .A(KEYINPUT35), .B(n712), .ZN(n718) );
  NAND2_X1 U783 ( .A1(G104), .A2(n877), .ZN(n714) );
  NAND2_X1 U784 ( .A1(G140), .A2(n878), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U786 ( .A(KEYINPUT94), .B(KEYINPUT34), .Z(n715) );
  XNOR2_X1 U787 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U789 ( .A(n720), .B(n719), .ZN(n894) );
  NOR2_X1 U790 ( .A1(n754), .A2(n894), .ZN(n1007) );
  NAND2_X1 U791 ( .A1(n756), .A2(n1007), .ZN(n752) );
  INV_X1 U792 ( .A(n752), .ZN(n741) );
  NAND2_X1 U793 ( .A1(G129), .A2(n881), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G117), .A2(n882), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U796 ( .A1(n877), .A2(G105), .ZN(n723) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(n723), .Z(n724) );
  NOR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U799 ( .A(KEYINPUT97), .B(n726), .Z(n728) );
  NAND2_X1 U800 ( .A1(n878), .A2(G141), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U802 ( .A(KEYINPUT98), .B(n729), .ZN(n896) );
  NAND2_X1 U803 ( .A1(n896), .A2(G1996), .ZN(n738) );
  NAND2_X1 U804 ( .A1(G119), .A2(n881), .ZN(n731) );
  NAND2_X1 U805 ( .A1(G107), .A2(n882), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U807 ( .A(KEYINPUT96), .B(n732), .Z(n736) );
  NAND2_X1 U808 ( .A1(n877), .A2(G95), .ZN(n734) );
  NAND2_X1 U809 ( .A1(G131), .A2(n878), .ZN(n733) );
  AND2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n889) );
  NAND2_X1 U812 ( .A1(G1991), .A2(n889), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U814 ( .A(n739), .B(KEYINPUT99), .ZN(n1020) );
  INV_X1 U815 ( .A(n756), .ZN(n740) );
  NOR2_X1 U816 ( .A1(n1020), .A2(n740), .ZN(n748) );
  NOR2_X1 U817 ( .A1(n741), .A2(n748), .ZN(n742) );
  AND2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n759) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n896), .ZN(n1015) );
  NOR2_X1 U821 ( .A1(G1991), .A2(n889), .ZN(n1003) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n746) );
  NOR2_X1 U823 ( .A1(n1003), .A2(n746), .ZN(n747) );
  NOR2_X1 U824 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U825 ( .A(n749), .B(KEYINPUT106), .ZN(n750) );
  NOR2_X1 U826 ( .A1(n1015), .A2(n750), .ZN(n751) );
  XNOR2_X1 U827 ( .A(n751), .B(KEYINPUT39), .ZN(n753) );
  NAND2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n754), .A2(n894), .ZN(n1008) );
  NAND2_X1 U830 ( .A1(n755), .A2(n1008), .ZN(n757) );
  NAND2_X1 U831 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U833 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U835 ( .A(G57), .ZN(G237) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U838 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U839 ( .A(G223), .ZN(n826) );
  NAND2_X1 U840 ( .A1(n826), .A2(G567), .ZN(n762) );
  XOR2_X1 U841 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U842 ( .A(G860), .ZN(n789) );
  OR2_X1 U843 ( .A1(n962), .A2(n789), .ZN(G153) );
  INV_X1 U844 ( .A(G868), .ZN(n767) );
  NOR2_X1 U845 ( .A1(n767), .A2(G171), .ZN(n763) );
  XNOR2_X1 U846 ( .A(n763), .B(KEYINPUT75), .ZN(n765) );
  NAND2_X1 U847 ( .A1(n767), .A2(n949), .ZN(n764) );
  NAND2_X1 U848 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U849 ( .A(KEYINPUT78), .B(n766), .ZN(G284) );
  NOR2_X1 U850 ( .A1(G286), .A2(n767), .ZN(n769) );
  NOR2_X1 U851 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U852 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U853 ( .A1(n789), .A2(G559), .ZN(n770) );
  INV_X1 U854 ( .A(n949), .ZN(n899) );
  NAND2_X1 U855 ( .A1(n770), .A2(n899), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(G868), .A2(n962), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G868), .A2(n899), .ZN(n772) );
  NOR2_X1 U859 ( .A1(G559), .A2(n772), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(G282) );
  XOR2_X1 U861 ( .A(G2100), .B(KEYINPUT84), .Z(n786) );
  NAND2_X1 U862 ( .A1(G123), .A2(n881), .ZN(n775) );
  XOR2_X1 U863 ( .A(KEYINPUT18), .B(n775), .Z(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT81), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G135), .A2(n878), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT82), .B(n779), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G99), .A2(n877), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G111), .A2(n882), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U872 ( .A(KEYINPUT83), .B(n784), .Z(n1002) );
  XNOR2_X1 U873 ( .A(G2096), .B(n1002), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(G156) );
  XNOR2_X1 U875 ( .A(n962), .B(KEYINPUT85), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n899), .A2(G559), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n788), .B(n787), .ZN(n806) );
  NAND2_X1 U878 ( .A1(n789), .A2(n806), .ZN(n800) );
  NAND2_X1 U879 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U880 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G93), .A2(n794), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G80), .A2(n795), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n809) );
  XOR2_X1 U886 ( .A(n800), .B(n809), .Z(G145) );
  XNOR2_X1 U887 ( .A(n809), .B(KEYINPUT19), .ZN(n805) );
  XNOR2_X1 U888 ( .A(n952), .B(G288), .ZN(n803) );
  XNOR2_X1 U889 ( .A(G290), .B(G303), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n801), .B(G305), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n805), .B(n804), .ZN(n898) );
  XNOR2_X1 U893 ( .A(n898), .B(n806), .ZN(n807) );
  NAND2_X1 U894 ( .A1(n807), .A2(G868), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(KEYINPUT88), .ZN(n811) );
  OR2_X1 U896 ( .A1(G868), .A2(n809), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U900 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U901 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U902 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U903 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U905 ( .A1(G661), .A2(G483), .ZN(n824) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n816) );
  XNOR2_X1 U907 ( .A(KEYINPUT22), .B(n816), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n817), .A2(G96), .ZN(n818) );
  NOR2_X1 U909 ( .A1(n818), .A2(G218), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT89), .ZN(n831) );
  NAND2_X1 U911 ( .A1(n831), .A2(G2106), .ZN(n823) );
  NAND2_X1 U912 ( .A1(G69), .A2(G120), .ZN(n820) );
  NOR2_X1 U913 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U914 ( .A1(G108), .A2(n821), .ZN(n832) );
  NAND2_X1 U915 ( .A1(n832), .A2(G567), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n853) );
  NOR2_X1 U917 ( .A1(n824), .A2(n853), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n825), .B(KEYINPUT90), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G36), .A2(n829), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U922 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n828) );
  XOR2_X1 U924 ( .A(KEYINPUT109), .B(n828), .Z(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U932 ( .A(G1981), .B(KEYINPUT112), .ZN(n842) );
  XOR2_X1 U933 ( .A(G1976), .B(G1971), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1966), .B(G1956), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U936 ( .A(G1961), .B(G1986), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2474), .B(KEYINPUT41), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2678), .B(KEYINPUT111), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U946 ( .A(KEYINPUT110), .B(G2072), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2100), .B(G2096), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U952 ( .A(G2078), .B(G2084), .Z(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G227) );
  INV_X1 U954 ( .A(n853), .ZN(G319) );
  NAND2_X1 U955 ( .A1(G124), .A2(n881), .ZN(n854) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(n854), .Z(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G100), .A2(n877), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G136), .A2(n878), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G112), .A2(n882), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U963 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G106), .A2(n877), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G142), .A2(n878), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT45), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G130), .A2(n881), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n882), .A2(G118), .ZN(n867) );
  XOR2_X1 U971 ( .A(KEYINPUT114), .B(n867), .Z(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n876) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT117), .B(KEYINPUT115), .ZN(n870) );
  XNOR2_X1 U975 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U976 ( .A(n872), .B(n1002), .Z(n874) );
  XNOR2_X1 U977 ( .A(G164), .B(G162), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G127), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(KEYINPUT116), .B(n885), .Z(n886) );
  XNOR2_X1 U987 ( .A(KEYINPUT47), .B(n886), .ZN(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n1010) );
  XNOR2_X1 U989 ( .A(n889), .B(n1010), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U991 ( .A(G160), .B(n892), .Z(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U993 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U995 ( .A(G286), .B(n898), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n962), .B(n899), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(G171), .B(n902), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n918) );
  XNOR2_X1 U1003 ( .A(G2451), .B(G2443), .ZN(n915) );
  XOR2_X1 U1004 ( .A(G2446), .B(G2454), .Z(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT107), .B(G2435), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1007 ( .A(KEYINPUT108), .B(G2438), .Z(n909) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1010 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G2430), .B(G2427), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n916), .A2(G14), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n921), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  INV_X1 U1021 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(G2084), .B(G34), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(n922), .B(KEYINPUT54), .ZN(n941) );
  XOR2_X1 U1024 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n936) );
  XNOR2_X1 U1025 ( .A(G1991), .B(G25), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(G32), .B(n923), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G2067), .B(G26), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(G27), .B(n924), .ZN(n925) );
  NOR2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(KEYINPUT119), .B(n931), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n934), .A2(G28), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n936), .B(n935), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(n939), .B(KEYINPUT121), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(n942), .Z(n943) );
  NOR2_X1 U1042 ( .A1(G29), .A2(n943), .ZN(n999) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .ZN(n968) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G168), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(n946), .B(KEYINPUT57), .ZN(n966) );
  NAND2_X1 U1047 ( .A1(G1971), .A2(G303), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G1348), .B(n949), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n952), .B(G1956), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(G1961), .B(G301), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT122), .B(n961), .Z(n964) );
  XNOR2_X1 U1058 ( .A(G1341), .B(n962), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n996) );
  INV_X1 U1062 ( .A(G16), .ZN(n994) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G1976), .B(G23), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1066 ( .A(KEYINPUT124), .B(n971), .Z(n973) );
  XNOR2_X1 U1067 ( .A(G1986), .B(G24), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT58), .B(n974), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G21), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G5), .B(G1961), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n990) );
  XOR2_X1 U1074 ( .A(n979), .B(G20), .Z(n984) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(G1981), .B(G6), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(n982), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT59), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(n985), .B(G4), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n988), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1085 ( .A(n991), .B(KEYINPUT125), .Z(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n992), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(KEYINPUT126), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(G11), .A2(n1000), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT127), .ZN(n1028) );
  XNOR2_X1 U1093 ( .A(G160), .B(G2084), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1022) );
  XOR2_X1 U1098 ( .A(G2072), .B(n1010), .Z(n1012) );
  XOR2_X1 U1099 ( .A(G164), .B(G2078), .Z(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT50), .B(n1013), .Z(n1018) );
  XOR2_X1 U1102 ( .A(G2090), .B(G162), .Z(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT51), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1023), .ZN(n1025) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(G29), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

