

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754;

  XNOR2_X1 U372 ( .A(n599), .B(n598), .ZN(n391) );
  XNOR2_X1 U373 ( .A(n471), .B(n470), .ZN(n669) );
  INV_X1 U374 ( .A(G953), .ZN(n742) );
  XNOR2_X1 U375 ( .A(KEYINPUT70), .B(KEYINPUT0), .ZN(n349) );
  NAND2_X1 U376 ( .A1(n545), .A2(n365), .ZN(n350) );
  XNOR2_X2 U377 ( .A(KEYINPUT38), .B(n622), .ZN(n682) );
  NOR2_X1 U378 ( .A1(n420), .A2(n418), .ZN(n417) );
  XNOR2_X1 U379 ( .A(n465), .B(n372), .ZN(n374) );
  NAND2_X1 U380 ( .A1(n569), .A2(n441), .ZN(n401) );
  NOR2_X1 U381 ( .A1(n587), .A2(n650), .ZN(n426) );
  NOR2_X1 U382 ( .A1(n583), .A2(n593), .ZN(n600) );
  XNOR2_X1 U383 ( .A(n492), .B(n491), .ZN(n604) );
  AND2_X1 U384 ( .A1(n684), .A2(n442), .ZN(n441) );
  XNOR2_X1 U385 ( .A(n405), .B(KEYINPUT4), .ZN(n478) );
  INV_X2 U386 ( .A(KEYINPUT80), .ZN(n413) );
  INV_X2 U387 ( .A(KEYINPUT71), .ZN(n410) );
  XNOR2_X2 U388 ( .A(n351), .B(n472), .ZN(n584) );
  NAND2_X2 U389 ( .A1(n489), .A2(n499), .ZN(n351) );
  XNOR2_X2 U390 ( .A(n352), .B(n485), .ZN(n489) );
  NAND2_X1 U391 ( .A1(n356), .A2(n355), .ZN(n352) );
  AND2_X1 U392 ( .A1(n569), .A2(n564), .ZN(n565) );
  XNOR2_X2 U393 ( .A(n429), .B(n349), .ZN(n569) );
  NAND2_X1 U394 ( .A1(n478), .A2(n724), .ZN(n355) );
  NAND2_X1 U395 ( .A1(n353), .A2(n354), .ZN(n356) );
  INV_X1 U396 ( .A(n478), .ZN(n353) );
  INV_X1 U397 ( .A(n724), .ZN(n354) );
  XNOR2_X2 U398 ( .A(n407), .B(n723), .ZN(n405) );
  XNOR2_X2 U399 ( .A(n410), .B(G101), .ZN(n548) );
  AND2_X1 U400 ( .A1(n400), .A2(n439), .ZN(n399) );
  NAND2_X1 U401 ( .A1(n398), .A2(n397), .ZN(n400) );
  XNOR2_X1 U402 ( .A(n503), .B(n502), .ZN(n533) );
  XNOR2_X1 U403 ( .A(G140), .B(KEYINPUT10), .ZN(n502) );
  NAND2_X1 U404 ( .A1(n448), .A2(n447), .ZN(n666) );
  AND2_X1 U405 ( .A1(n451), .A2(n449), .ZN(n448) );
  NAND2_X1 U406 ( .A1(n453), .A2(n458), .ZN(n447) );
  INV_X1 U407 ( .A(n666), .ZN(n561) );
  XNOR2_X1 U408 ( .A(n543), .B(n544), .ZN(n470) );
  OR2_X1 U409 ( .A1(n721), .A2(G902), .ZN(n471) );
  OR2_X1 U410 ( .A1(n656), .A2(n639), .ZN(n398) );
  NAND2_X1 U411 ( .A1(n387), .A2(KEYINPUT48), .ZN(n386) );
  XNOR2_X1 U412 ( .A(n419), .B(KEYINPUT79), .ZN(n418) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n507) );
  XNOR2_X1 U414 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n504) );
  XNOR2_X1 U415 ( .A(n506), .B(n422), .ZN(n421) );
  INV_X1 U416 ( .A(KEYINPUT11), .ZN(n422) );
  XNOR2_X1 U417 ( .A(G113), .B(G131), .ZN(n506) );
  XOR2_X1 U418 ( .A(n580), .B(KEYINPUT6), .Z(n611) );
  NAND2_X1 U419 ( .A1(n581), .A2(n681), .ZN(n396) );
  NOR2_X1 U420 ( .A1(n670), .A2(n669), .ZN(n564) );
  XNOR2_X1 U421 ( .A(n467), .B(n568), .ZN(n694) );
  INV_X1 U422 ( .A(KEYINPUT33), .ZN(n568) );
  NOR2_X1 U423 ( .A1(n567), .A2(n611), .ZN(n467) );
  XNOR2_X1 U424 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U425 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n585) );
  NAND2_X1 U426 ( .A1(n694), .A2(n569), .ZN(n446) );
  INV_X1 U427 ( .A(KEYINPUT34), .ZN(n445) );
  NAND2_X1 U428 ( .A1(n545), .A2(n364), .ZN(n406) );
  NAND2_X1 U429 ( .A1(n580), .A2(n669), .ZN(n464) );
  NAND2_X1 U430 ( .A1(n430), .A2(n350), .ZN(n439) );
  AND2_X1 U431 ( .A1(n431), .A2(n363), .ZN(n430) );
  AND2_X1 U432 ( .A1(n406), .A2(n403), .ZN(n402) );
  INV_X1 U433 ( .A(KEYINPUT44), .ZN(n403) );
  XNOR2_X1 U434 ( .A(n443), .B(G128), .ZN(n515) );
  INV_X1 U435 ( .A(G143), .ZN(n443) );
  NAND2_X1 U436 ( .A1(G469), .A2(n457), .ZN(n456) );
  INV_X1 U437 ( .A(G902), .ZN(n457) );
  NAND2_X1 U438 ( .A1(n461), .A2(G902), .ZN(n459) );
  NOR2_X1 U439 ( .A1(n384), .A2(n383), .ZN(n624) );
  INV_X1 U440 ( .A(n661), .ZN(n390) );
  XNOR2_X1 U441 ( .A(n527), .B(n528), .ZN(n738) );
  XNOR2_X1 U442 ( .A(G131), .B(KEYINPUT4), .ZN(n528) );
  NOR2_X1 U443 ( .A1(n573), .A2(n437), .ZN(n433) );
  XOR2_X1 U444 ( .A(G137), .B(KEYINPUT73), .Z(n534) );
  XNOR2_X1 U445 ( .A(n515), .B(G134), .ZN(n527) );
  XNOR2_X1 U446 ( .A(n548), .B(n408), .ZN(n407) );
  XNOR2_X1 U447 ( .A(n409), .B(KEYINPUT77), .ZN(n408) );
  INV_X1 U448 ( .A(KEYINPUT78), .ZN(n409) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n493) );
  OR2_X1 U450 ( .A1(n456), .A2(n454), .ZN(n450) );
  AND2_X1 U451 ( .A1(n455), .A2(n454), .ZN(n453) );
  XNOR2_X1 U452 ( .A(n594), .B(n428), .ZN(n680) );
  INV_X1 U453 ( .A(KEYINPUT110), .ZN(n428) );
  INV_X1 U454 ( .A(n670), .ZN(n442) );
  XNOR2_X1 U455 ( .A(G119), .B(G110), .ZN(n535) );
  XOR2_X1 U456 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n521) );
  XNOR2_X1 U457 ( .A(n512), .B(n511), .ZN(n714) );
  XNOR2_X1 U458 ( .A(n510), .B(n473), .ZN(n511) );
  XNOR2_X1 U459 ( .A(n505), .B(n421), .ZN(n512) );
  NAND2_X1 U460 ( .A1(n395), .A2(n393), .ZN(n583) );
  XNOR2_X1 U461 ( .A(n396), .B(n582), .ZN(n395) );
  XNOR2_X1 U462 ( .A(KEYINPUT19), .B(KEYINPUT69), .ZN(n491) );
  NOR2_X1 U463 ( .A1(n561), .A2(n669), .ZN(n440) );
  NAND2_X1 U464 ( .A1(n557), .A2(KEYINPUT88), .ZN(n432) );
  XNOR2_X1 U465 ( .A(n597), .B(n368), .ZN(n751) );
  XNOR2_X1 U466 ( .A(n469), .B(KEYINPUT35), .ZN(n749) );
  XNOR2_X1 U467 ( .A(n446), .B(n445), .ZN(n444) );
  XNOR2_X1 U468 ( .A(n563), .B(n562), .ZN(n656) );
  NOR2_X1 U469 ( .A1(n566), .A2(n593), .ZN(n639) );
  XNOR2_X1 U470 ( .A(n632), .B(KEYINPUT92), .ZN(n633) );
  XNOR2_X1 U471 ( .A(n717), .B(n718), .ZN(n375) );
  INV_X1 U472 ( .A(KEYINPUT56), .ZN(n378) );
  INV_X1 U473 ( .A(G119), .ZN(n414) );
  INV_X1 U474 ( .A(n406), .ZN(n644) );
  INV_X1 U475 ( .A(n439), .ZN(n637) );
  INV_X1 U476 ( .A(n669), .ZN(n394) );
  INV_X1 U477 ( .A(n545), .ZN(n558) );
  INV_X1 U478 ( .A(n679), .ZN(n397) );
  XNOR2_X1 U479 ( .A(n603), .B(KEYINPUT83), .ZN(n357) );
  XOR2_X2 U480 ( .A(KEYINPUT75), .B(KEYINPUT3), .Z(n358) );
  OR2_X1 U481 ( .A1(n617), .A2(n394), .ZN(n359) );
  AND2_X1 U482 ( .A1(n402), .A2(n374), .ZN(n360) );
  INV_X1 U483 ( .A(G469), .ZN(n461) );
  AND2_X1 U484 ( .A1(n547), .A2(G210), .ZN(n361) );
  AND2_X1 U485 ( .A1(n662), .A2(n625), .ZN(n362) );
  AND2_X1 U486 ( .A1(n432), .A2(n440), .ZN(n363) );
  NOR2_X1 U487 ( .A1(n561), .A2(n464), .ZN(n364) );
  NOR2_X1 U488 ( .A1(n557), .A2(KEYINPUT88), .ZN(n365) );
  XNOR2_X1 U489 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n366) );
  XOR2_X1 U490 ( .A(n488), .B(n487), .Z(n367) );
  INV_X1 U491 ( .A(KEYINPUT1), .ZN(n454) );
  XNOR2_X1 U492 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n368) );
  XOR2_X1 U493 ( .A(n709), .B(n708), .Z(n369) );
  INV_X1 U494 ( .A(KEYINPUT48), .ZN(n618) );
  XOR2_X1 U495 ( .A(n714), .B(n713), .Z(n370) );
  XOR2_X1 U496 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n371) );
  XNOR2_X1 U497 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n372) );
  NOR2_X1 U498 ( .A1(G952), .A2(n742), .ZN(n722) );
  INV_X1 U499 ( .A(n722), .ZN(n380) );
  XNOR2_X1 U500 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n373) );
  NAND2_X1 U501 ( .A1(n374), .A2(n406), .ZN(n404) );
  XNOR2_X1 U502 ( .A(n374), .B(n414), .ZN(n750) );
  XNOR2_X1 U503 ( .A(n720), .B(n721), .ZN(n376) );
  XNOR2_X1 U504 ( .A(n710), .B(n369), .ZN(n711) );
  XNOR2_X1 U505 ( .A(n415), .B(n371), .ZN(n732) );
  NOR2_X1 U506 ( .A1(n375), .A2(n722), .ZN(G63) );
  NAND2_X1 U507 ( .A1(n433), .A2(n434), .ZN(n416) );
  XNOR2_X1 U508 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X1 U509 ( .A1(n376), .A2(n722), .ZN(G66) );
  NAND2_X1 U510 ( .A1(n399), .A2(n572), .ZN(n573) );
  NAND2_X1 U511 ( .A1(n444), .A2(n357), .ZN(n469) );
  XNOR2_X1 U512 ( .A(n377), .B(n373), .ZN(G60) );
  NAND2_X1 U513 ( .A1(n382), .A2(n380), .ZN(n377) );
  XNOR2_X1 U514 ( .A(n379), .B(n378), .ZN(G51) );
  NAND2_X1 U515 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U516 ( .A(n630), .B(n367), .ZN(n381) );
  XNOR2_X1 U517 ( .A(n715), .B(n370), .ZN(n382) );
  XNOR2_X1 U518 ( .A(n556), .B(KEYINPUT65), .ZN(n438) );
  NAND2_X1 U519 ( .A1(n389), .A2(n390), .ZN(n383) );
  NAND2_X1 U520 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U521 ( .A1(n388), .A2(n391), .ZN(n385) );
  INV_X1 U522 ( .A(n391), .ZN(n387) );
  AND2_X1 U523 ( .A1(n392), .A2(n618), .ZN(n388) );
  OR2_X1 U524 ( .A1(n392), .A2(n618), .ZN(n389) );
  AND2_X1 U525 ( .A1(n609), .A2(n427), .ZN(n392) );
  AND2_X1 U526 ( .A1(n589), .A2(n394), .ZN(n393) );
  XNOR2_X2 U527 ( .A(n401), .B(n366), .ZN(n545) );
  NAND2_X1 U528 ( .A1(n404), .A2(KEYINPUT44), .ZN(n556) );
  XNOR2_X1 U529 ( .A(n405), .B(n531), .ZN(n532) );
  XNOR2_X2 U530 ( .A(n412), .B(n411), .ZN(n723) );
  XNOR2_X2 U531 ( .A(G104), .B(G107), .ZN(n411) );
  XNOR2_X2 U532 ( .A(n413), .B(G110), .ZN(n412) );
  NAND2_X1 U533 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U534 ( .A1(n360), .A2(n468), .ZN(n419) );
  NAND2_X1 U535 ( .A1(n436), .A2(n435), .ZN(n420) );
  XNOR2_X1 U536 ( .A(n423), .B(n615), .ZN(n616) );
  AND2_X1 U537 ( .A1(n584), .A2(n619), .ZN(n423) );
  INV_X1 U538 ( .A(n658), .ZN(n427) );
  INV_X1 U539 ( .A(KEYINPUT89), .ZN(n437) );
  XNOR2_X2 U540 ( .A(G119), .B(G116), .ZN(n475) );
  XNOR2_X1 U541 ( .A(n424), .B(n552), .ZN(n631) );
  XNOR2_X1 U542 ( .A(n551), .B(n474), .ZN(n424) );
  XNOR2_X2 U543 ( .A(n425), .B(n476), .ZN(n546) );
  XNOR2_X2 U544 ( .A(n358), .B(n475), .ZN(n425) );
  NAND2_X1 U545 ( .A1(n600), .A2(n682), .ZN(n586) );
  NAND2_X1 U546 ( .A1(n624), .A2(n662), .ZN(n741) );
  XNOR2_X1 U547 ( .A(n426), .B(n588), .ZN(n753) );
  XNOR2_X2 U548 ( .A(n546), .B(n477), .ZN(n724) );
  XNOR2_X1 U549 ( .A(n546), .B(n361), .ZN(n551) );
  NAND2_X1 U550 ( .A1(n545), .A2(n466), .ZN(n465) );
  NAND2_X1 U551 ( .A1(n753), .A2(n751), .ZN(n599) );
  NAND2_X1 U552 ( .A1(n680), .A2(n684), .ZN(n595) );
  NOR2_X2 U553 ( .A1(n604), .A2(n498), .ZN(n429) );
  NAND2_X1 U554 ( .A1(n558), .A2(KEYINPUT88), .ZN(n431) );
  INV_X1 U555 ( .A(n438), .ZN(n434) );
  NAND2_X1 U556 ( .A1(n573), .A2(n437), .ZN(n435) );
  NAND2_X1 U557 ( .A1(n438), .A2(n437), .ZN(n436) );
  OR2_X1 U558 ( .A1(n707), .A2(n456), .ZN(n455) );
  INV_X1 U559 ( .A(n452), .ZN(n458) );
  OR2_X1 U560 ( .A1(n707), .A2(n450), .ZN(n449) );
  NAND2_X1 U561 ( .A1(n452), .A2(KEYINPUT1), .ZN(n451) );
  NAND2_X1 U562 ( .A1(n460), .A2(n459), .ZN(n452) );
  NAND2_X1 U563 ( .A1(n458), .A2(n455), .ZN(n593) );
  NAND2_X1 U564 ( .A1(n707), .A2(n461), .ZN(n460) );
  NAND2_X1 U565 ( .A1(n462), .A2(n627), .ZN(n629) );
  OR2_X2 U566 ( .A1(n732), .A2(n463), .ZN(n462) );
  NAND2_X1 U567 ( .A1(n624), .A2(n362), .ZN(n463) );
  NOR2_X1 U568 ( .A1(n732), .A2(n741), .ZN(n663) );
  NOR2_X1 U569 ( .A1(n555), .A2(n359), .ZN(n466) );
  NAND2_X1 U570 ( .A1(n564), .A2(n561), .ZN(n567) );
  INV_X1 U571 ( .A(n749), .ZN(n468) );
  BUF_X1 U572 ( .A(n663), .Z(n699) );
  XNOR2_X1 U573 ( .A(n533), .B(n504), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n541), .B(n540), .ZN(n721) );
  AND2_X1 U575 ( .A1(G210), .A2(n490), .ZN(n472) );
  XOR2_X1 U576 ( .A(n509), .B(n508), .Z(n473) );
  XOR2_X1 U577 ( .A(n550), .B(n549), .Z(n474) );
  NOR2_X1 U578 ( .A1(n571), .A2(n570), .ZN(n684) );
  NAND2_X1 U579 ( .A1(n635), .A2(n380), .ZN(n636) );
  XNOR2_X1 U580 ( .A(n636), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U581 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n488) );
  XNOR2_X1 U582 ( .A(KEYINPUT16), .B(G122), .ZN(n477) );
  XOR2_X1 U583 ( .A(G113), .B(KEYINPUT76), .Z(n476) );
  XOR2_X2 U584 ( .A(G146), .B(G125), .Z(n503) );
  XOR2_X1 U585 ( .A(n515), .B(n503), .Z(n480) );
  NAND2_X1 U586 ( .A1(G224), .A2(n742), .ZN(n479) );
  XNOR2_X1 U587 ( .A(n480), .B(n479), .ZN(n484) );
  XOR2_X1 U588 ( .A(KEYINPUT94), .B(KEYINPUT18), .Z(n482) );
  XNOR2_X1 U589 ( .A(KEYINPUT17), .B(KEYINPUT82), .ZN(n481) );
  XNOR2_X1 U590 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U591 ( .A(n484), .B(n483), .Z(n485) );
  BUF_X1 U592 ( .A(n489), .Z(n486) );
  XNOR2_X1 U593 ( .A(n486), .B(KEYINPUT91), .ZN(n487) );
  XOR2_X1 U594 ( .A(KEYINPUT15), .B(G902), .Z(n625) );
  INV_X1 U595 ( .A(n625), .ZN(n499) );
  OR2_X1 U596 ( .A1(G237), .A2(G902), .ZN(n490) );
  NAND2_X1 U597 ( .A1(G214), .A2(n490), .ZN(n681) );
  NAND2_X1 U598 ( .A1(n584), .A2(n681), .ZN(n492) );
  XNOR2_X1 U599 ( .A(n493), .B(KEYINPUT95), .ZN(n494) );
  XOR2_X1 U600 ( .A(KEYINPUT14), .B(n494), .Z(n495) );
  NAND2_X1 U601 ( .A1(G952), .A2(n495), .ZN(n693) );
  NOR2_X1 U602 ( .A1(G953), .A2(n693), .ZN(n578) );
  AND2_X1 U603 ( .A1(G953), .A2(n495), .ZN(n496) );
  NAND2_X1 U604 ( .A1(G902), .A2(n496), .ZN(n574) );
  NOR2_X1 U605 ( .A1(G898), .A2(n574), .ZN(n497) );
  NOR2_X1 U606 ( .A1(n578), .A2(n497), .ZN(n498) );
  NAND2_X1 U607 ( .A1(n499), .A2(G234), .ZN(n500) );
  XNOR2_X1 U608 ( .A(n500), .B(KEYINPUT20), .ZN(n542) );
  NAND2_X1 U609 ( .A1(G221), .A2(n542), .ZN(n501) );
  XNOR2_X1 U610 ( .A(KEYINPUT21), .B(n501), .ZN(n670) );
  XNOR2_X1 U611 ( .A(KEYINPUT13), .B(G475), .ZN(n514) );
  XOR2_X1 U612 ( .A(KEYINPUT81), .B(n507), .Z(n547) );
  NAND2_X1 U613 ( .A1(G214), .A2(n547), .ZN(n510) );
  XOR2_X1 U614 ( .A(KEYINPUT101), .B(G104), .Z(n509) );
  XNOR2_X1 U615 ( .A(G143), .B(G122), .ZN(n508) );
  NOR2_X1 U616 ( .A1(G902), .A2(n714), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n514), .B(n513), .ZN(n571) );
  INV_X1 U618 ( .A(n527), .ZN(n519) );
  XOR2_X1 U619 ( .A(KEYINPUT103), .B(G107), .Z(n517) );
  XNOR2_X1 U620 ( .A(G116), .B(G122), .ZN(n516) );
  XNOR2_X1 U621 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U622 ( .A(n519), .B(n518), .Z(n523) );
  NAND2_X1 U623 ( .A1(G234), .A2(n742), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n537) );
  NAND2_X1 U625 ( .A1(G217), .A2(n537), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n524) );
  XNOR2_X1 U628 ( .A(n525), .B(n524), .ZN(n716) );
  NOR2_X1 U629 ( .A1(G902), .A2(n716), .ZN(n526) );
  XOR2_X1 U630 ( .A(G478), .B(n526), .Z(n570) );
  XNOR2_X1 U631 ( .A(G146), .B(n738), .ZN(n552) );
  XOR2_X1 U632 ( .A(n534), .B(G140), .Z(n530) );
  NAND2_X1 U633 ( .A1(G227), .A2(n742), .ZN(n529) );
  XNOR2_X1 U634 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n552), .B(n532), .ZN(n707) );
  XOR2_X1 U636 ( .A(n666), .B(KEYINPUT93), .Z(n617) );
  XNOR2_X1 U637 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n544) );
  XNOR2_X1 U638 ( .A(n534), .B(n533), .ZN(n740) );
  XNOR2_X1 U639 ( .A(n535), .B(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U640 ( .A(n740), .B(n536), .ZN(n541) );
  NAND2_X1 U641 ( .A1(G221), .A2(n537), .ZN(n539) );
  XOR2_X1 U642 ( .A(G128), .B(KEYINPUT24), .Z(n538) );
  XNOR2_X1 U643 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U644 ( .A1(n542), .A2(G217), .ZN(n543) );
  XOR2_X1 U645 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n550) );
  XNOR2_X1 U646 ( .A(n548), .B(G137), .ZN(n549) );
  NOR2_X1 U647 ( .A1(G902), .A2(n631), .ZN(n554) );
  XNOR2_X1 U648 ( .A(G472), .B(KEYINPUT98), .ZN(n553) );
  XNOR2_X2 U649 ( .A(n554), .B(n553), .ZN(n580) );
  INV_X1 U650 ( .A(n611), .ZN(n557) );
  XNOR2_X1 U651 ( .A(KEYINPUT84), .B(n557), .ZN(n555) );
  XNOR2_X1 U652 ( .A(KEYINPUT102), .B(n571), .ZN(n560) );
  INV_X1 U653 ( .A(n570), .ZN(n559) );
  NAND2_X1 U654 ( .A1(n560), .A2(n559), .ZN(n650) );
  INV_X1 U655 ( .A(n650), .ZN(n653) );
  NOR2_X1 U656 ( .A1(n560), .A2(n559), .ZN(n655) );
  NOR2_X1 U657 ( .A1(n653), .A2(n655), .ZN(n679) );
  NOR2_X1 U658 ( .A1(n580), .A2(n567), .ZN(n676) );
  NAND2_X1 U659 ( .A1(n569), .A2(n676), .ZN(n563) );
  XOR2_X1 U660 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n562) );
  INV_X1 U661 ( .A(n564), .ZN(n665) );
  NAND2_X1 U662 ( .A1(n580), .A2(n565), .ZN(n566) );
  NAND2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n603) );
  NAND2_X1 U664 ( .A1(n749), .A2(KEYINPUT44), .ZN(n572) );
  XNOR2_X1 U665 ( .A(KEYINPUT104), .B(n574), .ZN(n575) );
  NOR2_X1 U666 ( .A1(G900), .A2(n575), .ZN(n576) );
  XOR2_X1 U667 ( .A(KEYINPUT105), .B(n576), .Z(n577) );
  NOR2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U669 ( .A1(n670), .A2(n579), .ZN(n589) );
  XNOR2_X1 U670 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n582) );
  INV_X1 U671 ( .A(n580), .ZN(n581) );
  INV_X1 U672 ( .A(n584), .ZN(n622) );
  INV_X1 U673 ( .A(n655), .ZN(n645) );
  NOR2_X1 U674 ( .A1(n587), .A2(n645), .ZN(n661) );
  XNOR2_X1 U675 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n588) );
  XNOR2_X1 U676 ( .A(n589), .B(KEYINPUT74), .ZN(n612) );
  NAND2_X1 U677 ( .A1(n612), .A2(n669), .ZN(n590) );
  NOR2_X1 U678 ( .A1(n580), .A2(n590), .ZN(n591) );
  XOR2_X1 U679 ( .A(KEYINPUT28), .B(n591), .Z(n592) );
  NOR2_X1 U680 ( .A1(n593), .A2(n592), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n596) );
  NAND2_X1 U682 ( .A1(n682), .A2(n681), .ZN(n594) );
  XNOR2_X1 U683 ( .A(n596), .B(n595), .ZN(n695) );
  NAND2_X1 U684 ( .A1(n606), .A2(n695), .ZN(n597) );
  XOR2_X1 U685 ( .A(KEYINPUT46), .B(KEYINPUT86), .Z(n598) );
  AND2_X1 U686 ( .A1(n584), .A2(n600), .ZN(n601) );
  XOR2_X1 U687 ( .A(KEYINPUT108), .B(n601), .Z(n602) );
  NOR2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n648) );
  INV_X1 U689 ( .A(n604), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n649) );
  NOR2_X1 U691 ( .A1(n649), .A2(n679), .ZN(n607) );
  XOR2_X1 U692 ( .A(KEYINPUT47), .B(n607), .Z(n608) );
  NOR2_X1 U693 ( .A1(n648), .A2(n608), .ZN(n609) );
  XOR2_X1 U694 ( .A(KEYINPUT36), .B(KEYINPUT90), .Z(n615) );
  NAND2_X1 U695 ( .A1(n669), .A2(n681), .ZN(n610) );
  NOR2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n650), .A2(n614), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n658) );
  NAND2_X1 U700 ( .A1(n619), .A2(n666), .ZN(n620) );
  XNOR2_X1 U701 ( .A(n620), .B(KEYINPUT106), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT43), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n662) );
  NAND2_X1 U704 ( .A1(n625), .A2(KEYINPUT2), .ZN(n626) );
  XNOR2_X1 U705 ( .A(KEYINPUT68), .B(n626), .ZN(n627) );
  NAND2_X1 U706 ( .A1(KEYINPUT2), .A2(n663), .ZN(n628) );
  AND2_X2 U707 ( .A1(n629), .A2(n628), .ZN(n712) );
  NAND2_X1 U708 ( .A1(n712), .A2(G210), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n712), .A2(G472), .ZN(n634) );
  XOR2_X1 U710 ( .A(n631), .B(KEYINPUT62), .Z(n632) );
  XOR2_X1 U711 ( .A(G101), .B(n637), .Z(G3) );
  NAND2_X1 U712 ( .A1(n639), .A2(n653), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n638), .B(G104), .ZN(G6) );
  XOR2_X1 U714 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n641) );
  NAND2_X1 U715 ( .A1(n639), .A2(n655), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n641), .B(n640), .ZN(n643) );
  XOR2_X1 U717 ( .A(G107), .B(KEYINPUT27), .Z(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(G9) );
  XOR2_X1 U719 ( .A(G110), .B(n644), .Z(G12) );
  NOR2_X1 U720 ( .A1(n645), .A2(n649), .ZN(n647) );
  XNOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(G30) );
  XOR2_X1 U723 ( .A(G143), .B(n648), .Z(G45) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U725 ( .A(KEYINPUT114), .B(n651), .Z(n652) );
  XNOR2_X1 U726 ( .A(G146), .B(n652), .ZN(G48) );
  NAND2_X1 U727 ( .A1(n656), .A2(n653), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(G113), .ZN(G15) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(G116), .ZN(G18) );
  XOR2_X1 U731 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n660) );
  XNOR2_X1 U732 ( .A(G125), .B(n658), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(G27) );
  XOR2_X1 U734 ( .A(G134), .B(n661), .Z(G36) );
  XNOR2_X1 U735 ( .A(G140), .B(n662), .ZN(G42) );
  XNOR2_X1 U736 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n706) );
  XNOR2_X1 U737 ( .A(KEYINPUT85), .B(n699), .ZN(n664) );
  NOR2_X1 U738 ( .A1(KEYINPUT2), .A2(n664), .ZN(n704) );
  XOR2_X1 U739 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n668) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(n671), .Z(n672) );
  NAND2_X1 U744 ( .A1(n580), .A2(n672), .ZN(n673) );
  NOR2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n677), .B(KEYINPUT51), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n678), .A2(n695), .ZN(n690) );
  NAND2_X1 U749 ( .A1(n397), .A2(n680), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(KEYINPUT117), .B(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n688), .A2(n694), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U756 ( .A(KEYINPUT52), .B(n691), .Z(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n698) );
  NAND2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U759 ( .A1(n742), .A2(n696), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n699), .A2(KEYINPUT85), .ZN(n700) );
  NAND2_X1 U762 ( .A1(KEYINPUT2), .A2(n700), .ZN(n701) );
  NAND2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U765 ( .A(n706), .B(n705), .ZN(G75) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n709) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT119), .ZN(n708) );
  BUF_X2 U768 ( .A(n712), .Z(n719) );
  NAND2_X1 U769 ( .A1(n719), .A2(G469), .ZN(n710) );
  NOR2_X1 U770 ( .A1(n722), .A2(n711), .ZN(G54) );
  NAND2_X1 U771 ( .A1(n712), .A2(G475), .ZN(n715) );
  XOR2_X1 U772 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n713) );
  XNOR2_X1 U773 ( .A(n716), .B(KEYINPUT122), .ZN(n718) );
  NAND2_X1 U774 ( .A1(G478), .A2(n719), .ZN(n717) );
  NAND2_X1 U775 ( .A1(G217), .A2(n719), .ZN(n720) );
  XNOR2_X1 U776 ( .A(G101), .B(n723), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n725), .B(n724), .ZN(n727) );
  NOR2_X1 U778 ( .A1(G898), .A2(n742), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n737) );
  INV_X1 U780 ( .A(G898), .ZN(n731) );
  NAND2_X1 U781 ( .A1(G224), .A2(G953), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n728), .B(KEYINPUT61), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n729), .B(KEYINPUT123), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n735) );
  BUF_X1 U785 ( .A(n732), .Z(n733) );
  NOR2_X1 U786 ( .A1(G953), .A2(n733), .ZN(n734) );
  NOR2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U788 ( .A(n737), .B(n736), .Z(G69) );
  XOR2_X1 U789 ( .A(KEYINPUT124), .B(n738), .Z(n739) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(n744) );
  XNOR2_X1 U791 ( .A(n744), .B(n741), .ZN(n743) );
  NAND2_X1 U792 ( .A1(n743), .A2(n742), .ZN(n748) );
  XNOR2_X1 U793 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U795 ( .A1(G953), .A2(n746), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U797 ( .A(G122), .B(n749), .Z(G24) );
  XNOR2_X1 U798 ( .A(n750), .B(KEYINPUT125), .ZN(G21) );
  XNOR2_X1 U799 ( .A(G137), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(G39) );
  XOR2_X1 U801 ( .A(n753), .B(G131), .Z(n754) );
  XNOR2_X1 U802 ( .A(KEYINPUT127), .B(n754), .ZN(G33) );
endmodule

