//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  XOR2_X1   g000(.A(KEYINPUT26), .B(G101), .Z(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n187), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n198), .B2(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(new_n199), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G131), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n200), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n209), .A2(new_n211), .A3(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT64), .B1(new_n208), .B2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n210), .A3(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n217), .A3(new_n209), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n207), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT0), .B(G128), .Z(new_n224));
  AOI22_X1  g038(.A1(KEYINPUT0), .A2(new_n212), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n204), .A2(G131), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n206), .A2(new_n203), .A3(new_n199), .A4(new_n202), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n229), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(KEYINPUT71), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT71), .B1(new_n238), .B2(new_n239), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT77), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n239), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n240), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n213), .A2(new_n212), .B1(new_n218), .B2(new_n220), .ZN(new_n250));
  INV_X1    g064(.A(new_n200), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n227), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n207), .A2(new_n222), .A3(KEYINPUT68), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT67), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT67), .B1(new_n225), .B2(new_n228), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n236), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(KEYINPUT76), .A3(new_n236), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n257), .B2(new_n236), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n254), .A2(new_n253), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n229), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n264), .A2(new_n268), .A3(KEYINPUT75), .A4(new_n237), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n260), .A2(new_n261), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  AOI221_X4 g084(.A(new_n194), .B1(new_n243), .B2(new_n248), .C1(new_n270), .C2(KEYINPUT28), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT78), .B1(new_n271), .B2(G902), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n264), .A2(new_n268), .A3(new_n237), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n218), .A2(new_n224), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT0), .A4(G128), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n228), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n223), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n236), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n239), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n246), .A2(new_n240), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n193), .B(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n286), .B2(KEYINPUT73), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n281), .B1(new_n257), .B2(new_n236), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n241), .A2(new_n242), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n193), .B(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(new_n223), .C1(new_n278), .C2(new_n279), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(KEYINPUT30), .B2(new_n257), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n273), .B1(new_n297), .B2(new_n237), .ZN(new_n298));
  INV_X1    g112(.A(new_n193), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n292), .A2(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n287), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n257), .A2(KEYINPUT30), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n237), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  INV_X1    g118(.A(new_n273), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n286), .B2(KEYINPUT73), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n292), .B2(new_n293), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT74), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n311));
  INV_X1    g125(.A(new_n194), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n243), .A2(new_n248), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n272), .A2(new_n302), .A3(new_n310), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G472), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n285), .B1(new_n282), .B2(new_n283), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT72), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n322), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n304), .A2(new_n305), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT31), .B1(new_n324), .B2(new_n193), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n273), .B(new_n193), .C1(new_n297), .C2(new_n237), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT31), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n321), .B(new_n323), .C1(new_n325), .C2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n329), .A2(KEYINPUT32), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT32), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n319), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G214), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n189), .A2(G224), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n225), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n250), .A2(new_n338), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT7), .B(new_n337), .C1(new_n341), .C2(KEYINPUT94), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(KEYINPUT7), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n339), .A2(new_n343), .A3(new_n344), .A4(new_n340), .ZN(new_n345));
  XNOR2_X1  g159(.A(G110), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT8), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT89), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n231), .B2(KEYINPUT5), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT5), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(new_n230), .A3(KEYINPUT89), .A4(G116), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n349), .A2(new_n350), .A3(G113), .A4(new_n352), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n234), .A2(new_n235), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  INV_X1    g170(.A(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT85), .B1(new_n357), .B2(G104), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  OAI211_X1 g175(.A(G101), .B(new_n358), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n357), .A3(G104), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n360), .A2(G107), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n355), .B(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n342), .A2(new_n345), .B1(new_n347), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n362), .A2(new_n368), .A3(KEYINPUT87), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT87), .B1(new_n362), .B2(new_n368), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n372), .B1(new_n375), .B2(new_n355), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n353), .A2(new_n354), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(KEYINPUT90), .C1(new_n374), .C2(new_n373), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G101), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n368), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n382), .A3(G101), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n383), .A3(new_n236), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n376), .A2(new_n346), .A3(new_n378), .A4(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(G902), .B1(new_n371), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n337), .B(KEYINPUT92), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n341), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n376), .A2(new_n378), .A3(new_n384), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n346), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n385), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT6), .B1(new_n389), .B2(new_n391), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT93), .B(new_n388), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n369), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n362), .A2(new_n368), .A3(KEYINPUT87), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n355), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n384), .B1(new_n400), .B2(KEYINPUT90), .ZN(new_n401));
  INV_X1    g215(.A(new_n378), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n385), .A3(new_n392), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT93), .B1(new_n406), .B2(new_n388), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n386), .B1(new_n396), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT93), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n395), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n409), .A3(new_n386), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n336), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n250), .A2(new_n369), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n209), .A2(new_n211), .ZN(new_n419));
  INV_X1    g233(.A(G128), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(KEYINPUT1), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n219), .A2(G128), .B1(new_n209), .B2(new_n211), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n368), .B(new_n362), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n228), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT12), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(new_n228), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT10), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n212), .A2(new_n213), .B1(new_n220), .B2(new_n419), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(new_n369), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT10), .B(new_n222), .C1(new_n373), .C2(new_n374), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n423), .A2(KEYINPUT86), .A3(new_n430), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n381), .A2(new_n383), .A3(new_n225), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(new_n228), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT84), .B1(new_n429), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n189), .A2(G227), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n441), .B(new_n442), .Z(new_n443));
  XNOR2_X1  g257(.A(new_n438), .B(new_n228), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n429), .A2(new_n439), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G469), .ZN(new_n450));
  INV_X1    g264(.A(new_n429), .ZN(new_n451));
  INV_X1    g265(.A(new_n439), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n443), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n438), .A2(new_n228), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n446), .B1(new_n454), .B2(new_n439), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n447), .A2(KEYINPUT88), .A3(new_n443), .ZN(new_n458));
  INV_X1    g272(.A(G469), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n316), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n316), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n450), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G137), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n230), .A2(G128), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT23), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n420), .A2(G119), .ZN(new_n470));
  MUX2_X1   g284(.A(KEYINPUT23), .B(new_n469), .S(new_n470), .Z(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G110), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n468), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT24), .B(G110), .ZN(new_n474));
  OR3_X1    g288(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT79), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT79), .B1(new_n473), .B2(new_n474), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G125), .B(G140), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT80), .A3(KEYINPUT16), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n481));
  INV_X1    g295(.A(G140), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G125), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n478), .A2(KEYINPUT16), .B1(KEYINPUT80), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n480), .A2(new_n484), .A3(new_n210), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(KEYINPUT80), .ZN(new_n486));
  XOR2_X1   g300(.A(G125), .B(G140), .Z(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n481), .ZN(new_n488));
  AOI21_X1  g302(.A(G146), .B1(new_n488), .B2(new_n479), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n472), .B(new_n477), .C1(new_n485), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n473), .A2(new_n474), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n471), .B2(G110), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n478), .A2(new_n210), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(G146), .A3(new_n479), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n490), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n491), .B1(new_n490), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n467), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n496), .A3(new_n466), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n316), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G217), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(new_n316), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n503), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n499), .A2(KEYINPUT25), .A3(new_n316), .A4(new_n500), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT82), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n499), .A2(new_n500), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n506), .A2(G902), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT83), .Z(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT9), .B(G234), .ZN(new_n516));
  OAI21_X1  g330(.A(G221), .B1(new_n516), .B2(G902), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n463), .A2(new_n511), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G475), .ZN(new_n519));
  INV_X1    g333(.A(G214), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n520), .A2(G237), .A3(G953), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT96), .B1(new_n522), .B2(G143), .ZN(new_n523));
  OR2_X1    g337(.A1(KEYINPUT96), .A2(G143), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n208), .A2(KEYINPUT95), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(KEYINPUT96), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n206), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  INV_X1    g345(.A(new_n206), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(new_n532), .A3(new_n528), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n210), .B1(new_n480), .B2(new_n484), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n525), .A2(new_n532), .A3(new_n528), .A4(KEYINPUT17), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n495), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n360), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n487), .A2(G146), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n494), .ZN(new_n541));
  AND2_X1   g355(.A1(KEYINPUT18), .A2(G131), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n529), .A2(KEYINPUT97), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n529), .B2(KEYINPUT97), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n537), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n530), .A2(new_n533), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n478), .A2(KEYINPUT98), .A3(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT19), .B1(new_n478), .B2(KEYINPUT98), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n210), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n495), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n539), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n519), .B(new_n316), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n539), .B1(new_n537), .B2(new_n545), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n316), .B1(new_n546), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n545), .A2(new_n551), .ZN(new_n559));
  INV_X1    g373(.A(new_n539), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n537), .A2(new_n539), .A3(new_n545), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n519), .A4(new_n316), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n555), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n189), .A2(G952), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(G234), .B2(G237), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT21), .B(G898), .Z(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(G234), .A2(G237), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(G902), .A3(G953), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G478), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(KEYINPUT15), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT13), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n420), .B2(G143), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n208), .A2(G128), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT100), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n420), .A2(G143), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n208), .A2(KEYINPUT13), .A3(G128), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G134), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n586), .A3(new_n198), .ZN(new_n590));
  XNOR2_X1  g404(.A(G116), .B(G122), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n357), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n232), .A2(KEYINPUT14), .A3(G122), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  OAI211_X1 g409(.A(G107), .B(new_n594), .C1(new_n595), .C2(KEYINPUT14), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n357), .ZN(new_n597));
  INV_X1    g411(.A(new_n590), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n198), .B1(new_n584), .B2(new_n586), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n516), .A2(new_n505), .A3(G953), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n593), .A2(new_n600), .A3(new_n602), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n579), .B1(new_n606), .B2(new_n316), .ZN(new_n607));
  AOI211_X1 g421(.A(G902), .B(new_n578), .C1(new_n604), .C2(new_n605), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n555), .A2(new_n558), .A3(new_n564), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT99), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n567), .A2(new_n576), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n518), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n334), .A2(new_n417), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  NAND2_X1  g429(.A1(new_n329), .A2(new_n316), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n616), .A2(G472), .B1(new_n330), .B2(new_n329), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n463), .A2(new_n517), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n511), .A2(new_n515), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n617), .A2(new_n619), .A3(KEYINPUT101), .A4(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n409), .B1(new_n415), .B2(new_n386), .ZN(new_n623));
  INV_X1    g437(.A(new_n386), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n410), .B(new_n624), .C1(new_n414), .C2(new_n395), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n335), .B(new_n576), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(G478), .B(G902), .C1(new_n604), .C2(new_n605), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n606), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n604), .A2(KEYINPUT33), .A3(new_n605), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n316), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n627), .B1(new_n631), .B2(G478), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT102), .Z(new_n633));
  NAND2_X1  g447(.A1(new_n567), .A2(new_n611), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n329), .A2(new_n330), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n321), .A2(new_n323), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n326), .B(new_n327), .ZN(new_n640));
  AOI21_X1  g454(.A(G902), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G472), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n637), .B1(new_n643), .B2(new_n518), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n622), .A2(new_n636), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NOR2_X1   g461(.A1(new_n610), .A2(new_n609), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n622), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(new_n626), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n634), .A2(new_n607), .A3(new_n608), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n497), .A2(new_n498), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n467), .A2(KEYINPUT36), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n656), .B(new_n657), .Z(new_n658));
  AOI22_X1  g472(.A1(new_n507), .A2(new_n510), .B1(new_n514), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n618), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n654), .A2(new_n655), .A3(new_n660), .A4(new_n617), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  XOR2_X1   g477(.A(new_n569), .B(KEYINPUT103), .Z(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(new_n574), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n649), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n334), .A2(new_n417), .A3(new_n660), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  NAND2_X1  g483(.A1(new_n411), .A2(new_n416), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT38), .Z(new_n671));
  INV_X1    g485(.A(new_n634), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n671), .A2(new_n336), .A3(new_n609), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n326), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n285), .B2(new_n270), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n333), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n666), .B(KEYINPUT39), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n619), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n659), .A3(new_n677), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NOR2_X1   g497(.A1(new_n635), .A2(new_n666), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n334), .A2(new_n417), .A3(new_n660), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NAND3_X1  g500(.A1(new_n457), .A2(new_n316), .A3(new_n458), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n517), .A3(new_n460), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n334), .A2(new_n636), .A3(new_n621), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  AOI21_X1  g507(.A(new_n620), .B1(new_n319), .B2(new_n333), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n650), .A3(new_n690), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR3_X1   g510(.A1(new_n689), .A2(new_n659), .A3(new_n612), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n334), .A2(new_n417), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  AND2_X1   g513(.A1(new_n417), .A2(new_n690), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n641), .A2(new_n642), .ZN(new_n701));
  INV_X1    g515(.A(new_n330), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n270), .A2(KEYINPUT28), .B1(new_n243), .B2(new_n248), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n703), .A2(new_n291), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n704), .B2(new_n640), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n701), .A2(new_n620), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n672), .A2(new_n609), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n700), .A2(new_n706), .A3(new_n576), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NOR3_X1   g523(.A1(new_n701), .A2(new_n659), .A3(new_n705), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n700), .A2(new_n710), .A3(new_n684), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT105), .B(G125), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G27));
  NAND3_X1  g527(.A1(new_n411), .A2(new_n335), .A3(new_n416), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n618), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n334), .A2(new_n621), .A3(new_n684), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n684), .A4(new_n715), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G131), .ZN(G33));
  NAND4_X1  g535(.A1(new_n334), .A2(new_n621), .A3(new_n667), .A4(new_n715), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  NAND2_X1  g537(.A1(new_n672), .A2(new_n633), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT43), .ZN(new_n725));
  INV_X1    g539(.A(new_n659), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(KEYINPUT43), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(new_n643), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(KEYINPUT108), .Z(new_n731));
  INV_X1    g545(.A(new_n714), .ZN(new_n732));
  NAND2_X1  g546(.A1(KEYINPUT45), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n450), .A2(KEYINPUT106), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n449), .A2(KEYINPUT45), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(G469), .C1(new_n449), .C2(KEYINPUT45), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n462), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n460), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n743), .B(KEYINPUT46), .C1(new_n738), .C2(new_n462), .ZN(new_n744));
  OR3_X1    g558(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(new_n517), .A3(new_n678), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n728), .A2(new_n729), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n731), .A2(new_n732), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G137), .ZN(G39));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n750), .A3(new_n517), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n752));
  INV_X1    g566(.A(new_n517), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT47), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n333), .A2(new_n751), .A3(new_n319), .A4(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n620), .A3(new_n684), .A4(new_n732), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  OR2_X1    g571(.A1(G952), .A2(G953), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n710), .A2(new_n684), .A3(new_n715), .ZN(new_n760));
  INV_X1    g574(.A(new_n666), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n565), .A2(KEYINPUT109), .A3(new_n609), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n555), .A2(new_n609), .A3(new_n558), .A4(new_n564), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n666), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n335), .A2(new_n766), .A3(new_n411), .A4(new_n416), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n334), .A2(KEYINPUT110), .A3(new_n660), .A4(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n722), .A2(new_n768), .ZN(new_n769));
  AOI211_X1 g583(.A(KEYINPUT78), .B(G902), .C1(new_n703), .C2(new_n312), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT74), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n301), .B1(new_n287), .B2(new_n300), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n642), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT32), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n638), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n329), .A2(KEYINPUT32), .A3(new_n330), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n767), .B(new_n660), .C1(new_n776), .C2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n720), .A2(new_n760), .A3(new_n769), .A4(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n691), .A2(new_n708), .A3(new_n698), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n672), .A2(new_n633), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n655), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n622), .A2(new_n644), .A3(new_n787), .A4(new_n654), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(new_n614), .A3(new_n661), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n789), .A3(new_n695), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n759), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n783), .A2(new_n722), .A3(new_n768), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n718), .B2(new_n719), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n695), .A2(new_n691), .A3(new_n698), .A4(new_n708), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n788), .A2(new_n614), .A3(new_n661), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n796), .A4(new_n760), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n707), .A2(new_n335), .A3(new_n670), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n618), .A2(new_n666), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n677), .A3(new_n659), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n668), .A3(new_n685), .A4(new_n711), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n791), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n791), .A2(new_n797), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT54), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n725), .A2(new_n664), .A3(new_n727), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n706), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n700), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n806), .A2(new_n815), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n808), .A2(new_n790), .A3(new_n784), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n810), .B(new_n814), .C1(new_n819), .C2(KEYINPUT54), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n677), .A2(new_n620), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n569), .A2(new_n821), .A3(new_n690), .A4(new_n732), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n633), .A2(new_n634), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n811), .A2(new_n690), .A3(new_n732), .ZN(new_n826));
  INV_X1    g640(.A(new_n710), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n671), .A2(new_n336), .A3(new_n690), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n813), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n833), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT50), .B1(new_n833), .B2(KEYINPUT115), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n688), .A2(new_n460), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n751), .A2(new_n754), .B1(new_n753), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n714), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n841), .B2(new_n813), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n840), .A2(KEYINPUT113), .A3(new_n714), .A4(new_n812), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n829), .B(new_n836), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n694), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n826), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT48), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n822), .A2(new_n634), .A3(new_n633), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT116), .B1(new_n825), .B2(new_n828), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n824), .B(new_n852), .C1(new_n827), .C2(new_n826), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n834), .A3(new_n835), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n845), .B1(new_n841), .B2(new_n813), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n568), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n846), .A2(new_n849), .A3(new_n850), .A4(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n758), .B1(new_n820), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n838), .A2(KEYINPUT49), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n838), .A2(KEYINPUT49), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n860), .A2(new_n724), .A3(new_n861), .A4(new_n753), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n821), .A3(new_n335), .A4(new_n671), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(KEYINPUT117), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(G75));
  XNOR2_X1  g682(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n819), .A2(G210), .A3(G902), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n406), .B(new_n388), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n870), .A2(new_n871), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n872), .ZN(new_n878));
  INV_X1    g692(.A(new_n869), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n189), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n876), .A2(new_n881), .A3(new_n883), .ZN(G51));
  XNOR2_X1  g698(.A(new_n819), .B(KEYINPUT54), .ZN(new_n885));
  XOR2_X1   g699(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n461), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n886), .A2(new_n461), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n457), .A2(new_n458), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n819), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n738), .B(KEYINPUT120), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n882), .B1(new_n892), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n562), .A3(new_n561), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(new_n563), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n898), .A2(new_n883), .A3(new_n899), .ZN(G60));
  XNOR2_X1  g714(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n577), .A2(new_n316), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n629), .A2(new_n630), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT121), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n819), .A2(KEYINPUT54), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n819), .A2(KEYINPUT54), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n903), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n810), .B1(new_n819), .B2(KEYINPUT54), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n905), .B1(new_n911), .B2(new_n903), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n882), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n885), .A2(KEYINPUT123), .A3(new_n903), .A4(new_n905), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n819), .A2(new_n658), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n883), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n512), .B1(new_n819), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g737(.A(G224), .ZN(new_n924));
  OAI21_X1  g738(.A(G953), .B1(new_n571), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n796), .B2(G953), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT124), .ZN(new_n927));
  INV_X1    g741(.A(new_n406), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(G898), .B2(new_n189), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G69));
  NOR2_X1   g744(.A1(new_n548), .A2(new_n549), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT125), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n297), .B(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n756), .A2(new_n748), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n694), .A2(new_n678), .A3(new_n715), .A4(new_n787), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n668), .A2(new_n685), .A3(new_n711), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n682), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  AND3_X1   g753(.A1(new_n934), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n933), .B1(new_n940), .B2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n665), .A2(G953), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT126), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n934), .A2(new_n722), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n936), .B1(new_n718), .B2(new_n719), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n746), .A2(new_n694), .A3(new_n798), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n947), .B2(new_n189), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n948), .B2(new_n933), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n950), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n941), .B(new_n952), .C1(new_n948), .C2(new_n933), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(G72));
  NAND4_X1  g768(.A1(new_n944), .A2(new_n796), .A3(new_n945), .A4(new_n946), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  AOI21_X1  g771(.A(new_n193), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n940), .A2(new_n796), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n324), .B1(new_n959), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n306), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n306), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n962), .A2(new_n674), .A3(KEYINPUT127), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n809), .A2(new_n957), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n961), .A2(new_n883), .A3(new_n965), .ZN(G57));
endmodule


