

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(G160), .A2(G40), .ZN(n775) );
  NOR2_X2 U552 ( .A1(n530), .A2(n529), .ZN(G160) );
  XOR2_X1 U553 ( .A(KEYINPUT66), .B(n523), .Z(n516) );
  XOR2_X1 U554 ( .A(KEYINPUT31), .B(n696), .Z(n517) );
  OR2_X1 U555 ( .A1(n752), .A2(KEYINPUT33), .ZN(n518) );
  INV_X1 U556 ( .A(n690), .ZN(n715) );
  NOR2_X1 U557 ( .A1(G1966), .A2(n771), .ZN(n742) );
  NOR2_X1 U558 ( .A1(n751), .A2(n771), .ZN(n752) );
  AND2_X1 U559 ( .A1(n755), .A2(n987), .ZN(n756) );
  NAND2_X1 U560 ( .A1(n774), .A2(n681), .ZN(n690) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n774) );
  INV_X1 U562 ( .A(G2104), .ZN(n525) );
  NOR2_X2 U563 ( .A1(n633), .A2(n544), .ZN(n649) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n525), .ZN(n885) );
  NOR2_X1 U565 ( .A1(G651), .A2(n633), .ZN(n653) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n519), .Z(n886) );
  NAND2_X1 U568 ( .A1(G137), .A2(n886), .ZN(n520) );
  XNOR2_X1 U569 ( .A(n520), .B(KEYINPUT68), .ZN(n524) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(KEYINPUT67), .Z(n522) );
  NAND2_X1 U571 ( .A1(G101), .A2(n885), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n516), .ZN(n530) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U575 ( .A1(G113), .A2(n889), .ZN(n528) );
  NAND2_X1 U576 ( .A1(n525), .A2(G2105), .ZN(n526) );
  XNOR2_X2 U577 ( .A(n526), .B(KEYINPUT65), .ZN(n891) );
  NAND2_X1 U578 ( .A1(G125), .A2(n891), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n886), .A2(G138), .ZN(n531) );
  XOR2_X1 U581 ( .A(KEYINPUT93), .B(n531), .Z(n538) );
  NAND2_X1 U582 ( .A1(G126), .A2(n891), .ZN(n532) );
  XNOR2_X1 U583 ( .A(n532), .B(KEYINPUT92), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G114), .A2(n889), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G102), .A2(n885), .ZN(n533) );
  AND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(G164) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G82), .ZN(G220) );
  INV_X1 U591 ( .A(G57), .ZN(G237) );
  INV_X1 U592 ( .A(G108), .ZN(G238) );
  INV_X1 U593 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U594 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n543) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n648) );
  NAND2_X1 U596 ( .A1(G90), .A2(n648), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  INV_X1 U598 ( .A(G651), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G77), .A2(n649), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n541), .B(KEYINPUT9), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n543), .B(n542), .ZN(n549) );
  NOR2_X1 U603 ( .A1(G543), .A2(n544), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT1), .B(n545), .Z(n652) );
  NAND2_X1 U605 ( .A1(G64), .A2(n652), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G52), .A2(n653), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U608 ( .A1(n549), .A2(n548), .ZN(G171) );
  INV_X1 U609 ( .A(G171), .ZN(G301) );
  NAND2_X1 U610 ( .A1(n649), .A2(G76), .ZN(n550) );
  XNOR2_X1 U611 ( .A(KEYINPUT80), .B(n550), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n648), .A2(G89), .ZN(n551) );
  XNOR2_X1 U613 ( .A(KEYINPUT4), .B(n551), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G63), .A2(n652), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G51), .A2(n653), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U623 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n562) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n562), .B(n561), .ZN(G223) );
  INV_X1 U626 ( .A(G223), .ZN(n838) );
  NAND2_X1 U627 ( .A1(n838), .A2(G567), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U629 ( .A1(n648), .A2(G81), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G68), .A2(n649), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT13), .B(KEYINPUT78), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n652), .A2(G56), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n569), .Z(n570) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n653), .A2(G43), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n977) );
  INV_X1 U640 ( .A(G860), .ZN(n596) );
  OR2_X1 U641 ( .A1(n977), .A2(n596), .ZN(G153) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n653), .A2(G54), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G92), .A2(n648), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G66), .A2(n652), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G79), .A2(n649), .ZN(n576) );
  XNOR2_X1 U648 ( .A(KEYINPUT79), .B(n576), .ZN(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X2 U651 ( .A(KEYINPUT15), .B(n581), .Z(n969) );
  INV_X1 U652 ( .A(G868), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n969), .A2(n592), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U655 ( .A1(n649), .A2(G78), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n584), .B(KEYINPUT74), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G91), .A2(n648), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(n587), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G65), .A2(n652), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G53), .A2(n653), .ZN(n588) );
  AND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(G299) );
  NOR2_X1 U664 ( .A1(G286), .A2(n592), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT81), .B(n593), .Z(n595) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n596), .A2(G559), .ZN(n597) );
  INV_X1 U669 ( .A(n969), .ZN(n643) );
  NAND2_X1 U670 ( .A1(n597), .A2(n643), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U672 ( .A1(n643), .A2(G868), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G559), .A2(n599), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT82), .ZN(n602) );
  NOR2_X1 U675 ( .A1(n977), .A2(G868), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G111), .A2(n889), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G99), .A2(n885), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n611) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n606) );
  NAND2_X1 U681 ( .A1(G123), .A2(n891), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U683 ( .A(KEYINPUT83), .B(n607), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n886), .A2(G135), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n1003) );
  XNOR2_X1 U687 ( .A(n1003), .B(G2096), .ZN(n613) );
  INV_X1 U688 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G85), .A2(n648), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G72), .A2(n649), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U693 ( .A(KEYINPUT69), .B(n616), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G47), .A2(n653), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT71), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G60), .A2(n652), .ZN(n618) );
  XOR2_X1 U697 ( .A(KEYINPUT70), .B(n618), .Z(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G290) );
  NAND2_X1 U700 ( .A1(G62), .A2(n652), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G50), .A2(n653), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U703 ( .A(KEYINPUT86), .B(n625), .Z(n629) );
  NAND2_X1 U704 ( .A1(G88), .A2(n648), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G75), .A2(n649), .ZN(n626) );
  AND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G303) );
  INV_X1 U708 ( .A(G303), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G49), .A2(n653), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U712 ( .A1(n652), .A2(n632), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n633), .A2(G87), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G86), .A2(n648), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G61), .A2(n652), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n649), .A2(G73), .ZN(n638) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n653), .A2(G48), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G559), .A2(n643), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(n977), .ZN(n845) );
  XNOR2_X1 U725 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n646) );
  XNOR2_X1 U726 ( .A(G288), .B(KEYINPUT19), .ZN(n645) );
  XNOR2_X1 U727 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U728 ( .A(G166), .B(n647), .ZN(n661) );
  INV_X1 U729 ( .A(G299), .ZN(n986) );
  NAND2_X1 U730 ( .A1(G93), .A2(n648), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G80), .A2(n649), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U733 ( .A1(G67), .A2(n652), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G55), .A2(n653), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U737 ( .A(KEYINPUT85), .B(n658), .Z(n846) );
  XNOR2_X1 U738 ( .A(n986), .B(n846), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n659), .B(G305), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U741 ( .A(G290), .B(n662), .Z(n911) );
  XNOR2_X1 U742 ( .A(n845), .B(n911), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G868), .ZN(n665) );
  OR2_X1 U744 ( .A1(G868), .A2(n846), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U752 ( .A(KEYINPUT76), .B(G132), .Z(G219) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U754 ( .A1(G236), .A2(G238), .ZN(n670) );
  NAND2_X1 U755 ( .A1(G69), .A2(n670), .ZN(n671) );
  NOR2_X1 U756 ( .A1(n671), .A2(G237), .ZN(n672) );
  XNOR2_X1 U757 ( .A(n672), .B(KEYINPUT89), .ZN(n843) );
  NAND2_X1 U758 ( .A1(n843), .A2(G567), .ZN(n677) );
  NOR2_X1 U759 ( .A1(G219), .A2(G220), .ZN(n673) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U761 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U762 ( .A1(G96), .A2(n675), .ZN(n844) );
  NAND2_X1 U763 ( .A1(n844), .A2(G2106), .ZN(n676) );
  NAND2_X1 U764 ( .A1(n677), .A2(n676), .ZN(n848) );
  NOR2_X1 U765 ( .A1(n678), .A2(n848), .ZN(n679) );
  XNOR2_X1 U766 ( .A(n679), .B(KEYINPUT90), .ZN(n841) );
  NAND2_X1 U767 ( .A1(n841), .A2(G36), .ZN(n680) );
  XOR2_X1 U768 ( .A(KEYINPUT91), .B(n680), .Z(G176) );
  INV_X1 U769 ( .A(n775), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G8), .A2(n690), .ZN(n771) );
  INV_X1 U771 ( .A(n742), .ZN(n685) );
  NOR2_X1 U772 ( .A1(n775), .A2(G2084), .ZN(n682) );
  AND2_X1 U773 ( .A1(n682), .A2(n774), .ZN(n683) );
  XOR2_X1 U774 ( .A(KEYINPUT103), .B(n683), .Z(n741) );
  INV_X1 U775 ( .A(n741), .ZN(n684) );
  NAND2_X1 U776 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n686), .B(KEYINPUT105), .ZN(n687) );
  NAND2_X1 U778 ( .A1(n687), .A2(G8), .ZN(n688) );
  XNOR2_X1 U779 ( .A(n688), .B(KEYINPUT30), .ZN(n689) );
  NOR2_X1 U780 ( .A1(G168), .A2(n689), .ZN(n695) );
  XOR2_X1 U781 ( .A(KEYINPUT25), .B(G2078), .Z(n952) );
  NAND2_X1 U782 ( .A1(n715), .A2(n952), .ZN(n692) );
  INV_X1 U783 ( .A(n715), .ZN(n728) );
  NAND2_X1 U784 ( .A1(G1961), .A2(n728), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U786 ( .A(KEYINPUT104), .B(n693), .Z(n697) );
  NOR2_X1 U787 ( .A1(G171), .A2(n697), .ZN(n694) );
  NOR2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(G171), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n728), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n715), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n969), .A2(n700), .ZN(n714) );
  NAND2_X1 U794 ( .A1(G1348), .A2(n969), .ZN(n701) );
  XNOR2_X1 U795 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n701), .A2(n706), .ZN(n702) );
  NOR2_X1 U797 ( .A1(G1341), .A2(n702), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n715), .A2(n703), .ZN(n705) );
  NOR2_X1 U799 ( .A1(G1996), .A2(n706), .ZN(n704) );
  NOR2_X1 U800 ( .A1(n705), .A2(n704), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n969), .A2(G2067), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G1996), .A2(n706), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n709), .A2(n715), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n977), .A2(n712), .ZN(n713) );
  NOR2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n715), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U809 ( .A(n716), .B(KEYINPUT27), .ZN(n718) );
  AND2_X1 U810 ( .A1(G1956), .A2(n728), .ZN(n717) );
  NOR2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n721), .A2(n986), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n724) );
  NOR2_X1 U814 ( .A1(n721), .A2(n986), .ZN(n722) );
  XOR2_X1 U815 ( .A(n722), .B(KEYINPUT28), .Z(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U817 ( .A(KEYINPUT29), .B(n725), .Z(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n740) );
  INV_X1 U819 ( .A(G8), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n771), .ZN(n730) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U823 ( .A1(n731), .A2(G303), .ZN(n732) );
  OR2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n735) );
  AND2_X1 U825 ( .A1(n740), .A2(n735), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n517), .A2(n734), .ZN(n738) );
  INV_X1 U827 ( .A(n735), .ZN(n736) );
  OR2_X1 U828 ( .A1(n736), .A2(G286), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U830 ( .A(n739), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n517), .A2(n740), .ZN(n745) );
  AND2_X1 U832 ( .A1(G8), .A2(n741), .ZN(n743) );
  NOR2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n759) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n975) );
  AND2_X1 U836 ( .A1(n759), .A2(n975), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n758), .A2(n746), .ZN(n750) );
  INV_X1 U838 ( .A(n975), .ZN(n748) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U841 ( .A1(n753), .A2(n747), .ZN(n981) );
  OR2_X1 U842 ( .A1(n748), .A2(n981), .ZN(n749) );
  AND2_X1 U843 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  OR2_X1 U845 ( .A1(n771), .A2(n754), .ZN(n755) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n987) );
  NAND2_X1 U847 ( .A1(n518), .A2(n756), .ZN(n757) );
  XNOR2_X1 U848 ( .A(n757), .B(KEYINPUT106), .ZN(n766) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n762) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U851 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U853 ( .A(KEYINPUT107), .B(n763), .Z(n764) );
  NAND2_X1 U854 ( .A1(n764), .A2(n771), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n773) );
  XNOR2_X1 U856 ( .A(KEYINPUT24), .B(KEYINPUT102), .ZN(n767) );
  XNOR2_X1 U857 ( .A(n767), .B(KEYINPUT101), .ZN(n769) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n780) );
  NOR2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U863 ( .A(n776), .B(KEYINPUT94), .ZN(n824) );
  NOR2_X1 U864 ( .A1(G290), .A2(G1986), .ZN(n813) );
  INV_X1 U865 ( .A(n813), .ZN(n976) );
  NAND2_X1 U866 ( .A1(G1986), .A2(G290), .ZN(n972) );
  NAND2_X1 U867 ( .A1(n976), .A2(n972), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n824), .A2(n777), .ZN(n778) );
  XNOR2_X1 U869 ( .A(n778), .B(KEYINPUT95), .ZN(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n811) );
  NAND2_X1 U871 ( .A1(G107), .A2(n889), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G95), .A2(n885), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G131), .A2(n886), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G119), .A2(n891), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n904) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n904), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT96), .ZN(n799) );
  NAND2_X1 U880 ( .A1(G117), .A2(n889), .ZN(n789) );
  NAND2_X1 U881 ( .A1(G129), .A2(n891), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U883 ( .A(KEYINPUT97), .B(n790), .Z(n793) );
  NAND2_X1 U884 ( .A1(n885), .A2(G105), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n794), .B(KEYINPUT98), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G141), .A2(n886), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U890 ( .A(KEYINPUT99), .B(n797), .Z(n907) );
  NAND2_X1 U891 ( .A1(G1996), .A2(n907), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n1016) );
  NAND2_X1 U893 ( .A1(n824), .A2(n1016), .ZN(n812) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n821) );
  NAND2_X1 U895 ( .A1(G104), .A2(n885), .ZN(n801) );
  NAND2_X1 U896 ( .A1(G140), .A2(n886), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n802), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G116), .A2(n889), .ZN(n804) );
  NAND2_X1 U900 ( .A1(G128), .A2(n891), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n805), .Z(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n808), .ZN(n899) );
  NOR2_X1 U905 ( .A1(n821), .A2(n899), .ZN(n1005) );
  NAND2_X1 U906 ( .A1(n1005), .A2(n824), .ZN(n819) );
  NAND2_X1 U907 ( .A1(n812), .A2(n819), .ZN(n809) );
  XOR2_X1 U908 ( .A(KEYINPUT100), .B(n809), .Z(n810) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n826) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n907), .ZN(n1009) );
  INV_X1 U911 ( .A(n812), .ZN(n816) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n904), .ZN(n1004) );
  NOR2_X1 U913 ( .A1(n813), .A2(n1004), .ZN(n814) );
  XNOR2_X1 U914 ( .A(n814), .B(KEYINPUT108), .ZN(n815) );
  NOR2_X1 U915 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n1009), .A2(n817), .ZN(n818) );
  XNOR2_X1 U917 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n821), .A2(n899), .ZN(n1013) );
  NAND2_X1 U920 ( .A1(n822), .A2(n1013), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U924 ( .A(KEYINPUT109), .B(G2427), .Z(n829) );
  XNOR2_X1 U925 ( .A(G2435), .B(G2438), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n836) );
  XOR2_X1 U927 ( .A(G2443), .B(G2430), .Z(n831) );
  XNOR2_X1 U928 ( .A(G2454), .B(G2446), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U930 ( .A(n832), .B(G2451), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1348), .B(G1341), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n837), .A2(G14), .ZN(n915) );
  XOR2_X1 U935 ( .A(KEYINPUT110), .B(n915), .Z(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U938 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT111), .B(n840), .Z(n842) );
  NAND2_X1 U941 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  NOR2_X1 U944 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  NOR2_X1 U946 ( .A1(n845), .A2(G860), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G145) );
  INV_X1 U948 ( .A(n848), .ZN(G319) );
  XNOR2_X1 U949 ( .A(G1996), .B(KEYINPUT41), .ZN(n858) );
  XOR2_X1 U950 ( .A(G1981), .B(G1966), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1991), .B(G1986), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U954 ( .A(G1961), .B(G1956), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(G2474), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(G229) );
  XOR2_X1 U960 ( .A(G2678), .B(KEYINPUT42), .Z(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U963 ( .A(KEYINPUT112), .B(G2090), .Z(n862) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2072), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U966 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U967 ( .A(G2096), .B(G2100), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U969 ( .A(G2078), .B(G2084), .Z(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(G227) );
  NAND2_X1 U971 ( .A1(G112), .A2(n889), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G100), .A2(n885), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G124), .A2(n891), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT44), .B(n871), .Z(n872) );
  XNOR2_X1 U976 ( .A(n872), .B(KEYINPUT115), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G136), .A2(n886), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G118), .A2(n889), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G130), .A2(n891), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G106), .A2(n885), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G142), .A2(n886), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U986 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U988 ( .A(KEYINPUT48), .B(n884), .Z(n903) );
  NAND2_X1 U989 ( .A1(G103), .A2(n885), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G139), .A2(n886), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n896) );
  NAND2_X1 U992 ( .A1(n889), .A2(G115), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n890), .B(KEYINPUT116), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n998) );
  XNOR2_X1 U998 ( .A(n998), .B(G162), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n897), .B(n1003), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(G164), .B(G160), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n904), .B(KEYINPUT46), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1006 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1008 ( .A(G286), .B(G301), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n910), .B(n977), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n969), .B(n911), .Z(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n914), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1021 ( .A(G24), .B(G1986), .Z(n923) );
  XNOR2_X1 U1022 ( .A(G1971), .B(G22), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(n921), .B(KEYINPUT125), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G23), .B(G1976), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1027 ( .A(KEYINPUT58), .B(n926), .Z(n943) );
  XOR2_X1 U1028 ( .A(G1966), .B(G21), .Z(n937) );
  XOR2_X1 U1029 ( .A(KEYINPUT123), .B(G4), .Z(n928) );
  XNOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .ZN(n927) );
  XNOR2_X1 U1031 ( .A(n928), .B(n927), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(G6), .B(G1981), .ZN(n929) );
  NOR2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(G20), .B(G1956), .ZN(n933) );
  NOR2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1038 ( .A(KEYINPUT60), .B(n935), .ZN(n936) );
  NAND2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(G5), .B(G1961), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(KEYINPUT122), .B(n938), .ZN(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1043 ( .A(KEYINPUT124), .B(n941), .Z(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1045 ( .A(n944), .B(KEYINPUT61), .Z(n945) );
  XNOR2_X1 U1046 ( .A(KEYINPUT126), .B(n945), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(G16), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(n947), .ZN(n1029) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n1021) );
  XNOR2_X1 U1050 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(n948), .B(KEYINPUT54), .ZN(n961) );
  XOR2_X1 U1052 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1053 ( .A1(n949), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G1996), .B(G32), .ZN(n951) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1056 ( .A1(n951), .A2(n950), .ZN(n956) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1058 ( .A(G27), .B(n952), .ZN(n953) );
  NOR2_X1 U1059 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1060 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1062 ( .A(n959), .B(KEYINPUT53), .ZN(n960) );
  NOR2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1064 ( .A(G2090), .B(KEYINPUT118), .Z(n962) );
  XNOR2_X1 U1065 ( .A(G35), .B(n962), .ZN(n963) );
  NAND2_X1 U1066 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1067 ( .A(n1021), .B(n965), .ZN(n967) );
  INV_X1 U1068 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1069 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n968), .ZN(n1027) );
  XNOR2_X1 U1071 ( .A(G1348), .B(KEYINPUT120), .ZN(n970) );
  XNOR2_X1 U1072 ( .A(n970), .B(n969), .ZN(n974) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1074 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1075 ( .A1(n974), .A2(n973), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G301), .B(G1961), .ZN(n979) );
  XNOR2_X1 U1078 ( .A(n977), .B(G1341), .ZN(n978) );
  NOR2_X1 U1079 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1080 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n986), .B(G1956), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(n989), .B(KEYINPUT57), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(n994), .B(KEYINPUT121), .ZN(n997) );
  XOR2_X1 U1090 ( .A(G16), .B(KEYINPUT56), .Z(n995) );
  XNOR2_X1 U1091 ( .A(KEYINPUT119), .B(n995), .ZN(n996) );
  NAND2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n1025) );
  XOR2_X1 U1093 ( .A(G2072), .B(n998), .Z(n1000) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1001), .Z(n1019) );
  XOR2_X1 U1097 ( .A(G2084), .B(G160), .Z(n1002) );
  NOR2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(G2090), .B(G162), .Z(n1008) );
  NOR2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(n1010), .B(KEYINPUT51), .ZN(n1011) );
  NOR2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT117), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

