//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1383,
    new_n1384, new_n1385;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n217), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n216), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n207), .A2(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n202), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT73), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n213), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n254), .B1(new_n253), .B2(new_n256), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT11), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT11), .B1(new_n257), .B2(new_n258), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n213), .A3(new_n255), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n207), .A2(G1), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n264), .A2(new_n217), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT12), .B1(new_n263), .B2(G68), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n261), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n206), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G238), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n276), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G226), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n226), .A2(G1698), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n287), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G97), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n285), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT71), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n298), .B(new_n285), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n284), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n271), .B1(new_n300), .B2(KEYINPUT13), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n284), .B(new_n302), .C1(new_n297), .C2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G226), .A2(G1698), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n226), .B2(G1698), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT3), .B(G33), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(new_n307), .B1(G33), .B2(G97), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n298), .B1(new_n308), .B2(new_n285), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n302), .A4(new_n284), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n301), .A2(new_n304), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n303), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n302), .B1(new_n311), .B2(new_n284), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT13), .B(new_n283), .C1(new_n309), .C2(new_n310), .ZN(new_n321));
  OAI21_X1  g0121(.A(G169), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n270), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n304), .A2(new_n316), .A3(new_n313), .A4(G190), .ZN(new_n325));
  INV_X1    g0125(.A(new_n270), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n277), .A2(G226), .B1(new_n280), .B2(new_n281), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n289), .A2(G223), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G222), .A2(G1698), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n287), .B(new_n292), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n291), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n202), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n285), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT69), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n330), .A2(new_n338), .A3(new_n339), .A4(G190), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n330), .A2(new_n338), .A3(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT69), .ZN(new_n342));
  INV_X1    g0142(.A(G200), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n330), .B2(new_n338), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT10), .B1(new_n345), .B2(KEYINPUT68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G50), .B1(new_n207), .B2(G1), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n264), .A2(new_n349), .B1(G50), .B2(new_n263), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n250), .A2(G150), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT8), .B(G58), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n351), .B1(new_n201), .B2(new_n207), .C1(new_n352), .C2(new_n252), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n353), .B2(new_n256), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT67), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n348), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n256), .ZN(new_n359));
  INV_X1    g0159(.A(new_n350), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n355), .A3(new_n356), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n345), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n346), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n357), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n347), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n354), .A2(KEYINPUT67), .A3(KEYINPUT9), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n345), .C1(KEYINPUT68), .C2(KEYINPUT10), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n330), .A2(new_n338), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n271), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n361), .C1(G169), .C2(new_n372), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n264), .A2(new_n202), .A3(new_n265), .ZN(new_n375));
  INV_X1    g0175(.A(new_n263), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n202), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n207), .A2(new_n286), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n352), .A2(new_n378), .B1(new_n207), .B2(new_n202), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n252), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n256), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G232), .A2(G1698), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n289), .A2(G238), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n307), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n337), .C1(G107), .C2(new_n307), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n277), .A2(G244), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n282), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n384), .B(new_n391), .C1(new_n392), .C2(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n315), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n383), .C1(G179), .C2(new_n390), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n396), .A2(new_n364), .A3(new_n369), .A4(new_n374), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n329), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT75), .B1(new_n291), .B2(G33), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(new_n286), .A3(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n404), .A3(new_n292), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G20), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n307), .B2(G20), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n217), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT74), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G58), .A2(G68), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n207), .B1(new_n218), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n250), .A2(G159), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(G58), .A2(G68), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G58), .A2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n401), .B1(new_n410), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n419), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT74), .B1(new_n419), .B2(new_n414), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n307), .A2(new_n406), .A3(G20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n287), .A2(new_n292), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT7), .B1(new_n427), .B2(new_n207), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n429), .A3(KEYINPUT16), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n430), .A3(new_n256), .ZN(new_n431));
  INV_X1    g0231(.A(new_n264), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n352), .A2(new_n265), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n432), .A2(new_n433), .B1(new_n376), .B2(new_n352), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n274), .A2(new_n206), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G232), .A3(new_n285), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n282), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(G223), .A2(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n288), .A2(G1698), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n287), .A2(new_n440), .A3(new_n292), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G87), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n285), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n315), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n438), .A2(new_n444), .A3(new_n271), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n435), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT18), .ZN(new_n451));
  INV_X1    g0251(.A(new_n434), .ZN(new_n452));
  INV_X1    g0252(.A(new_n256), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n427), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n217), .B1(new_n409), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n421), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n456), .B2(KEYINPUT16), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n452), .B1(new_n457), .B2(new_n422), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n439), .A2(new_n445), .A3(new_n392), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n343), .B1(new_n438), .B2(new_n444), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n431), .A2(new_n461), .A3(KEYINPUT76), .A4(new_n434), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT17), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n435), .A2(new_n466), .A3(new_n449), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n451), .A2(new_n462), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT77), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n463), .B(KEYINPUT17), .ZN(new_n470));
  AOI211_X1 g0270(.A(KEYINPUT18), .B(new_n448), .C1(new_n431), .C2(new_n434), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n435), .B2(new_n449), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT77), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n400), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT78), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT78), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n400), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n206), .A2(G33), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n263), .A2(new_n483), .A3(new_n213), .A4(new_n255), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n376), .A2(KEYINPUT25), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT25), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n263), .B2(G107), .ZN(new_n489));
  AOI22_X1  g0289(.A1(G107), .A2(new_n485), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n287), .A2(new_n292), .A3(new_n207), .A4(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n307), .A2(new_n494), .A3(new_n207), .A4(G87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT84), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G116), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n286), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT23), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n207), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n486), .A2(KEYINPUT23), .A3(G20), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n501), .A2(new_n207), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n496), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n491), .B1(new_n510), .B2(new_n256), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT82), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(G41), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n272), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n273), .A2(G1), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(G41), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G264), .A3(new_n285), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n206), .A2(G45), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n513), .B2(G41), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(new_n280), .A3(new_n515), .A4(new_n514), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n228), .B2(G1698), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n307), .B1(G33), .B2(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n519), .B(new_n522), .C1(new_n525), .C2(new_n285), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n315), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n228), .A2(G1698), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G250), .B2(G1698), .ZN(new_n529));
  INV_X1    g0329(.A(G294), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n529), .A2(new_n427), .B1(new_n286), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n337), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n271), .A3(new_n522), .A4(new_n519), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n482), .B1(new_n511), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n496), .A2(new_n508), .A3(new_n505), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n508), .B1(new_n496), .B2(new_n505), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n256), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n490), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(KEYINPUT87), .A3(new_n533), .A4(new_n527), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n526), .A2(new_n343), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n532), .A2(new_n392), .A3(new_n522), .A4(new_n519), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(new_n543), .A3(new_n490), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n535), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G283), .ZN(new_n546));
  AND2_X1   g0346(.A1(G250), .A2(G1698), .ZN(new_n547));
  INV_X1    g0347(.A(G244), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n549), .B2(KEYINPUT4), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n546), .B1(new_n550), .B2(new_n427), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT4), .B1(new_n307), .B2(new_n549), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n337), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n554));
  INV_X1    g0354(.A(new_n546), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G250), .A2(G1698), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n555), .B1(new_n558), .B2(new_n307), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n289), .A2(G244), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n427), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n285), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT81), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n518), .A2(G257), .A3(new_n285), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n566), .A2(new_n522), .A3(new_n271), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n554), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n566), .A2(new_n522), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n553), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n315), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n378), .A2(new_n202), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n408), .A2(new_n409), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT79), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(KEYINPUT6), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n227), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(KEYINPUT6), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g0383(.A(G97), .B(G107), .Z(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g0385(.A(G97), .B(G107), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(G20), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n453), .B1(new_n574), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n376), .A2(new_n227), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n484), .B2(new_n227), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n568), .B(new_n571), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n589), .A2(new_n591), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n554), .A2(new_n565), .A3(new_n569), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n566), .A2(new_n522), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n563), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n599), .B2(G190), .ZN(new_n600));
  NOR4_X1   g0400(.A1(new_n598), .A2(new_n563), .A3(KEYINPUT83), .A4(new_n392), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n592), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n228), .A2(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n287), .A3(new_n292), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n307), .A2(KEYINPUT86), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n427), .A2(G303), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n287), .A2(new_n292), .A3(G264), .A4(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n337), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n518), .A2(G270), .A3(new_n285), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n522), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n498), .A2(new_n500), .A3(G20), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n546), .B(new_n207), .C1(G33), .C2(new_n227), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n256), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT20), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n616), .A2(KEYINPUT20), .A3(new_n256), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n498), .A2(new_n500), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n484), .A2(new_n497), .B1(new_n263), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n615), .A2(new_n626), .A3(G169), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n612), .A2(new_n614), .A3(G179), .ZN(new_n630));
  NAND2_X1  g0430(.A1(KEYINPUT21), .A2(G169), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n612), .B2(new_n614), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n626), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n499), .A2(G116), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n635));
  OAI21_X1  g0435(.A(G33), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n221), .A2(new_n289), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n548), .A2(G1698), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n287), .A2(new_n637), .A3(new_n292), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n285), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n516), .A2(new_n279), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n520), .A2(new_n223), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n285), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n315), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(G238), .A2(G1698), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n548), .B2(G1698), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n307), .B1(new_n623), .B2(G33), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n271), .B(new_n643), .C1(new_n648), .C2(new_n285), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n380), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n263), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n287), .A2(new_n292), .A3(new_n207), .A4(G68), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT19), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n207), .B1(new_n295), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n222), .A2(new_n227), .A3(new_n486), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT85), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n658), .B2(new_n654), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n653), .B(new_n657), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n652), .B1(new_n662), .B2(new_n256), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n484), .A2(new_n380), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n484), .A2(new_n222), .ZN(new_n667));
  AOI211_X1 g0467(.A(new_n652), .B(new_n667), .C1(new_n662), .C2(new_n256), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n343), .B1(new_n640), .B2(new_n644), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n392), .B(new_n643), .C1(new_n648), .C2(new_n285), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n650), .A2(new_n666), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n626), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n612), .A2(new_n614), .A3(G190), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n613), .A2(new_n522), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n337), .B2(new_n611), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n673), .B(new_n674), .C1(new_n676), .C2(new_n343), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n629), .A2(new_n633), .A3(new_n672), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n603), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n481), .A2(new_n545), .A3(new_n679), .ZN(G372));
  NAND2_X1  g0480(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n317), .A2(new_n318), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(new_n314), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT90), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n395), .B(new_n684), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n683), .A2(new_n270), .B1(new_n685), .B2(new_n328), .ZN(new_n686));
  INV_X1    g0486(.A(new_n470), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n473), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n370), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(new_n374), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  INV_X1    g0493(.A(new_n671), .ZN(new_n694));
  INV_X1    g0494(.A(new_n667), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n663), .A2(new_n695), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n652), .B(new_n664), .C1(new_n662), .C2(new_n256), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n645), .A2(new_n649), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n694), .A2(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n693), .B1(new_n592), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(G169), .B1(new_n569), .B2(new_n553), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n559), .A2(new_n562), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n564), .B1(new_n702), .B2(new_n337), .ZN(new_n703));
  AOI211_X1 g0503(.A(KEYINPUT81), .B(new_n285), .C1(new_n559), .C2(new_n562), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n701), .B1(new_n705), .B2(new_n567), .ZN(new_n706));
  INV_X1    g0506(.A(new_n572), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n427), .A2(new_n207), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n708), .A2(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n707), .B1(new_n709), .B2(new_n486), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n586), .B1(new_n579), .B2(new_n582), .ZN(new_n711));
  INV_X1    g0511(.A(new_n587), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n207), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n256), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n591), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n672), .A2(new_n706), .A3(KEYINPUT26), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n700), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n697), .A2(new_n698), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n692), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI211_X1 g0521(.A(KEYINPUT89), .B(new_n719), .C1(new_n700), .C2(new_n717), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT88), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n633), .A2(new_n629), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n534), .B1(new_n538), .B2(new_n490), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n544), .B(new_n672), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n727), .B2(new_n603), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n544), .A2(new_n672), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n612), .A2(new_n614), .A3(G179), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n676), .B2(new_n631), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n732));
  INV_X1    g0532(.A(new_n726), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n343), .B1(new_n705), .B2(new_n569), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n716), .ZN(new_n736));
  INV_X1    g0536(.A(new_n602), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(new_n716), .B2(new_n706), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n738), .A3(KEYINPUT88), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n728), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n723), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n691), .B1(new_n481), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT91), .ZN(G369));
  AOI21_X1  g0543(.A(KEYINPUT94), .B1(new_n732), .B2(new_n677), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT27), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n745), .B(KEYINPUT92), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT27), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n751), .A3(G213), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n748), .A2(new_n751), .A3(KEYINPUT93), .A4(G213), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G343), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n673), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n744), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n732), .A2(KEYINPUT94), .A3(new_n677), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n732), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G330), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n758), .A2(new_n539), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n535), .A2(new_n768), .A3(new_n540), .A4(new_n544), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n726), .A2(new_n758), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT95), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n733), .A2(new_n758), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n732), .A2(new_n758), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n779), .ZN(G399));
  INV_X1    g0580(.A(new_n210), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G41), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n656), .A2(G116), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(G1), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n219), .B2(new_n783), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n719), .B1(new_n700), .B2(new_n717), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n738), .A2(new_n544), .A3(new_n672), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n535), .A2(new_n540), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n725), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(KEYINPUT29), .A3(new_n759), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n758), .B1(new_n723), .B2(new_n740), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n794), .B2(KEYINPUT29), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n679), .A2(new_n545), .A3(new_n759), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT30), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n676), .A2(G179), .A3(new_n599), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n643), .B1(new_n648), .B2(new_n285), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n519), .B1(new_n525), .B2(new_n285), .ZN(new_n801));
  OAI21_X1  g0601(.A(KEYINPUT96), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n640), .A2(new_n644), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT96), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n803), .A2(new_n804), .A3(new_n519), .A4(new_n532), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n730), .A2(new_n570), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n808), .A2(KEYINPUT30), .A3(new_n805), .A4(new_n802), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n803), .A2(G179), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n594), .A2(new_n526), .A3(new_n615), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n807), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT31), .B1(new_n812), .B2(new_n758), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(KEYINPUT31), .A3(new_n758), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n797), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G330), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n796), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n787), .B1(new_n819), .B2(G1), .ZN(G364));
  INV_X1    g0620(.A(G13), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n206), .B1(new_n822), .B2(G45), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n782), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n767), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(G330), .B1(new_n763), .B2(new_n764), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OR3_X1    g0630(.A1(new_n830), .A2(KEYINPUT97), .A3(G20), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT97), .B1(new_n830), .B2(G20), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n765), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n825), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n213), .B1(G20), .B2(new_n315), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n210), .A2(G355), .A3(new_n307), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n781), .A2(new_n307), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(G45), .B2(new_n219), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n248), .A2(new_n273), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n840), .B1(G116), .B2(new_n210), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n835), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  INV_X1    g0646(.A(new_n836), .ZN(new_n847));
  NOR4_X1   g0647(.A1(new_n207), .A2(new_n392), .A3(new_n343), .A4(G179), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G87), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n207), .A2(new_n343), .A3(G179), .A4(G190), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G107), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n307), .A3(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT100), .Z(new_n853));
  NOR2_X1   g0653(.A1(G190), .A2(G200), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(G20), .A3(new_n271), .ZN(new_n855));
  INV_X1    g0655(.A(G159), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT32), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n207), .A2(new_n271), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n392), .A3(G200), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n854), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n862), .A2(G68), .B1(new_n864), .B2(G77), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(G190), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(G200), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n868), .A2(new_n216), .B1(new_n858), .B2(new_n857), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n343), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(G50), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n271), .A2(new_n343), .A3(G190), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(G20), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n871), .A2(new_n872), .B1(new_n227), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n853), .A2(new_n859), .A3(new_n865), .A4(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(G322), .ZN(new_n879));
  INV_X1    g0679(.A(G283), .ZN(new_n880));
  INV_X1    g0680(.A(new_n850), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n868), .A2(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G294), .B2(new_n874), .ZN(new_n883));
  XNOR2_X1  g0683(.A(KEYINPUT33), .B(G317), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n307), .B1(new_n862), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n855), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n864), .A2(G311), .B1(new_n886), .B2(G329), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n870), .A2(G326), .B1(G303), .B2(new_n848), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n883), .A2(new_n885), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n847), .B1(new_n878), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n846), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n826), .A2(new_n828), .B1(new_n834), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(G396));
  NAND2_X1  g0693(.A1(new_n396), .A2(new_n759), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n788), .B(new_n692), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n727), .A2(new_n724), .A3(new_n603), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT88), .B1(new_n734), .B2(new_n738), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n895), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n685), .A2(new_n383), .A3(new_n758), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n396), .B1(new_n384), .B2(new_n759), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n794), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n817), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT101), .Z(new_n906));
  AOI21_X1  g0706(.A(new_n825), .B1(new_n904), .B2(new_n817), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n836), .A2(new_n829), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n825), .B1(G77), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(G303), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n868), .A2(new_n530), .B1(new_n871), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(G107), .B2(new_n848), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n307), .B1(new_n862), .B2(G283), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n864), .A2(new_n623), .B1(new_n886), .B2(G311), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n881), .A2(new_n222), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(G97), .B2(new_n874), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n881), .A2(new_n217), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n427), .B(new_n920), .C1(G132), .C2(new_n886), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n848), .A2(G50), .B1(new_n874), .B2(G58), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n862), .A2(G150), .B1(new_n864), .B2(G159), .ZN(new_n923));
  INV_X1    g0723(.A(G143), .ZN(new_n924));
  INV_X1    g0724(.A(G137), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n923), .B1(new_n868), .B2(new_n924), .C1(new_n925), .C2(new_n871), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT34), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n921), .B(new_n922), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n919), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n911), .B1(new_n930), .B2(new_n836), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n903), .B2(new_n830), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n908), .A2(new_n932), .ZN(G384));
  NOR2_X1   g0733(.A1(new_n822), .A2(new_n206), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n431), .A2(new_n461), .A3(new_n434), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n421), .B2(new_n455), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n425), .A2(new_n429), .A3(KEYINPUT105), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n939), .A3(new_n401), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n452), .B1(new_n940), .B2(new_n457), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n936), .B1(new_n941), .B2(new_n756), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n448), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT37), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n435), .A2(new_n754), .A3(new_n755), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT37), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(new_n450), .A3(new_n946), .A4(new_n936), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(KEYINPUT106), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n941), .A2(new_n756), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n468), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT106), .B1(new_n944), .B2(new_n947), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n935), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n944), .A2(new_n947), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n956), .A2(KEYINPUT38), .A3(new_n950), .A4(new_n948), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n758), .A2(new_n270), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n324), .A2(new_n328), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n328), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n270), .B(new_n758), .C1(new_n683), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n816), .A2(new_n903), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT40), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n816), .A2(new_n903), .A3(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT109), .ZN(new_n969));
  INV_X1    g0769(.A(new_n945), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n468), .A2(KEYINPUT108), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n945), .A2(new_n936), .A3(new_n450), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT37), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n947), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT108), .B1(new_n468), .B2(new_n970), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n935), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n957), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT109), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n816), .A2(new_n979), .A3(new_n963), .A4(new_n903), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n969), .A2(new_n978), .A3(KEYINPUT40), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n967), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n481), .A2(new_n816), .ZN(new_n983));
  OAI21_X1  g0783(.A(G330), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n982), .B2(new_n983), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT110), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n963), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n758), .A2(new_n395), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT103), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n900), .A2(KEYINPUT104), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT104), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n894), .B1(new_n723), .B2(new_n740), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n990), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n988), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n958), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT39), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n978), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n683), .A2(new_n270), .A3(new_n759), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT107), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n953), .A2(KEYINPUT39), .A3(new_n957), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n756), .B1(new_n471), .B2(new_n472), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n997), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n796), .A2(new_n481), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n690), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1006), .B(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n934), .B1(new_n987), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n987), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n585), .A2(new_n587), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT35), .ZN(new_n1013));
  OAI211_X1 g0813(.A(G116), .B(new_n214), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT36), .Z(new_n1016));
  NOR3_X1   g0816(.A1(new_n219), .A2(new_n202), .A3(new_n417), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1017), .A2(KEYINPUT102), .B1(new_n872), .B2(G68), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT102), .B2(new_n1017), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(G1), .A3(new_n821), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1011), .A2(new_n1016), .A3(new_n1020), .ZN(G367));
  NOR2_X1   g0821(.A1(new_n759), .A2(new_n593), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1022), .A2(new_n603), .A3(KEYINPUT112), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT112), .B1(new_n1022), .B2(new_n603), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n758), .A2(new_n716), .A3(new_n706), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n774), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT95), .B1(new_n769), .B2(new_n770), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n778), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1028), .A2(KEYINPUT42), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n790), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n592), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n759), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT42), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n758), .A2(new_n696), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n672), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n720), .B2(new_n1038), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT43), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(KEYINPUT43), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n776), .A2(new_n1028), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1042), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n782), .B(KEYINPUT41), .Z(new_n1051));
  INV_X1    g0851(.A(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1031), .B1(new_n733), .B2(new_n758), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n779), .A2(KEYINPUT45), .A3(new_n1027), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(KEYINPUT44), .A3(new_n1028), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT44), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n779), .B2(new_n1027), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n776), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n775), .A2(new_n778), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n1031), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(new_n767), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1056), .A2(new_n1060), .A3(new_n776), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1063), .A2(new_n819), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1051), .B1(new_n1069), .B2(new_n819), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1049), .B(new_n1050), .C1(new_n1070), .C2(new_n824), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n837), .B1(new_n210), .B2(new_n380), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n841), .A2(new_n240), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n825), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n848), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n871), .A2(new_n924), .B1(new_n216), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G150), .B2(new_n867), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n863), .A2(new_n872), .B1(new_n855), .B2(new_n925), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n427), .B(new_n1078), .C1(G159), .C2(new_n862), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n874), .A2(G68), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n850), .A2(G77), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT46), .B1(new_n1075), .B2(new_n497), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n623), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT46), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1085), .B2(new_n1075), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n307), .B1(new_n862), .B2(G294), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n864), .A2(G283), .B1(new_n886), .B2(G317), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n850), .A2(G97), .B1(new_n874), .B2(G107), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G303), .A2(new_n867), .B1(new_n870), .B2(G311), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT113), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1082), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT47), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1074), .B1(new_n1094), .B2(new_n836), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n833), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n1040), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1071), .A2(new_n1097), .ZN(G387));
  NAND2_X1  g0898(.A1(new_n867), .A2(G317), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n912), .B2(new_n863), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT115), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT115), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G322), .A2(new_n870), .B1(new_n862), .B2(G311), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT48), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1075), .A2(new_n530), .B1(new_n880), .B2(new_n875), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n307), .B1(new_n886), .B2(G326), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n1084), .C2(new_n881), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT49), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n875), .A2(new_n380), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n202), .B2(new_n1075), .C1(new_n872), .C2(new_n868), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n307), .B1(new_n861), .B2(new_n352), .ZN(new_n1117));
  INV_X1    g0917(.A(G150), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n863), .A2(new_n217), .B1(new_n855), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n871), .A2(new_n856), .B1(new_n227), .B2(new_n881), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n836), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n784), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n210), .A3(new_n307), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(G107), .B2(new_n210), .ZN(new_n1125));
  AOI211_X1 g0925(.A(G45), .B(new_n1123), .C1(G68), .C2(G77), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n352), .A2(G50), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT50), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n781), .B(new_n307), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n237), .A2(G45), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1125), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT114), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(KEYINPUT114), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n839), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1122), .B(new_n825), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n775), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n833), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1067), .B2(new_n824), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1067), .A2(new_n819), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n782), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1067), .A2(new_n819), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(G393));
  NAND3_X1  g0942(.A1(new_n1063), .A2(new_n824), .A3(new_n1068), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n245), .A2(new_n841), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n837), .B1(new_n227), .B2(new_n210), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n825), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G150), .A2(new_n870), .B1(new_n867), .B2(G159), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT51), .Z(new_n1148));
  NOR2_X1   g0948(.A1(new_n875), .A2(new_n202), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1149), .B(new_n917), .C1(G68), .C2(new_n848), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n863), .A2(new_n352), .B1(new_n855), .B2(new_n924), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n427), .B(new_n1151), .C1(G50), .C2(new_n862), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G311), .A2(new_n867), .B1(new_n870), .B2(G317), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT52), .Z(new_n1155));
  OAI221_X1 g0955(.A(new_n851), .B1(new_n875), .B2(new_n1084), .C1(new_n1075), .C2(new_n880), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n427), .B1(new_n861), .B2(new_n912), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n863), .A2(new_n530), .B1(new_n855), .B2(new_n879), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1153), .A2(KEYINPUT116), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(KEYINPUT116), .B2(new_n1153), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1146), .B1(new_n1161), .B2(new_n836), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT117), .Z(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1096), .B2(new_n1027), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1143), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1068), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n776), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1139), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n1069), .A3(new_n782), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT118), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1168), .A2(new_n1069), .A3(new_n1171), .A4(new_n782), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1165), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(G390));
  NAND2_X1  g0974(.A1(new_n397), .A2(new_n399), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n329), .ZN(new_n1176));
  AND4_X1   g0976(.A1(new_n479), .A2(new_n1175), .A3(new_n1176), .A4(new_n476), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n479), .B1(new_n400), .B2(new_n476), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n818), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n690), .C1(new_n1180), .C2(new_n795), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT119), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1007), .A2(KEYINPUT119), .A3(new_n690), .A4(new_n1179), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n816), .A2(G330), .A3(new_n903), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n988), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n812), .A2(KEYINPUT31), .A3(new_n758), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1187), .A2(new_n813), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1188), .A2(new_n797), .B1(new_n901), .B2(new_n902), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(G330), .A3(new_n963), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT104), .B1(new_n900), .B2(new_n991), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n994), .A2(new_n993), .A3(new_n990), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n792), .A2(new_n759), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n989), .B1(new_n1195), .B2(new_n903), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n1186), .A3(new_n1190), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1183), .A2(new_n1184), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n999), .A2(new_n1003), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n996), .B2(new_n1002), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n978), .B(new_n1001), .C1(new_n1196), .C2(new_n988), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1201), .A2(new_n1190), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1190), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1183), .A2(new_n1184), .A3(new_n1198), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1190), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n963), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1208), .A2(new_n1001), .B1(new_n999), .B2(new_n1003), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1202), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1201), .A2(new_n1190), .A3(new_n1202), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1206), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1205), .A2(new_n1213), .A3(new_n782), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1200), .A2(new_n829), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT54), .B(G143), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n861), .A2(new_n925), .B1(new_n863), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT120), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n848), .A2(G150), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT53), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n427), .B1(new_n886), .B2(G125), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n856), .B2(new_n875), .C1(new_n872), .C2(new_n881), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1219), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G128), .A2(new_n870), .B1(new_n867), .B2(G132), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT121), .Z(new_n1226));
  OAI22_X1  g1026(.A1(new_n863), .A2(new_n227), .B1(new_n855), .B2(new_n530), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n307), .B(new_n1227), .C1(G107), .C2(new_n862), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1228), .B(new_n849), .C1(new_n217), .C2(new_n881), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1149), .B1(G116), .B2(new_n867), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n880), .B2(new_n871), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1224), .A2(new_n1226), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n836), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n835), .B1(new_n352), .B2(new_n909), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1216), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1215), .A2(new_n824), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1214), .A2(new_n1238), .ZN(G378));
  NAND2_X1  g1039(.A1(new_n370), .A2(new_n374), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n756), .A2(new_n354), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1240), .B(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1242), .B(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n980), .A2(KEYINPUT40), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n979), .B1(new_n1189), .B2(new_n963), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1248), .A2(new_n978), .B1(new_n966), .B2(new_n965), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1245), .B1(new_n1249), .B2(G330), .ZN(new_n1250));
  AND4_X1   g1050(.A1(G330), .A2(new_n967), .A3(new_n1245), .A4(new_n981), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1006), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1244), .B1(new_n982), .B2(new_n766), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n967), .A2(new_n1245), .A3(G330), .A4(new_n981), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n997), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1244), .A2(new_n829), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n825), .B1(G50), .B2(new_n910), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT123), .ZN(new_n1260));
  INV_X1    g1060(.A(G132), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n861), .A2(new_n1261), .B1(new_n863), .B2(new_n925), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n870), .A2(G125), .B1(G150), .B2(new_n874), .ZN(new_n1263));
  INV_X1    g1063(.A(G128), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n868), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1217), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1262), .B(new_n1265), .C1(new_n848), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT59), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n850), .A2(G159), .ZN(new_n1271));
  AOI211_X1 g1071(.A(G33), .B(G41), .C1(new_n886), .C2(G124), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n872), .B1(G33), .B2(G41), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n427), .B2(new_n272), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n871), .A2(new_n497), .B1(new_n216), .B2(new_n881), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G107), .B2(new_n867), .ZN(new_n1277));
  AOI211_X1 g1077(.A(G41), .B(new_n307), .C1(new_n862), .C2(G97), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n864), .A2(new_n651), .B1(new_n886), .B2(G283), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n848), .A2(G77), .B1(new_n874), .B2(G68), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT58), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1275), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1273), .B(new_n1283), .C1(new_n1282), .C2(new_n1281), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1260), .B1(new_n1284), .B2(new_n836), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1257), .A2(new_n824), .B1(new_n1258), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1215), .B2(new_n1198), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1250), .A2(new_n1006), .A3(new_n1251), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1253), .A2(new_n1255), .B1(new_n997), .B2(new_n1254), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT57), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n782), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1213), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT57), .B1(new_n1294), .B2(new_n1257), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1286), .B1(new_n1292), .B2(new_n1295), .ZN(G375));
  NAND2_X1  g1096(.A1(new_n988), .A2(new_n829), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n871), .A2(new_n530), .B1(new_n227), .B2(new_n1075), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(G283), .B2(new_n867), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1084), .A2(new_n861), .B1(new_n912), .B2(new_n855), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n307), .B(new_n1300), .C1(G107), .C2(new_n864), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1299), .A2(new_n1081), .A3(new_n1301), .A4(new_n1115), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n868), .A2(new_n925), .B1(new_n872), .B2(new_n875), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(G159), .B2(new_n848), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n863), .A2(new_n1118), .B1(new_n855), .B2(new_n1264), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n427), .B(new_n1305), .C1(new_n862), .C2(new_n1266), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n870), .A2(G132), .B1(G58), .B2(new_n850), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n847), .B1(new_n1302), .B2(new_n1308), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n835), .B(new_n1309), .C1(new_n217), .C2(new_n909), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1198), .A2(new_n824), .B1(new_n1297), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1206), .A2(new_n1051), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1198), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1312), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(G381));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G375), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(KEYINPUT124), .B(new_n1286), .C1(new_n1292), .C2(new_n1295), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1165), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1321), .A2(new_n1322), .A3(new_n1238), .A4(new_n1214), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n892), .B(new_n1138), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(G384), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1071), .A2(new_n1097), .A3(new_n1325), .A4(new_n1316), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1319), .A2(new_n1320), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1319), .A2(KEYINPUT125), .A3(new_n1327), .A4(new_n1320), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(G407));
  INV_X1    g1132(.A(G213), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(G378), .A2(G343), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1333), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G407), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(G407), .A2(new_n1336), .A3(KEYINPUT126), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G409));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  OAI211_X1 g1142(.A(G378), .B(new_n1286), .C1(new_n1292), .C2(new_n1295), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1294), .A2(new_n1257), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1286), .B1(new_n1344), .B2(new_n1051), .ZN(new_n1345));
  INV_X1    g1145(.A(G378), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  AOI22_X1  g1147(.A1(new_n1343), .A2(new_n1347), .B1(G213), .B2(new_n757), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1314), .B1(KEYINPUT60), .B2(new_n1199), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1198), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1287), .A2(KEYINPUT60), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n782), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1311), .B1(new_n1349), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(G384), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  OAI211_X1 g1155(.A(G384), .B(new_n1311), .C1(new_n1349), .C2(new_n1352), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n757), .A2(G213), .A3(G2897), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1355), .A2(new_n1356), .A3(new_n1358), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1342), .B1(new_n1348), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1357), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1348), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT63), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(G390), .A2(new_n1071), .A3(new_n1097), .ZN(new_n1369));
  OAI21_X1  g1169(.A(KEYINPUT127), .B1(G387), .B2(new_n1173), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(G387), .A2(new_n1173), .ZN(new_n1371));
  XNOR2_X1  g1171(.A(G393), .B(new_n892), .ZN(new_n1372));
  AND4_X1   g1172(.A1(new_n1369), .A2(new_n1370), .A3(new_n1371), .A4(new_n1372), .ZN(new_n1373));
  AOI22_X1  g1173(.A1(new_n1369), .A2(new_n1371), .B1(new_n1370), .B2(new_n1372), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1365), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1364), .A2(new_n1368), .A3(new_n1375), .A4(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT62), .ZN(new_n1378));
  AND3_X1   g1178(.A1(new_n1348), .A2(new_n1378), .A3(new_n1365), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1378), .B1(new_n1348), .B2(new_n1365), .ZN(new_n1380));
  NOR3_X1   g1180(.A1(new_n1379), .A2(new_n1363), .A3(new_n1380), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1377), .B1(new_n1381), .B2(new_n1375), .ZN(G405));
  NAND2_X1  g1182(.A1(G375), .A2(new_n1346), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1383), .A2(new_n1343), .ZN(new_n1384));
  XNOR2_X1  g1184(.A(new_n1384), .B(new_n1357), .ZN(new_n1385));
  XNOR2_X1  g1185(.A(new_n1385), .B(new_n1375), .ZN(G402));
endmodule


