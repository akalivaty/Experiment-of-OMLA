//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT65), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n217), .A2(G1), .A3(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(new_n207), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n202), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G107), .A2(G264), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n214), .B(new_n224), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT67), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G97), .B(G107), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(G264), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT86), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n257), .A2(KEYINPUT86), .A3(G264), .A4(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n252), .A2(new_n253), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G303), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(G257), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n256), .A2(new_n258), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n219), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT5), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n269), .B(G45), .C1(new_n270), .C2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT69), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT69), .A2(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT69), .A2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT69), .A2(G41), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT5), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n271), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n276), .A2(G270), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n266), .A2(new_n283), .A3(KEYINPUT87), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT87), .B1(new_n266), .B2(new_n283), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(G20), .B1(G33), .B2(G283), .ZN(new_n288));
  INV_X1    g0088(.A(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G97), .ZN(new_n290));
  INV_X1    g0090(.A(G116), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n290), .B1(G20), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n216), .A2(new_n218), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT20), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G116), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(G1), .B2(new_n289), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(new_n301), .B2(G116), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT88), .B1(new_n287), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G190), .B1(new_n284), .B2(new_n285), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n266), .A2(new_n283), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT87), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n266), .A2(new_n283), .A3(KEYINPUT87), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G200), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT88), .ZN(new_n311));
  INV_X1    g0111(.A(new_n303), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n304), .A2(new_n305), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n294), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G1), .B2(new_n221), .ZN(new_n316));
  MUX2_X1   g0116(.A(new_n298), .B(new_n316), .S(G77), .Z(new_n317));
  NAND2_X1  g0117(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT8), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G58), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G20), .A2(G33), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n322), .B1(G20), .B2(G77), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n221), .A2(G33), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n294), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n267), .A2(KEYINPUT70), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT70), .B1(new_n267), .B2(new_n330), .ZN(new_n332));
  OAI21_X1  g0132(.A(G244), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n273), .A2(new_n274), .A3(G45), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n281), .A2(G1), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n219), .A2(new_n264), .ZN(new_n340));
  OR2_X1    g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n261), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT66), .B(G238), .Z(new_n344));
  AOI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(G107), .B2(new_n259), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n257), .A2(G232), .A3(new_n261), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT77), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n346), .ZN(new_n349));
  OAI21_X1  g0149(.A(G1698), .B1(new_n252), .B2(new_n253), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n350), .A2(new_n225), .B1(new_n257), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n265), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT77), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n353), .A2(new_n354), .A3(new_n338), .A4(new_n333), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n355), .A3(G200), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n348), .B2(new_n355), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n329), .B(new_n356), .C1(new_n358), .C2(KEYINPUT78), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n348), .A2(new_n355), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n348), .A2(new_n355), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n366), .A3(new_n328), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT72), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n201), .A3(KEYINPUT8), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n298), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n316), .B2(new_n372), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n259), .B2(new_n221), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NOR4_X1   g0177(.A1(new_n252), .A2(new_n253), .A3(new_n377), .A4(G20), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n203), .A2(new_n205), .A3(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n322), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n315), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n375), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(G223), .B(new_n261), .C1(new_n252), .C2(new_n253), .ZN(new_n388));
  OAI211_X1 g0188(.A(G226), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n265), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n267), .A2(new_n330), .ZN(new_n393));
  INV_X1    g0193(.A(G45), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n277), .A2(new_n394), .A3(new_n278), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n393), .A2(G232), .B1(new_n395), .B2(new_n335), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n357), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n267), .A2(G232), .A3(new_n330), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n334), .B2(new_n336), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n265), .B2(new_n391), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n397), .B(KEYINPUT82), .C1(G200), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT82), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n402), .A3(new_n357), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n387), .A2(KEYINPUT17), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n377), .B1(new_n257), .B2(G20), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n202), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n381), .A2(G20), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n322), .A2(G159), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n384), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(new_n386), .A3(new_n294), .ZN(new_n412));
  INV_X1    g0212(.A(new_n375), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n401), .A2(new_n412), .A3(new_n413), .A4(new_n403), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n413), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT81), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT81), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n420), .A3(new_n413), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n400), .A2(G179), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n365), .B2(new_n400), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n417), .B1(KEYINPUT18), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n419), .A2(new_n426), .A3(new_n421), .A4(new_n423), .ZN(new_n427));
  OAI211_X1 g0227(.A(G232), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n428));
  OAI211_X1 g0228(.A(G226), .B(new_n261), .C1(new_n252), .C2(new_n253), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n265), .ZN(new_n432));
  OAI21_X1  g0232(.A(G238), .B1(new_n331), .B2(new_n332), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n338), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G190), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n433), .A3(new_n338), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT79), .A4(new_n338), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n316), .A2(new_n202), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n373), .A2(new_n202), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT12), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n443), .B(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT80), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n443), .B(KEYINPUT12), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n448), .C1(new_n202), .C2(new_n316), .ZN(new_n449));
  OR3_X1    g0249(.A1(new_n289), .A2(KEYINPUT73), .A3(G20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(G77), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n322), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n315), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n454), .A2(KEYINPUT11), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(KEYINPUT11), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n446), .A2(new_n449), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n286), .B1(new_n458), .B2(new_n435), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n441), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n435), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G169), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT14), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n464), .A3(G169), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n435), .A2(G179), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n439), .B2(new_n440), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n460), .B1(new_n469), .B2(new_n457), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n368), .A2(new_n425), .A3(new_n427), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n259), .A2(G1698), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(G222), .B1(G77), .B2(new_n259), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT71), .B(G223), .Z(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n350), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n265), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n267), .A2(new_n330), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n267), .A2(KEYINPUT70), .A3(new_n330), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G226), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n476), .A2(new_n482), .A3(new_n338), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G179), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n373), .A2(new_n207), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n316), .B2(new_n207), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n369), .A2(new_n450), .A3(new_n371), .A4(new_n451), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n322), .A2(G150), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(KEYINPUT74), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n208), .A2(G20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT74), .B1(new_n487), .B2(new_n488), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n294), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n493), .B2(KEYINPUT75), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT75), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n294), .C1(new_n491), .C2(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n483), .A2(new_n365), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n484), .B1(new_n499), .B2(KEYINPUT76), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT76), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT10), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(KEYINPUT9), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT9), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n494), .A2(new_n506), .A3(new_n496), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n483), .A2(G200), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n476), .A2(G190), .A3(new_n482), .A4(new_n338), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n504), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(KEYINPUT10), .B(new_n511), .C1(new_n505), .C2(new_n507), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n471), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n365), .B1(new_n297), .B2(new_n302), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n308), .A2(new_n517), .A3(new_n309), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n266), .A2(new_n283), .A3(G179), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n303), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n308), .A2(new_n517), .A3(KEYINPUT21), .A4(new_n309), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n301), .A2(G107), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n269), .A2(new_n351), .A3(G13), .A4(G20), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT25), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT89), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT89), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n294), .A2(new_n300), .A3(new_n351), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n527), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n289), .A2(new_n291), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n536), .A2(new_n221), .A3(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT23), .B1(new_n351), .B2(G20), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n535), .A2(G20), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n257), .A2(new_n221), .A3(G87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n257), .A2(new_n542), .A3(new_n221), .A4(G87), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n294), .B1(new_n544), .B2(KEYINPUT24), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT24), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n546), .B(new_n539), .C1(new_n541), .C2(new_n543), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n533), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G250), .A2(G1698), .ZN(new_n549));
  INV_X1    g0349(.A(G257), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G1698), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n257), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G294), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(new_n265), .B1(new_n276), .B2(G264), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n272), .A2(new_n275), .A3(G274), .A4(new_n267), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n363), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(new_n267), .C1(new_n279), .C2(new_n271), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n551), .A2(new_n257), .B1(G33), .B2(G294), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n556), .C1(new_n559), .C2(new_n340), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n365), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n548), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  AND4_X1   g0362(.A1(new_n520), .A2(new_n523), .A3(new_n524), .A4(new_n562), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n545), .A2(new_n547), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(new_n286), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n565), .B(KEYINPUT90), .C1(G190), .C2(new_n560), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT90), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n567), .A3(new_n286), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n564), .A2(new_n566), .A3(new_n533), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G244), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n252), .B2(new_n253), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G283), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n571), .B(KEYINPUT4), .C1(new_n253), .C2(new_n252), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n265), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n276), .A2(G257), .B1(new_n280), .B2(new_n282), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G190), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n322), .A2(G77), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  INV_X1    g0384(.A(G97), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n584), .A2(new_n585), .A3(G107), .ZN(new_n586));
  XNOR2_X1  g0386(.A(G97), .B(G107), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n588), .B2(new_n221), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n351), .B1(new_n405), .B2(new_n406), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n294), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n298), .A2(G97), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n301), .B2(G97), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n580), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n579), .A2(KEYINPUT83), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n578), .A2(new_n597), .A3(new_n265), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n582), .B(new_n594), .C1(new_n599), .C2(new_n286), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n394), .A2(G1), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n281), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n267), .C1(G250), .C2(new_n601), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G238), .A2(G1698), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n570), .B2(G1698), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n534), .B1(new_n605), .B2(new_n257), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(new_n340), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G200), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT84), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT84), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G87), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G97), .A2(G107), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n221), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n221), .B(G68), .C1(new_n252), .C2(new_n253), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n324), .B2(new_n585), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n294), .B1(new_n373), .B2(new_n325), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n301), .A2(G87), .ZN(new_n623));
  OAI211_X1 g0423(.A(G190), .B(new_n603), .C1(new_n606), .C2(new_n340), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n608), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n620), .ZN(new_n626));
  XNOR2_X1  g0426(.A(KEYINPUT84), .B(G87), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(new_n613), .B1(new_n221), .B2(new_n615), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n294), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n325), .A2(KEYINPUT85), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n325), .A2(KEYINPUT85), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n301), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n325), .A2(new_n373), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n607), .A2(new_n365), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n363), .B(new_n603), .C1(new_n606), .C2(new_n340), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n579), .A2(new_n580), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n365), .B1(new_n591), .B2(new_n593), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n578), .A2(new_n597), .A3(new_n265), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n597), .B1(new_n578), .B2(new_n265), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n363), .B(new_n580), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n569), .A2(new_n600), .A3(new_n638), .A4(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n314), .A2(new_n516), .A3(new_n563), .A4(new_n645), .ZN(G372));
  NAND4_X1  g0446(.A1(new_n569), .A2(new_n600), .A3(new_n638), .A4(new_n644), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n637), .B1(new_n563), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n640), .A2(new_n643), .A3(new_n637), .A4(new_n625), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT91), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n638), .A2(KEYINPUT26), .A3(new_n643), .A4(new_n640), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n654), .B2(KEYINPUT91), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n516), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n418), .A2(new_n423), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT18), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n418), .A2(new_n423), .A3(new_n426), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT92), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n367), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n460), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n364), .A2(KEYINPUT92), .A3(new_n366), .A4(new_n328), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n469), .A2(new_n457), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n660), .B1(new_n667), .B2(new_n417), .ZN(new_n668));
  INV_X1    g0468(.A(new_n507), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n506), .B1(new_n494), .B2(new_n496), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n512), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT10), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n508), .A2(new_n504), .A3(new_n512), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n668), .A2(new_n674), .B1(new_n502), .B2(new_n500), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n656), .A2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n269), .A2(new_n221), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n312), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n677), .A2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n314), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n548), .A2(new_n557), .A3(new_n561), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n548), .A2(new_n683), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n569), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n562), .A2(new_n683), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  INV_X1    g0497(.A(new_n694), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n677), .A2(new_n684), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n697), .B(new_n698), .C1(new_n699), .C2(new_n693), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n568), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n548), .A2(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n703), .A2(new_n566), .B1(new_n548), .B2(new_n683), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n677), .A2(new_n704), .A3(new_n562), .A4(new_n684), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n697), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n696), .B1(new_n701), .B2(new_n706), .ZN(G399));
  NOR2_X1   g0507(.A1(new_n614), .A2(G116), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT94), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n273), .A2(new_n274), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n212), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n709), .A2(new_n269), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n223), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  INV_X1    g0515(.A(new_n637), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n520), .A2(new_n523), .A3(new_n524), .A4(new_n562), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n645), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n683), .B1(new_n718), .B2(new_n654), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n684), .B1(new_n648), .B2(new_n655), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n580), .B1(new_n641), .B2(new_n642), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n560), .A2(new_n363), .A3(new_n607), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n308), .A3(new_n309), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n607), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n728), .A2(new_n555), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n522), .A2(new_n729), .A3(KEYINPUT30), .A4(new_n581), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n728), .A2(new_n555), .A3(new_n579), .A4(new_n580), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n521), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n683), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n563), .A2(new_n645), .A3(new_n314), .A4(new_n684), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n724), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n715), .B1(new_n745), .B2(G1), .ZN(G364));
  AND2_X1   g0546(.A1(new_n221), .A2(G13), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n269), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n712), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n212), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n259), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G355), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G116), .B2(new_n212), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n247), .A2(new_n394), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n751), .A2(new_n257), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n223), .B2(new_n394), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n220), .B1(G20), .B2(new_n365), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n750), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n363), .A2(new_n357), .A3(G20), .A4(G200), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n363), .A2(new_n286), .A3(KEYINPUT97), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT97), .B1(new_n363), .B2(new_n286), .ZN(new_n773));
  OAI211_X1 g0573(.A(G20), .B(new_n357), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n771), .A2(G283), .B1(new_n775), .B2(G329), .ZN(new_n776));
  NAND2_X1  g0576(.A1(G20), .A2(G179), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n286), .A3(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT33), .B(G317), .Z(new_n780));
  NOR3_X1   g0580(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n777), .A2(new_n357), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n357), .A2(new_n286), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(G20), .A3(G179), .ZN(new_n789));
  INV_X1    g0589(.A(G326), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n786), .A2(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n788), .A2(G20), .A3(new_n363), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n259), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n784), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n772), .A2(new_n773), .ZN(new_n797));
  OAI21_X1  g0597(.A(G20), .B1(new_n797), .B2(new_n357), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n776), .B(new_n795), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n799), .A2(new_n585), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n774), .A2(KEYINPUT32), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n257), .B1(new_n792), .B2(new_n627), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n779), .A2(new_n202), .B1(new_n789), .B2(new_n207), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G58), .C2(new_n785), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n781), .A2(KEYINPUT96), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n781), .A2(KEYINPUT96), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n812), .A2(G77), .B1(new_n771), .B2(G107), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n774), .B2(new_n803), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n805), .A2(new_n808), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT100), .B1(new_n801), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n760), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n801), .A2(KEYINPUT100), .A3(new_n815), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n766), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n763), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n689), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT101), .Z(new_n823));
  NOR2_X1   g0623(.A1(new_n689), .A2(G330), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n824), .B(new_n690), .C1(new_n711), .C2(new_n748), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n823), .A2(new_n825), .ZN(G396));
  NOR2_X1   g0626(.A1(new_n760), .A2(new_n761), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT102), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n771), .A2(G87), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n291), .B2(new_n811), .C1(new_n783), .C2(new_n774), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n259), .B1(new_n786), .B2(new_n796), .ZN(new_n831));
  INV_X1    g0631(.A(new_n789), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G303), .B1(G283), .B2(new_n778), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n351), .B2(new_n792), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n830), .A2(new_n802), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n771), .A2(G68), .ZN(new_n836));
  INV_X1    g0636(.A(new_n792), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n259), .B1(new_n837), .B2(G50), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n838), .C1(new_n839), .C2(new_n774), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G58), .B2(new_n798), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n832), .A2(G137), .B1(G150), .B2(new_n778), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n786), .C1(new_n811), .C2(new_n803), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n835), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n750), .B1(G77), .B2(new_n828), .C1(new_n846), .C2(new_n817), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT103), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n329), .A2(new_n684), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n662), .A2(new_n664), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n849), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n367), .B(new_n851), .C1(new_n359), .C2(new_n360), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n848), .B1(new_n762), .B2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT104), .Z(new_n855));
  OAI211_X1 g0655(.A(new_n684), .B(new_n853), .C1(new_n648), .C2(new_n655), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT105), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n850), .A2(KEYINPUT105), .A3(new_n852), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n861));
  INV_X1    g0661(.A(new_n651), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n683), .B1(new_n863), .B2(new_n718), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n856), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(new_n743), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n750), .B1(new_n865), .B2(new_n743), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n855), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G384));
  INV_X1    g0670(.A(new_n588), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(KEYINPUT35), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(KEYINPUT35), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(G116), .A3(new_n222), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT106), .B(KEYINPUT36), .Z(new_n875));
  XNOR2_X1  g0675(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n223), .A2(G77), .A3(new_n380), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n207), .A2(G68), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n269), .B(G13), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(G330), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n404), .A2(new_n416), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n424), .A2(KEYINPUT18), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n427), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n387), .A2(new_n681), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT107), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n414), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n681), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n419), .A2(new_n421), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n424), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n657), .A2(new_n414), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n893), .B2(new_n885), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT38), .A4(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AOI221_X4 g0697(.A(new_n897), .B1(new_n892), .B2(new_n894), .C1(new_n884), .C2(new_n885), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n412), .A2(new_n420), .A3(new_n413), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n420), .B1(new_n412), .B2(new_n413), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n899), .A2(new_n900), .A3(new_n681), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n901), .B2(new_n893), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n658), .A2(new_n404), .A3(new_n416), .A4(new_n659), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n902), .A2(new_n892), .B1(new_n903), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT107), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n896), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n736), .A2(new_n735), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n739), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n457), .A2(new_n683), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n464), .B1(new_n461), .B2(G169), .ZN(new_n910));
  AOI211_X1 g0710(.A(KEYINPUT14), .B(new_n365), .C1(new_n458), .C2(new_n435), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n910), .A2(new_n911), .A3(new_n467), .ZN(new_n912));
  INV_X1    g0712(.A(new_n457), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n663), .B(new_n909), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n457), .B(new_n683), .C1(new_n469), .C2(new_n460), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(new_n850), .B2(new_n852), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n916), .A3(KEYINPUT40), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n906), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n886), .B2(new_n895), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n908), .B(new_n916), .C1(new_n898), .C2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n516), .A2(new_n908), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n881), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n896), .C1(new_n898), .C2(new_n905), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n666), .A2(new_n683), .ZN(new_n928));
  INV_X1    g0728(.A(new_n885), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n425), .B2(new_n427), .ZN(new_n930));
  INV_X1    g0730(.A(new_n895), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n897), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(new_n928), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n660), .A2(new_n890), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n914), .A2(new_n915), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n367), .A2(new_n683), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n856), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n936), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n935), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n516), .A2(new_n723), .A3(new_n720), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n675), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n925), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n269), .B2(new_n747), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n925), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n880), .B1(new_n949), .B2(new_n950), .ZN(G367));
  OAI211_X1 g0751(.A(new_n600), .B(new_n644), .C1(new_n594), .C2(new_n684), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n640), .A2(new_n643), .A3(new_n683), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n705), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n691), .A2(new_n600), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n683), .B1(new_n958), .B2(new_n644), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n956), .B2(KEYINPUT42), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n622), .A2(new_n623), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n683), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n638), .A2(new_n962), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n963), .A2(KEYINPUT108), .B1(new_n637), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(KEYINPUT108), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n957), .A2(new_n960), .B1(KEYINPUT43), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n967), .B(new_n968), .Z(new_n969));
  NOR2_X1   g0769(.A1(new_n696), .A2(new_n955), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n711), .B(KEYINPUT41), .ZN(new_n972));
  XNOR2_X1  g0772(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n701), .A2(new_n706), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n955), .ZN(new_n976));
  NOR4_X1   g0776(.A1(new_n701), .A2(new_n706), .A3(KEYINPUT110), .A4(new_n954), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n954), .B1(new_n701), .B2(new_n706), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n706), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(new_n700), .A3(new_n955), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n975), .A2(new_n974), .A3(new_n955), .ZN(new_n985));
  INV_X1    g0785(.A(new_n973), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n978), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n696), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n695), .B(new_n699), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n690), .B(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n744), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n978), .A2(new_n981), .A3(new_n696), .A4(new_n987), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n972), .B1(new_n995), .B2(new_n745), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n971), .B1(new_n996), .B2(new_n749), .ZN(new_n997));
  INV_X1    g0797(.A(new_n750), .ZN(new_n998));
  INV_X1    g0798(.A(new_n325), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n765), .B1(new_n751), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n242), .A2(new_n756), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n257), .B1(new_n779), .B2(new_n803), .ZN(new_n1003));
  INV_X1    g0803(.A(G150), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n786), .A2(new_n1004), .B1(new_n792), .B2(new_n201), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G143), .C2(new_n832), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n799), .A2(new_n202), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n771), .A2(G77), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n812), .A2(G50), .B1(G137), .B2(new_n775), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n837), .A2(G116), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT46), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1012), .A2(new_n1013), .B1(G294), .B2(new_n778), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT111), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(KEYINPUT111), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n259), .B1(new_n789), .B2(new_n783), .C1(new_n793), .C2(new_n786), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n770), .A2(new_n585), .B1(new_n1021), .B2(new_n774), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(G283), .C2(new_n812), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1019), .B(new_n1023), .C1(new_n351), .C2(new_n799), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1011), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT47), .Z(new_n1027));
  OAI221_X1 g0827(.A(new_n1002), .B1(new_n821), .B2(new_n966), .C1(new_n1027), .C2(new_n817), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n997), .A2(new_n1029), .ZN(G387));
  AOI22_X1  g0830(.A1(new_n832), .A2(G322), .B1(G311), .B2(new_n778), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n1021), .B2(new_n786), .C1(new_n811), .C2(new_n793), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n798), .A2(G283), .B1(G294), .B2(new_n837), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT49), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n259), .B1(new_n774), .B2(new_n790), .C1(new_n770), .C2(new_n291), .ZN(new_n1041));
  OR3_X1    g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n257), .B1(new_n782), .B2(new_n202), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n786), .A2(new_n207), .B1(new_n789), .B2(new_n803), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G77), .C2(new_n837), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n775), .A2(G150), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n372), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n771), .A2(G97), .B1(new_n1047), .B2(new_n778), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n798), .A2(new_n630), .A3(new_n631), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n817), .B1(new_n1042), .B2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n239), .A2(new_n394), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1052), .A2(new_n756), .B1(new_n709), .B2(new_n752), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n321), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT50), .B1(new_n1054), .B2(G50), .ZN(new_n1055));
  INV_X1    g0855(.A(G77), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n394), .C1(new_n202), .C2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1054), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n709), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1053), .A2(new_n1059), .B1(G107), .B2(new_n212), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n998), .B(new_n1051), .C1(new_n764), .C2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n763), .B1(new_n693), .B2(new_n694), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n712), .B1(new_n992), .B2(new_n744), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n992), .A2(new_n744), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1063), .B1(new_n748), .B2(new_n992), .C1(new_n1064), .C2(new_n1065), .ZN(G393));
  AND2_X1   g0866(.A1(new_n995), .A2(new_n712), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n990), .A2(new_n994), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n993), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n250), .A2(new_n757), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n764), .B1(new_n585), .B2(new_n212), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n832), .A2(G317), .B1(G311), .B2(new_n785), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  INV_X1    g0873(.A(G283), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n782), .A2(new_n796), .B1(new_n792), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n257), .B(new_n1075), .C1(G303), .C2(new_n778), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n351), .B2(new_n770), .C1(new_n787), .C2(new_n774), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(G116), .C2(new_n798), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n832), .A2(G150), .B1(G159), .B2(new_n785), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n259), .B1(new_n837), .B2(G68), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n829), .B(new_n1081), .C1(new_n843), .C2(new_n774), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(G77), .C2(new_n798), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n811), .A2(new_n1054), .B1(new_n207), .B2(new_n779), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n1078), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n750), .B1(new_n1070), .B2(new_n1071), .C1(new_n1086), .C2(new_n817), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n763), .B2(new_n955), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1068), .B2(new_n749), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1069), .A2(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(KEYINPUT115), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n928), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n940), .B1(new_n864), .B2(new_n853), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1092), .C1(new_n1093), .C2(new_n939), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n927), .A2(new_n934), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT115), .B1(new_n942), .B2(new_n928), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n906), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n940), .B1(new_n719), .B2(new_n853), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1092), .C1(new_n939), .C2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n742), .A2(G330), .A3(new_n853), .A4(new_n938), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n881), .B1(new_n739), .B2(new_n907), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n916), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n742), .A2(G330), .A3(new_n853), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1107), .A2(new_n939), .B1(new_n916), .B2(new_n1104), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n938), .B1(new_n860), .B2(new_n1104), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1108), .A2(new_n1093), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n516), .A2(new_n1104), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n945), .A2(new_n675), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT116), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT116), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1106), .A2(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1105), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT116), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(new_n1127), .A3(new_n712), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n786), .A2(new_n839), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n259), .B(new_n1129), .C1(G128), .C2(new_n832), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n771), .A2(G50), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n792), .A2(new_n1004), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n775), .A2(G125), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G159), .B2(new_n798), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  INV_X1    g0937(.A(G137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n811), .A2(new_n1137), .B1(new_n1138), .B2(new_n779), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT117), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n798), .A2(G77), .B1(G116), .B2(new_n785), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT118), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n812), .A2(G97), .B1(G294), .B2(new_n775), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n257), .B1(new_n837), .B2(G87), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n832), .A2(G283), .B1(G107), .B2(new_n778), .ZN(new_n1145));
  AND4_X1   g0945(.A1(new_n836), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1136), .A2(new_n1140), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n750), .B1(new_n1047), .B2(new_n828), .C1(new_n1147), .C2(new_n817), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1095), .B2(new_n761), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT119), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1121), .A2(new_n749), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1128), .A2(new_n1150), .A3(new_n1151), .ZN(G378));
  INV_X1    g0952(.A(new_n944), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n908), .A2(new_n916), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n933), .B2(new_n932), .ZN(new_n1155));
  OAI21_X1  g0955(.A(G330), .B1(new_n1155), .B2(KEYINPUT40), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n497), .A2(new_n890), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n515), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n674), .A2(new_n503), .A3(new_n1157), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1156), .A2(new_n1166), .A3(new_n918), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n881), .B1(new_n921), .B2(new_n919), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n917), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n896), .C1(new_n898), .C2(new_n905), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1170), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1153), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT123), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1166), .B1(new_n1156), .B2(new_n918), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1171), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n944), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT123), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1177), .A2(new_n944), .A3(new_n1178), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1176), .A2(new_n1181), .A3(KEYINPUT122), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT122), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1180), .B1(new_n1185), .B2(new_n1153), .ZN(new_n1186));
  AOI211_X1 g0986(.A(KEYINPUT123), .B(new_n944), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1114), .B1(new_n1106), .B2(new_n1117), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT57), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1113), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1182), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1179), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n712), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1183), .A2(new_n1188), .A3(new_n749), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n771), .A2(G58), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n630), .A2(new_n631), .A3(new_n781), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n1074), .C2(new_n774), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n259), .B(new_n710), .C1(new_n792), .C2(new_n1056), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n832), .A2(G116), .B1(G107), .B2(new_n785), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n585), .B2(new_n779), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1202), .A2(new_n1007), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G33), .A2(G41), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT120), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n710), .A2(new_n259), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n207), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1207), .A2(new_n1208), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n832), .A2(G125), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n1138), .B2(new_n782), .C1(new_n792), .C2(new_n1137), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G128), .A2(new_n785), .B1(new_n778), .B2(G132), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n1004), .C2(new_n799), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1210), .B1(new_n775), .B2(G124), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n803), .B2(new_n770), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n760), .B1(new_n1213), .B2(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT121), .Z(new_n1225));
  AOI211_X1 g1025(.A(new_n998), .B(new_n1225), .C1(new_n207), .C2(new_n827), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1170), .A2(new_n761), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1199), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1198), .A2(new_n1230), .ZN(G375));
  NAND2_X1  g1031(.A1(new_n1111), .A2(new_n749), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n750), .B1(new_n828), .B2(G68), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n782), .A2(new_n1004), .B1(new_n792), .B2(new_n803), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n779), .A2(new_n1137), .B1(new_n789), .B2(new_n839), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n257), .B1(new_n786), .B2(new_n1138), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n798), .A2(G50), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n775), .A2(G128), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1237), .A2(new_n1200), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1049), .B1(new_n1074), .B2(new_n786), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT124), .Z(new_n1242));
  AOI22_X1  g1042(.A1(new_n812), .A2(G107), .B1(G303), .B2(new_n775), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n257), .B1(new_n837), .B2(G97), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n832), .A2(G294), .B1(G116), .B2(new_n778), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1009), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1233), .B1(new_n1247), .B2(new_n760), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n938), .B2(new_n762), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1232), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n972), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1251), .B1(new_n1255), .B2(new_n1126), .ZN(G381));
  NOR2_X1   g1056(.A1(G375), .A2(G378), .ZN(new_n1257));
  OR3_X1    g1057(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(G407));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n682), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(G213), .ZN(G409));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G343), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1253), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n711), .B1(new_n1252), .B2(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1270), .B2(new_n1251), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1269), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1267), .B2(new_n1253), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1273), .A2(new_n869), .A3(new_n1250), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1266), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1270), .A2(G384), .A3(new_n1251), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n869), .B1(new_n1273), .B2(new_n1250), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1265), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1198), .A2(G378), .A3(new_n1230), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1183), .A2(new_n1188), .A3(new_n1189), .A4(new_n1254), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n748), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1227), .B2(new_n1226), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G378), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1280), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1264), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1279), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1196), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1128), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1229), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1287), .B(new_n1290), .C1(new_n1293), .C2(new_n1284), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1288), .A2(KEYINPUT125), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(G387), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n997), .B2(new_n1029), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1296), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1298), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT126), .B1(new_n997), .B2(new_n1029), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1303), .B(G390), .C1(new_n1304), .C2(new_n1298), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1229), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1284), .B1(new_n1310), .B2(G378), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1311), .B2(new_n1264), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1308), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1294), .A2(new_n1289), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1295), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1286), .A2(new_n1318), .A3(new_n1287), .A4(new_n1290), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1317), .A2(new_n1312), .A3(new_n1319), .A4(new_n1307), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1306), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1316), .A2(new_n1322), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1292), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1290), .A2(new_n1325), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1324), .A2(new_n1280), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1326), .B1(new_n1324), .B2(new_n1280), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1306), .ZN(G402));
endmodule


