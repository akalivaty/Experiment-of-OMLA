//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(new_n217), .B2(new_n216), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AND3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n212), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n219), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(G232), .Z(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  OAI21_X1  g0044(.A(KEYINPUT68), .B1(new_n211), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT68), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n247), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT67), .B(G1), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n249), .B1(G20), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n257), .A2(new_n259), .A3(G13), .A4(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n253), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT75), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n266));
  AOI21_X1  g0066(.A(G20), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n263), .B1(new_n267), .B2(KEYINPUT7), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(KEYINPUT75), .B(new_n269), .C1(new_n270), .C2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT74), .B(G33), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n266), .B1(new_n273), .B2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G20), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G68), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G58), .A2(G68), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n280), .A2(G20), .B1(G159), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT16), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n244), .A2(KEYINPUT74), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT74), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT3), .ZN(new_n287));
  AOI21_X1  g0087(.A(G20), .B1(new_n287), .B2(new_n265), .ZN(new_n288));
  OAI21_X1  g0088(.A(G68), .B1(new_n288), .B2(new_n269), .ZN(new_n289));
  INV_X1    g0089(.A(new_n265), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n273), .B2(KEYINPUT3), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(KEYINPUT7), .A3(G20), .ZN(new_n292));
  OAI211_X1 g0092(.A(KEYINPUT16), .B(new_n282), .C1(new_n289), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n249), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n262), .B1(new_n283), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n208), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G226), .A2(G1698), .ZN(new_n298));
  INV_X1    g0098(.A(G223), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(G1698), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n287), .A2(new_n265), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G87), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n257), .A2(new_n259), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G41), .A2(G45), .ZN(new_n305));
  OAI211_X1 g0105(.A(G232), .B(new_n297), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n208), .B2(new_n296), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT66), .B1(new_n305), .B2(G1), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT66), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n256), .C1(G41), .C2(G45), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n314), .A2(KEYINPUT76), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT76), .B1(new_n314), .B2(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n315), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n295), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT18), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n295), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR4_X1   g0124(.A1(new_n303), .A2(new_n313), .A3(KEYINPUT77), .A4(G190), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT77), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n314), .B2(G200), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OR3_X1    g0130(.A1(new_n295), .A2(KEYINPUT17), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT78), .B1(new_n295), .B2(new_n330), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n329), .ZN(new_n333));
  INV_X1    g0133(.A(new_n325), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT78), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n272), .B2(new_n276), .ZN(new_n339));
  INV_X1    g0139(.A(new_n282), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(new_n293), .A3(new_n249), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n335), .A2(new_n336), .A3(new_n342), .A4(new_n262), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n332), .A2(KEYINPUT17), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n324), .B1(new_n331), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n312), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n304), .A2(new_n305), .ZN(new_n347));
  INV_X1    g0147(.A(new_n297), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(G226), .ZN(new_n350));
  INV_X1    g0150(.A(G1698), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n270), .A2(G222), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n270), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n270), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n299), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n348), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G169), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n315), .B2(new_n358), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n275), .A2(G33), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n253), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n275), .B1(new_n201), .B2(new_n202), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT69), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n281), .A2(G150), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n363), .A2(KEYINPUT69), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n249), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n260), .A2(G50), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n251), .B2(G50), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G20), .A2(G77), .ZN(new_n373));
  INV_X1    g0173(.A(new_n281), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  OAI221_X1 g0175(.A(new_n373), .B1(new_n253), .B2(new_n374), .C1(new_n361), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n249), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n251), .A2(G77), .ZN(new_n378));
  INV_X1    g0178(.A(new_n260), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n353), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n270), .A2(G232), .A3(new_n351), .ZN(new_n383));
  INV_X1    g0183(.A(G107), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n383), .B1(new_n384), .B2(new_n270), .C1(new_n355), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n348), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n346), .B1(new_n349), .B2(G244), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G169), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(G179), .A3(new_n388), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n382), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n389), .A2(G190), .ZN(new_n394));
  AOI21_X1  g0194(.A(G200), .B1(new_n387), .B2(new_n388), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n382), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT71), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n358), .B2(G200), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT9), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n371), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n350), .A2(new_n357), .A3(G190), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT10), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT9), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT70), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n406), .B(KEYINPUT70), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT10), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n372), .B(new_n397), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n379), .A2(new_n338), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT12), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT11), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n374), .A2(new_n202), .B1(new_n275), .B2(G68), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n361), .A2(new_n353), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n249), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n414), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n415), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n252), .B2(new_n338), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n312), .A2(KEYINPUT73), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT73), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n308), .A2(new_n309), .A3(new_n426), .A4(new_n311), .ZN(new_n427));
  OAI211_X1 g0227(.A(G238), .B(new_n297), .C1(new_n304), .C2(new_n305), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G97), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n265), .A2(new_n266), .A3(G226), .A4(new_n351), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT72), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n270), .A2(new_n435), .A3(G226), .A4(new_n351), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n424), .B(new_n429), .C1(new_n438), .C2(new_n297), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n297), .B1(new_n432), .B2(new_n437), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT13), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(G179), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G169), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n439), .B2(new_n442), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT14), .B(new_n444), .C1(new_n439), .C2(new_n442), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n423), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n439), .A2(new_n328), .A3(new_n442), .ZN(new_n450));
  AOI21_X1  g0250(.A(G200), .B1(new_n439), .B2(new_n442), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n422), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n345), .A2(new_n412), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT79), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n345), .A2(new_n412), .A3(new_n457), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n291), .A2(new_n275), .A3(G68), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n275), .B1(new_n431), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(G87), .A2(G97), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n384), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n275), .A2(G33), .A3(G97), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n464), .A2(new_n466), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n461), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n375), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n260), .ZN(new_n471));
  AND3_X1   g0271(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n208), .B1(new_n472), .B2(new_n247), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n257), .A2(new_n259), .A3(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n260), .A3(new_n245), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G87), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n469), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n287), .A2(G244), .A3(G1698), .A4(new_n265), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n385), .A2(G1698), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n287), .A2(new_n265), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n284), .A2(new_n286), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G116), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n348), .ZN(new_n485));
  INV_X1    g0285(.A(new_n296), .ZN(new_n486));
  OAI21_X1  g0286(.A(G274), .B1(new_n486), .B2(new_n246), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n257), .A2(new_n259), .A3(G45), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT82), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n308), .A2(new_n490), .A3(new_n250), .A4(G45), .ZN(new_n491));
  INV_X1    g0291(.A(G250), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n348), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n489), .A2(new_n491), .B1(new_n493), .B2(new_n488), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n485), .A2(G190), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n485), .A2(new_n494), .ZN(new_n496));
  INV_X1    g0296(.A(G200), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n478), .B(new_n495), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n469), .ZN(new_n500));
  INV_X1    g0300(.A(new_n475), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n470), .ZN(new_n502));
  INV_X1    g0302(.A(new_n471), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n485), .A2(G179), .A3(new_n494), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n444), .B1(new_n485), .B2(new_n494), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT83), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT83), .B1(new_n505), .B2(new_n506), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n461), .A2(G116), .A3(new_n260), .A4(new_n474), .ZN(new_n512));
  INV_X1    g0312(.A(G116), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n379), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G33), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n275), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n275), .A2(new_n513), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n521), .A2(KEYINPUT20), .A3(new_n249), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT20), .B1(new_n521), .B2(new_n249), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n512), .B(new_n514), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G270), .B(new_n297), .C1(new_n488), .C2(new_n527), .ZN(new_n528));
  XNOR2_X1  g0328(.A(KEYINPUT5), .B(G41), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n308), .A2(new_n250), .A3(new_n529), .A4(G45), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G264), .A2(G1698), .ZN(new_n533));
  INV_X1    g0333(.A(G257), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n287), .A2(new_n265), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n265), .A2(new_n266), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G303), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n348), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n524), .A2(KEYINPUT21), .A3(G169), .A4(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n514), .B1(new_n475), .B2(new_n513), .ZN(new_n544));
  INV_X1    g0344(.A(new_n523), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n521), .A2(KEYINPUT20), .A3(new_n249), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n297), .B1(new_n536), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g0348(.A(G169), .B1(new_n548), .B2(new_n531), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n543), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n548), .A2(new_n531), .A3(new_n315), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n524), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n524), .B2(new_n551), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n542), .B(new_n550), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n541), .A2(new_n497), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n548), .A2(new_n531), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n328), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n547), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT81), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n297), .C1(new_n488), .C2(new_n527), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n564), .A2(new_n530), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n265), .A2(new_n266), .A3(G250), .A4(G1698), .ZN(new_n566));
  AND2_X1   g0366(.A1(KEYINPUT4), .A2(G244), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n265), .A2(new_n266), .A3(new_n567), .A4(new_n351), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n568), .A3(new_n515), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n287), .A2(G244), .A3(new_n351), .A4(new_n265), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n565), .B1(new_n572), .B2(new_n297), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n563), .B1(new_n573), .B2(G179), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n571), .A2(new_n570), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n348), .B1(new_n575), .B2(new_n569), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(KEYINPUT81), .A3(new_n315), .A4(new_n565), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n384), .B1(new_n272), .B2(new_n276), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  AND2_X1   g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G97), .A2(G107), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n384), .A2(KEYINPUT6), .A3(G97), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n275), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n374), .A2(new_n353), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT80), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  INV_X1    g0388(.A(new_n586), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT6), .A2(G97), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(G107), .ZN(new_n591));
  XNOR2_X1  g0391(.A(G97), .B(G107), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n580), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n588), .B(new_n589), .C1(new_n593), .C2(new_n275), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n249), .B1(new_n579), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n260), .A2(new_n516), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n501), .B2(new_n516), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n596), .A2(new_n598), .B1(new_n444), .B2(new_n573), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n596), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n573), .A2(new_n497), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(G190), .B2(new_n573), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n578), .A2(new_n599), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G264), .B(new_n297), .C1(new_n488), .C2(new_n527), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n530), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G257), .A2(G1698), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n492), .B2(G1698), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n287), .A2(new_n265), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n482), .A2(G294), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n297), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(KEYINPUT85), .B2(new_n610), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n328), .ZN(new_n613));
  INV_X1    g0413(.A(new_n610), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n530), .A3(new_n604), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n497), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT22), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n476), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n287), .A2(new_n275), .A3(new_n265), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n275), .A2(G87), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n537), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT23), .B1(new_n275), .B2(G107), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT23), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n384), .A3(G20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n482), .A2(new_n275), .A3(G116), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n620), .A2(new_n622), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT24), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n273), .A2(new_n513), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n626), .B1(new_n632), .B2(new_n275), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(KEYINPUT24), .A3(new_n620), .A4(new_n622), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n634), .A3(new_n249), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n475), .A2(new_n384), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT25), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n379), .B2(new_n384), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n260), .A2(KEYINPUT25), .A3(G107), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n617), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n640), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n444), .B1(new_n611), .B2(new_n612), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n615), .A2(new_n315), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n511), .A2(new_n562), .A3(new_n603), .A4(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n460), .A2(new_n648), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n344), .A2(new_n331), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n452), .A2(new_n392), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n449), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n321), .A2(new_n323), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n409), .A2(new_n411), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n372), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n555), .A2(new_n642), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n646), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n505), .B2(new_n506), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n499), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n603), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT86), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n578), .A2(new_n599), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n511), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n578), .A2(new_n599), .A3(new_n661), .A4(new_n498), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n661), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n666), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n578), .A2(new_n599), .A3(new_n661), .A4(new_n498), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n662), .B1(new_n674), .B2(new_n667), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n485), .A2(G179), .A3(new_n494), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n508), .B(new_n676), .C1(new_n496), .C2(new_n444), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n510), .A3(new_n660), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n498), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT26), .B1(new_n679), .B2(new_n668), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(new_n680), .A3(KEYINPUT86), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n665), .B1(new_n673), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n657), .B1(new_n460), .B2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(new_n555), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n213), .A2(G20), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n250), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n524), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT87), .B1(new_n684), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n562), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n684), .A2(KEYINPUT87), .A3(new_n692), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT88), .B1(new_n695), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n691), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n647), .B1(new_n641), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n646), .A2(new_n701), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n659), .A2(new_n691), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT89), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(G399));
  NOR2_X1   g0510(.A1(new_n214), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G1), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n465), .A2(new_n384), .A3(new_n513), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n207), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n511), .A2(new_n667), .A3(new_n669), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n662), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n717), .B(new_n718), .C1(new_n659), .C2(new_n664), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .A3(new_n701), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n682), .A2(new_n691), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  AND4_X1   g0522(.A1(new_n614), .A2(new_n532), .A3(new_n540), .A4(new_n604), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n505), .A3(new_n576), .A4(new_n565), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n557), .A2(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n485), .A2(new_n494), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n573), .A3(new_n728), .A4(new_n615), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n691), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT31), .B(new_n691), .C1(new_n726), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT90), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n648), .B2(new_n691), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n532), .A2(new_n540), .A3(G179), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT84), .B1(new_n547), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n524), .A2(new_n551), .A3(new_n552), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(new_n560), .A3(new_n542), .A4(new_n550), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n642), .A2(new_n646), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n679), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(KEYINPUT90), .A3(new_n603), .A4(new_n701), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n735), .B1(new_n737), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n722), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n716), .B1(new_n751), .B2(G1), .ZN(G364));
  NAND2_X1  g0552(.A1(new_n685), .A2(G45), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT91), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n712), .A2(G1), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n697), .A2(new_n747), .A3(new_n698), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n700), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n214), .A2(new_n537), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n513), .B2(new_n214), .ZN(new_n759));
  AOI21_X1  g0559(.A(G45), .B1(new_n206), .B2(G50), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n239), .B2(G45), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n214), .A2(new_n291), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n759), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT92), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n246), .B1(G20), .B2(new_n444), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n755), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n275), .A2(new_n328), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n315), .A3(G200), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n270), .B1(new_n772), .B2(new_n476), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT93), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n275), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(G190), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n516), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G58), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n315), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n771), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n315), .A2(new_n497), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n775), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n786), .B1(new_n787), .B2(new_n789), .C1(new_n338), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n775), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n793), .A2(G179), .A3(new_n497), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n384), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n771), .A2(new_n790), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n775), .A2(new_n788), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n202), .B1(new_n798), .B2(new_n353), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n781), .A2(new_n792), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n802));
  INV_X1    g0602(.A(G326), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n797), .A2(new_n803), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G294), .B2(new_n783), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT95), .Z(new_n807));
  OR2_X1    g0607(.A1(new_n777), .A2(KEYINPUT96), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n777), .A2(KEYINPUT96), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G329), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT33), .B(G317), .Z(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n772), .B1(new_n814), .B2(new_n791), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n537), .B1(new_n795), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n789), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n815), .B(new_n817), .C1(G322), .C2(new_n818), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n807), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n801), .A2(new_n802), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n768), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n770), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n695), .A2(new_n696), .ZN(new_n825));
  INV_X1    g0625(.A(new_n767), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n757), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  OAI21_X1  g0629(.A(new_n396), .B1(new_n382), .B2(new_n701), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n393), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n392), .A2(new_n701), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n721), .B(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(new_n749), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n749), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n755), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n766), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n768), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT98), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n755), .B1(new_n842), .B2(new_n353), .ZN(new_n843));
  INV_X1    g0643(.A(new_n797), .ZN(new_n844));
  INV_X1    g0644(.A(new_n798), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n844), .A2(G137), .B1(new_n845), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  INV_X1    g0647(.A(G150), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n847), .B2(new_n789), .C1(new_n848), .C2(new_n791), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT34), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n784), .A2(new_n787), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n291), .B1(new_n202), .B2(new_n772), .C1(new_n795), .C2(new_n338), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(G132), .C2(new_n811), .ZN(new_n853));
  INV_X1    g0653(.A(new_n772), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n854), .A2(G107), .B1(new_n818), .B2(G294), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n794), .A2(G87), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n537), .A3(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n785), .B(new_n857), .C1(G311), .C2(new_n811), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n844), .A2(G303), .B1(new_n845), .B2(G116), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n816), .B2(new_n791), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n850), .A2(new_n853), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n843), .B1(new_n822), .B2(new_n862), .C1(new_n834), .C2(new_n766), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n838), .A2(new_n863), .ZN(G384));
  NAND2_X1  g0664(.A1(new_n279), .A2(G77), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n207), .A2(new_n865), .B1(G50), .B2(new_n338), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n213), .A3(new_n304), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT35), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n513), .B(new_n209), .C1(new_n593), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n868), .B2(new_n593), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT36), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  XOR2_X1   g0673(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n874));
  AND2_X1   g0674(.A1(new_n293), .A2(new_n249), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(new_n341), .B1(new_n261), .B2(new_n255), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT100), .B1(new_n876), .B2(new_n689), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT100), .ZN(new_n878));
  INV_X1    g0678(.A(new_n689), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n295), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n335), .A2(new_n342), .A3(new_n262), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT102), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n882), .A2(new_n883), .B1(new_n295), .B2(new_n319), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n876), .A2(KEYINPUT102), .A3(new_n335), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT37), .B1(new_n295), .B2(new_n319), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n332), .A2(new_n887), .A3(new_n343), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n886), .A2(KEYINPUT37), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n881), .B1(new_n650), .B2(new_n654), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n874), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT7), .B1(new_n291), .B2(G20), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n288), .A2(new_n269), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(G68), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT16), .B1(new_n894), .B2(new_n282), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n262), .B1(new_n294), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n319), .B2(new_n879), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n332), .A2(new_n343), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  AOI211_X1 g0699(.A(KEYINPUT100), .B(new_n689), .C1(new_n342), .C2(new_n262), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n878), .B1(new_n295), .B2(new_n879), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n332), .A2(new_n887), .A3(new_n343), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n898), .A2(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n896), .A2(new_n879), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n904), .B(KEYINPUT38), .C1(new_n345), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n891), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT104), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT104), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n891), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n423), .A2(new_n691), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n449), .A2(new_n452), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n449), .B2(new_n452), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n834), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n746), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n905), .B1(new_n650), .B2(new_n654), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n332), .A2(new_n897), .A3(new_n343), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n888), .A2(new_n881), .B1(KEYINPUT37), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n906), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n737), .A2(new_n745), .ZN(new_n925));
  INV_X1    g0725(.A(new_n735), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n915), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n918), .B1(new_n928), .B2(new_n911), .ZN(new_n929));
  AOI211_X1 g0729(.A(KEYINPUT103), .B(KEYINPUT40), .C1(new_n924), .C2(new_n927), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n917), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n746), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n459), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n747), .ZN(new_n935));
  INV_X1    g0735(.A(new_n665), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n675), .A2(new_n680), .A3(KEYINPUT86), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT86), .B1(new_n675), .B2(new_n680), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n701), .A3(new_n834), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n832), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n913), .A2(new_n914), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n924), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n654), .A2(new_n879), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n449), .A2(new_n691), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n923), .B2(new_n906), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n891), .A2(new_n949), .A3(new_n906), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n459), .B(new_n720), .C1(new_n721), .C2(KEYINPUT29), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n657), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n935), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT106), .Z(new_n959));
  INV_X1    g0759(.A(KEYINPUT105), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n250), .A2(new_n685), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n935), .B2(new_n957), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n962), .A2(new_n960), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n873), .B1(new_n963), .B2(new_n964), .ZN(G367));
  NAND2_X1  g0765(.A1(new_n754), .A2(G1), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n603), .B1(new_n600), .B2(new_n701), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n669), .A2(new_n691), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT44), .B1(new_n709), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n707), .B(KEYINPUT89), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n973), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT45), .B1(new_n709), .B2(new_n971), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n706), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n972), .A2(new_n976), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n705), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n700), .A2(new_n704), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n706), .A2(new_n555), .A3(new_n701), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n555), .A2(new_n701), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n700), .A2(new_n704), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n705), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n750), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n711), .B(KEYINPUT41), .Z(new_n993));
  OAI21_X1  g0793(.A(new_n967), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n706), .A2(new_n973), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT111), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n702), .A2(new_n988), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n971), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT42), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n701), .A2(new_n478), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT107), .ZN(new_n1003));
  MUX2_X1   g0803(.A(new_n663), .B(new_n662), .S(new_n1003), .Z(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n668), .B1(new_n969), .B2(new_n646), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT109), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g0808(.A(KEYINPUT109), .B(new_n668), .C1(new_n969), .C2(new_n646), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n701), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1001), .A2(new_n1005), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1004), .B(KEYINPUT43), .Z(new_n1013));
  AOI22_X1  g0813(.A1(new_n1011), .A2(KEYINPUT110), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT110), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1001), .A2(new_n1015), .A3(new_n1005), .A4(new_n1010), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n997), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1019));
  AND4_X1   g0819(.A1(new_n997), .A2(new_n1018), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n996), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1014), .A2(new_n997), .A3(new_n1016), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n995), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n994), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n755), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n769), .B1(new_n215), .B2(new_n375), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n763), .A2(new_n235), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n854), .A2(G116), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT46), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(KEYINPUT112), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(G317), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n795), .A2(new_n516), .B1(new_n777), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1031), .B2(KEYINPUT112), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n789), .A2(new_n813), .B1(new_n798), .B2(new_n816), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(G294), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n797), .A2(new_n804), .B1(new_n791), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n291), .B(new_n1041), .C1(G107), .C2(new_n783), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n848), .A2(new_n789), .B1(new_n791), .B2(new_n778), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n795), .A2(new_n353), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n777), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1044), .C1(G137), .C2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n270), .B1(new_n797), .B2(new_n847), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n772), .A2(new_n787), .B1(new_n798), .B2(new_n202), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G68), .C2(new_n783), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1039), .A2(new_n1042), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT47), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n822), .B1(new_n1050), .B2(KEYINPUT47), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1030), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1004), .B2(new_n826), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1026), .A2(new_n1054), .ZN(G387));
  NAND3_X1  g0855(.A1(new_n987), .A2(new_n751), .A3(new_n990), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n711), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n751), .B2(new_n991), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n763), .B1(new_n232), .B2(G45), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n714), .B2(new_n758), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n254), .A2(new_n202), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n338), .A2(new_n353), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1062), .A2(G45), .A3(new_n1063), .A4(new_n714), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1060), .A2(new_n1064), .B1(G107), .B2(new_n215), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n769), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n291), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n470), .B2(new_n783), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n789), .A2(new_n202), .B1(new_n777), .B2(new_n848), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G77), .B2(new_n854), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n794), .A2(G97), .B1(new_n844), .B2(G159), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n791), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1072), .A2(new_n254), .B1(new_n845), .B2(G68), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n798), .A2(new_n813), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n804), .A2(new_n791), .B1(new_n789), .B2(new_n1035), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G322), .C2(new_n844), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(KEYINPUT48), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n854), .A2(G294), .B1(G283), .B2(new_n783), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(KEYINPUT113), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1077), .A2(KEYINPUT48), .B1(new_n1082), .B2(new_n1079), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n794), .A2(G116), .B1(G326), .B2(new_n1045), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n1067), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT49), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1074), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n755), .B1(new_n1088), .B2(new_n768), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n704), .B2(new_n767), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n991), .B2(new_n966), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1058), .A2(new_n1092), .ZN(G393));
  NAND2_X1  g0893(.A1(new_n973), .A2(new_n767), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n769), .B1(new_n516), .B2(new_n215), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n763), .A2(new_n242), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1027), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n856), .B1(new_n202), .B2(new_n791), .C1(new_n253), .C2(new_n798), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1067), .B(new_n1098), .C1(G77), .C2(new_n783), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n797), .A2(new_n848), .B1(new_n789), .B2(new_n778), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n772), .A2(new_n338), .B1(new_n777), .B2(new_n847), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT114), .Z(new_n1103));
  NAND3_X1  g0903(.A1(new_n1099), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n797), .A2(new_n1035), .B1(new_n789), .B2(new_n804), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT52), .Z(new_n1106));
  AOI211_X1 g0906(.A(new_n270), .B(new_n796), .C1(G116), .C2(new_n783), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1072), .A2(G303), .B1(new_n1045), .B2(G322), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n854), .A2(G283), .B1(new_n845), .B2(G294), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1104), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1097), .B1(new_n1111), .B2(new_n768), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n985), .A2(new_n966), .B1(new_n1094), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n981), .A2(new_n984), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1056), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n711), .B1(new_n1056), .B2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT115), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1113), .B(KEYINPUT115), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(G390));
  NAND3_X1  g0921(.A1(new_n459), .A2(G330), .A3(new_n932), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n955), .A2(new_n657), .A3(new_n1122), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n746), .A2(new_n747), .A3(new_n833), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n943), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n746), .A2(new_n747), .A3(new_n915), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n941), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n719), .A2(new_n701), .A3(new_n831), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n832), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n914), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT116), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n449), .A2(new_n452), .A3(new_n912), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT116), .B1(new_n913), .B2(new_n914), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1130), .B1(new_n1136), .B2(new_n1124), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1123), .B1(new_n1127), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n942), .B1(new_n940), .B2(new_n832), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n948), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n951), .B(new_n952), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n908), .A2(new_n1143), .A3(new_n910), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1126), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1139), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1141), .B1(new_n941), .B2(new_n943), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n951), .A2(new_n952), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1126), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n1138), .A3(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n711), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n966), .A3(new_n1146), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n795), .A2(new_n338), .B1(new_n384), .B2(new_n791), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n270), .B(new_n1157), .C1(G87), .C2(new_n854), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n783), .A2(G77), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n811), .A2(G294), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n789), .A2(new_n513), .B1(new_n798), .B2(new_n516), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G283), .B2(new_n844), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n795), .A2(new_n202), .B1(new_n1164), .B2(new_n797), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n537), .B(new_n1165), .C1(G132), .C2(new_n818), .ZN(new_n1166));
  INV_X1    g0966(.A(G137), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n791), .A2(new_n1167), .B1(new_n798), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT117), .Z(new_n1170));
  INV_X1    g0970(.A(G125), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1166), .B(new_n1170), .C1(new_n1171), .C2(new_n810), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1173));
  OR3_X1    g0973(.A1(new_n772), .A2(new_n1173), .A3(new_n848), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n772), .B2(new_n848), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n778), .C2(new_n784), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1163), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n768), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n755), .B1(new_n842), .B2(new_n253), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(new_n1151), .C2(new_n766), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1155), .A2(new_n1156), .A3(new_n1180), .ZN(G378));
  OAI211_X1 g0981(.A(G330), .B(new_n917), .C1(new_n929), .C2(new_n930), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n372), .B1(new_n409), .B2(new_n411), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n371), .A2(new_n879), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1184), .B(new_n1185), .Z(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n945), .B1(new_n1140), .B2(new_n924), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n891), .A2(new_n949), .A3(new_n906), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1141), .B1(new_n1190), .B2(new_n950), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1188), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n1191), .A2(new_n944), .A3(new_n946), .A4(new_n1188), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1188), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n947), .B2(new_n953), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1189), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1182), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n967), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G41), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n772), .B2(new_n353), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G116), .A2(new_n844), .B1(new_n818), .B2(G107), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n516), .B2(new_n791), .C1(new_n810), .C2(new_n816), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n795), .A2(new_n787), .B1(new_n798), .B2(new_n375), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1067), .B1(new_n784), .B2(new_n338), .ZN(new_n1205));
  OR4_X1    g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1200), .B1(new_n1067), .B2(new_n244), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1206), .A2(new_n1207), .B1(new_n202), .B2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  INV_X1    g1010(.A(G132), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n797), .A2(new_n1171), .B1(new_n791), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1168), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n854), .A2(new_n1213), .B1(new_n818), .B2(G128), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1167), .B2(new_n798), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1212), .B(new_n1215), .C1(G150), .C2(new_n783), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n244), .B(new_n1200), .C1(new_n795), .C2(new_n778), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G124), .B2(new_n1045), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT59), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1218), .A2(new_n1222), .B1(new_n1207), .B2(new_n1206), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n768), .B1(new_n1210), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n755), .B1(new_n202), .B2(new_n840), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1195), .C2(new_n766), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT120), .Z(new_n1227));
  NOR2_X1   g1027(.A1(new_n1199), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1123), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1154), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT57), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1230), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1229), .B1(new_n1237), .B2(new_n711), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n1127), .A2(new_n1137), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n966), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1027), .B1(new_n841), .B2(G68), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT121), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n795), .A2(new_n787), .B1(new_n778), .B2(new_n772), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G150), .B2(new_n845), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1067), .B1(G50), .B2(new_n783), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n1164), .C2(new_n810), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT122), .Z(new_n1248));
  AOI22_X1  g1048(.A1(G132), .A2(new_n844), .B1(new_n1072), .B2(new_n1213), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1167), .B2(new_n789), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1044), .A2(new_n270), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G116), .A2(new_n1072), .B1(new_n818), .B2(G283), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n375), .C2(new_n784), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n854), .A2(G97), .B1(new_n845), .B2(G107), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n1040), .B2(new_n797), .C1(new_n810), .C2(new_n813), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1248), .A2(new_n1250), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1243), .B1(new_n1256), .B2(new_n768), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1136), .B2(new_n766), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1241), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n993), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1127), .A2(new_n1123), .A3(new_n1137), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1139), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT123), .Z(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(G381));
  NOR2_X1   g1066(.A1(G375), .A2(G378), .ZN(new_n1267));
  AND4_X1   g1067(.A1(new_n1026), .A2(new_n1119), .A3(new_n1054), .A4(new_n1120), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1058), .A2(new_n1092), .A3(new_n828), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(G381), .A2(G384), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1270), .ZN(G407));
  INV_X1    g1071(.A(G213), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(G343), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1267), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(G213), .A3(new_n1274), .ZN(G409));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1269), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1026), .A2(new_n1054), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1268), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(G390), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1026), .A2(new_n1119), .A3(new_n1054), .A4(new_n1120), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1277), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1230), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1235), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n711), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G378), .A3(new_n1228), .ZN(new_n1288));
  INV_X1    g1088(.A(G378), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1230), .A2(new_n1232), .A3(new_n1261), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1228), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1273), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT124), .B1(new_n1240), .B2(new_n1231), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1262), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(new_n1296), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1139), .A2(new_n1262), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n712), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1295), .B1(new_n1303), .B2(new_n1259), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1262), .B1(new_n1138), .B2(KEYINPUT124), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1301), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1138), .A2(new_n1306), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1305), .A2(new_n1296), .B1(new_n1307), .B2(new_n1262), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1260), .C1(new_n1308), .C2(new_n712), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1304), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1293), .A2(new_n1294), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT62), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1273), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1315));
  INV_X1    g1115(.A(G2897), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1294), .A2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1304), .A2(new_n1309), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1304), .B2(new_n1309), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(KEYINPUT127), .B(new_n1314), .C1(new_n1315), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1315), .A2(new_n1322), .A3(new_n1311), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1313), .A2(new_n1321), .A3(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1319), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1304), .A2(new_n1309), .A3(new_n1317), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(G378), .B1(new_n1290), .B2(new_n1228), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1238), .B2(G378), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1327), .B1(new_n1329), .B2(new_n1273), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT127), .B1(new_n1330), .B2(new_n1314), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1284), .B1(new_n1324), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1325), .A2(new_n1333), .A3(new_n1326), .ZN(new_n1334));
  OAI21_X1  g1134(.A(KEYINPUT126), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1315), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1280), .A2(new_n1314), .A3(new_n1283), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT125), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1312), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1312), .A2(new_n1339), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT63), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1338), .A2(new_n1341), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1332), .A2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(new_n1284), .A2(new_n1310), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1280), .A2(new_n1283), .A3(new_n1311), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(G375), .B(G378), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1348), .B(new_n1349), .ZN(G402));
endmodule


