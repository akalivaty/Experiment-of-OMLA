

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U554 ( .A(n700), .B(KEYINPUT95), .ZN(n702) );
  INV_X1 U555 ( .A(KEYINPUT83), .ZN(n547) );
  NAND2_X1 U556 ( .A1(n876), .A2(G137), .ZN(n524) );
  XOR2_X1 U557 ( .A(n722), .B(KEYINPUT29), .Z(n519) );
  NOR2_X1 U558 ( .A1(n814), .A2(n744), .ZN(n520) );
  NOR2_X1 U559 ( .A1(n754), .A2(n752), .ZN(n695) );
  INV_X1 U560 ( .A(n695), .ZN(n704) );
  INV_X1 U561 ( .A(n922), .ZN(n701) );
  AND2_X1 U562 ( .A1(n702), .A2(n701), .ZN(n709) );
  BUF_X1 U563 ( .A(n695), .Z(n713) );
  XNOR2_X1 U564 ( .A(KEYINPUT99), .B(KEYINPUT32), .ZN(n730) );
  INV_X1 U565 ( .A(KEYINPUT64), .ZN(n746) );
  INV_X1 U566 ( .A(KEYINPUT17), .ZN(n521) );
  INV_X1 U567 ( .A(KEYINPUT33), .ZN(n748) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n643) );
  NOR2_X1 U569 ( .A1(G651), .A2(n630), .ZN(n644) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n528), .ZN(n872) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n532), .Z(n642) );
  NOR2_X1 U572 ( .A1(n531), .A2(n530), .ZN(G160) );
  XNOR2_X2 U573 ( .A(n522), .B(n521), .ZN(n876) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n873) );
  NAND2_X1 U575 ( .A1(G113), .A2(n873), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n525), .B(KEYINPUT67), .ZN(n527) );
  INV_X1 U578 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G125), .A2(n872), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n531) );
  AND2_X1 U581 ( .A1(n528), .A2(G2104), .ZN(n877) );
  NAND2_X1 U582 ( .A1(G101), .A2(n877), .ZN(n529) );
  XNOR2_X1 U583 ( .A(KEYINPUT23), .B(n529), .ZN(n530) );
  INV_X1 U584 ( .A(G651), .ZN(n536) );
  NOR2_X1 U585 ( .A1(G543), .A2(n536), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G64), .A2(n642), .ZN(n535) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n533) );
  XNOR2_X1 U588 ( .A(KEYINPUT68), .B(n533), .ZN(n630) );
  NAND2_X1 U589 ( .A1(G52), .A2(n644), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G90), .A2(n643), .ZN(n539) );
  OR2_X1 U592 ( .A1(n536), .A2(n630), .ZN(n537) );
  XNOR2_X1 U593 ( .A(KEYINPUT69), .B(n537), .ZN(n649) );
  NAND2_X1 U594 ( .A1(G77), .A2(n649), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U597 ( .A1(n542), .A2(n541), .ZN(G171) );
  INV_X1 U598 ( .A(G171), .ZN(G301) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G132), .ZN(G219) );
  INV_X1 U601 ( .A(G82), .ZN(G220) );
  NAND2_X1 U602 ( .A1(G138), .A2(n876), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G102), .A2(n877), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G126), .A2(n872), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G114), .A2(n873), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U608 ( .A(n548), .B(n547), .ZN(n549) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n676) );
  BUF_X1 U610 ( .A(n676), .Z(G164) );
  NAND2_X1 U611 ( .A1(G62), .A2(n642), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G50), .A2(n644), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U614 ( .A(KEYINPUT81), .B(n553), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G88), .A2(n643), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G75), .A2(n649), .ZN(n554) );
  AND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(G303) );
  NAND2_X1 U619 ( .A1(n643), .A2(G89), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G76), .A2(n649), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G63), .A2(n642), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G51), .A2(n644), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G94), .A2(G452), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT70), .B(n568), .Z(G173) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U634 ( .A(n569), .B(KEYINPUT10), .Z(n828) );
  NAND2_X1 U635 ( .A1(n828), .A2(G567), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n642), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U639 ( .A1(n643), .A2(G81), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G68), .A2(n649), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n644), .A2(G43), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n922) );
  INV_X1 U647 ( .A(G860), .ZN(n600) );
  OR2_X1 U648 ( .A1(n922), .A2(n600), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT73), .B(n580), .Z(G153) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G66), .A2(n642), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G92), .A2(n643), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G79), .A2(n649), .ZN(n584) );
  NAND2_X1 U655 ( .A1(G54), .A2(n644), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n587), .Z(n921) );
  OR2_X1 U659 ( .A1(n921), .A2(G868), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G53), .A2(n644), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT72), .B(n590), .Z(n595) );
  NAND2_X1 U663 ( .A1(G91), .A2(n643), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G78), .A2(n649), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT71), .B(n593), .Z(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n642), .A2(G65), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(G299) );
  INV_X1 U670 ( .A(G868), .ZN(n659) );
  NOR2_X1 U671 ( .A1(G286), .A2(n659), .ZN(n599) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n601), .A2(n921), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT16), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n603), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n922), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G868), .A2(n921), .ZN(n604) );
  NOR2_X1 U680 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n872), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT18), .B(n607), .Z(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT75), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G111), .A2(n873), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G135), .A2(n876), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G99), .A2(n877), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n977) );
  XNOR2_X1 U691 ( .A(n977), .B(G2096), .ZN(n615) );
  INV_X1 U692 ( .A(G2100), .ZN(n847) );
  NAND2_X1 U693 ( .A1(n615), .A2(n847), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G67), .A2(n642), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G93), .A2(n643), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G80), .A2(n649), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G55), .A2(n644), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n660) );
  XNOR2_X1 U701 ( .A(n922), .B(KEYINPUT76), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n921), .A2(G559), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n623), .B(n622), .ZN(n657) );
  NOR2_X1 U704 ( .A1(n657), .A2(G860), .ZN(n624) );
  XOR2_X1 U705 ( .A(KEYINPUT77), .B(n624), .Z(n625) );
  XOR2_X1 U706 ( .A(n660), .B(n625), .Z(G145) );
  NAND2_X1 U707 ( .A1(n644), .A2(G49), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT78), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n642), .A2(n629), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n630), .A2(G87), .ZN(n631) );
  XOR2_X1 U713 ( .A(KEYINPUT79), .B(n631), .Z(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G73), .A2(n649), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G86), .A2(n643), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G48), .A2(n644), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n642), .A2(G61), .ZN(n637) );
  XOR2_X1 U721 ( .A(KEYINPUT80), .B(n637), .Z(n638) );
  NOR2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(G305) );
  AND2_X1 U724 ( .A1(n642), .A2(G60), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G85), .A2(n643), .ZN(n646) );
  NAND2_X1 U726 ( .A1(G47), .A2(n644), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n649), .A2(G72), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G290) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(G288), .ZN(n656) );
  XOR2_X1 U732 ( .A(G299), .B(G303), .Z(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(G305), .ZN(n653) );
  XOR2_X1 U734 ( .A(n660), .B(n653), .Z(n654) );
  XNOR2_X1 U735 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n656), .B(n655), .ZN(n900) );
  XOR2_X1 U737 ( .A(n900), .B(n657), .Z(n658) );
  NOR2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U739 ( .A1(G868), .A2(n660), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U743 ( .A1(n664), .A2(G2090), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n665), .B(KEYINPUT21), .ZN(n666) );
  XNOR2_X1 U745 ( .A(KEYINPUT82), .B(n666), .ZN(n667) );
  NAND2_X1 U746 ( .A1(G2072), .A2(n667), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U750 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G96), .A2(n670), .ZN(n832) );
  NAND2_X1 U752 ( .A1(n832), .A2(G2106), .ZN(n674) );
  NAND2_X1 U753 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U754 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U755 ( .A1(G108), .A2(n672), .ZN(n833) );
  NAND2_X1 U756 ( .A1(n833), .A2(G567), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n674), .A2(n673), .ZN(n855) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U759 ( .A1(n855), .A2(n675), .ZN(n831) );
  NAND2_X1 U760 ( .A1(n831), .A2(G36), .ZN(G176) );
  NOR2_X1 U761 ( .A1(n676), .A2(G1384), .ZN(n677) );
  XNOR2_X1 U762 ( .A(KEYINPUT65), .B(n677), .ZN(n754) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n752) );
  NAND2_X1 U764 ( .A1(G8), .A2(n704), .ZN(n814) );
  NOR2_X1 U765 ( .A1(G1966), .A2(n814), .ZN(n737) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n704), .ZN(n734) );
  NOR2_X1 U767 ( .A1(n737), .A2(n734), .ZN(n678) );
  NAND2_X1 U768 ( .A1(G8), .A2(n678), .ZN(n679) );
  XNOR2_X1 U769 ( .A(KEYINPUT30), .B(n679), .ZN(n680) );
  NOR2_X1 U770 ( .A1(G168), .A2(n680), .ZN(n681) );
  XNOR2_X1 U771 ( .A(n681), .B(KEYINPUT97), .ZN(n687) );
  XOR2_X1 U772 ( .A(G2078), .B(KEYINPUT25), .Z(n682) );
  XNOR2_X1 U773 ( .A(KEYINPUT92), .B(n682), .ZN(n1010) );
  NAND2_X1 U774 ( .A1(n713), .A2(n1010), .ZN(n684) );
  NAND2_X1 U775 ( .A1(G1961), .A2(n704), .ZN(n683) );
  NAND2_X1 U776 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U777 ( .A(KEYINPUT93), .B(n685), .ZN(n723) );
  OR2_X1 U778 ( .A1(n723), .A2(G171), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U780 ( .A(KEYINPUT31), .B(n688), .ZN(n732) );
  INV_X1 U781 ( .A(G8), .ZN(n694) );
  NOR2_X1 U782 ( .A1(G2090), .A2(n704), .ZN(n689) );
  XNOR2_X1 U783 ( .A(n689), .B(KEYINPUT98), .ZN(n691) );
  NOR2_X1 U784 ( .A1(n814), .A2(G1971), .ZN(n690) );
  NOR2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n692), .A2(G303), .ZN(n693) );
  OR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n726) );
  AND2_X1 U788 ( .A1(n732), .A2(n726), .ZN(n725) );
  XOR2_X1 U789 ( .A(G1996), .B(KEYINPUT94), .Z(n1011) );
  NOR2_X1 U790 ( .A1(n704), .A2(n1011), .ZN(n697) );
  XOR2_X1 U791 ( .A(KEYINPUT66), .B(KEYINPUT26), .Z(n696) );
  XNOR2_X1 U792 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n704), .A2(G1341), .ZN(n698) );
  NAND2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n921), .A2(n709), .ZN(n708) );
  AND2_X1 U796 ( .A1(n713), .A2(G2067), .ZN(n703) );
  XOR2_X1 U797 ( .A(n703), .B(KEYINPUT96), .Z(n706) );
  NAND2_X1 U798 ( .A1(n704), .A2(G1348), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n711) );
  OR2_X1 U801 ( .A1(n921), .A2(n709), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n717) );
  INV_X1 U803 ( .A(G299), .ZN(n927) );
  NAND2_X1 U804 ( .A1(n713), .A2(G2072), .ZN(n712) );
  XNOR2_X1 U805 ( .A(n712), .B(KEYINPUT27), .ZN(n715) );
  INV_X1 U806 ( .A(G1956), .ZN(n836) );
  NOR2_X1 U807 ( .A1(n836), .A2(n713), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n927), .A2(n718), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n927), .A2(n718), .ZN(n719) );
  XOR2_X1 U812 ( .A(n719), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U814 ( .A1(G171), .A2(n723), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n519), .A2(n724), .ZN(n733) );
  NAND2_X1 U816 ( .A1(n725), .A2(n733), .ZN(n729) );
  INV_X1 U817 ( .A(n726), .ZN(n727) );
  OR2_X1 U818 ( .A1(n727), .A2(G286), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U820 ( .A(n731), .B(n730), .ZN(n740) );
  NAND2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U822 ( .A1(G8), .A2(n734), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n738) );
  NOR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n806) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U828 ( .A1(n750), .A2(n741), .ZN(n930) );
  XOR2_X1 U829 ( .A(n930), .B(KEYINPUT100), .Z(n742) );
  NOR2_X1 U830 ( .A1(n806), .A2(n742), .ZN(n743) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT101), .ZN(n745) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n929) );
  INV_X1 U833 ( .A(n929), .ZN(n744) );
  AND2_X1 U834 ( .A1(n745), .A2(n520), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n805) );
  NAND2_X1 U837 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n751), .A2(n814), .ZN(n803) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n942) );
  INV_X1 U840 ( .A(n752), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n785) );
  INV_X1 U842 ( .A(n785), .ZN(n799) );
  XNOR2_X1 U843 ( .A(G2067), .B(KEYINPUT37), .ZN(n795) );
  NAND2_X1 U844 ( .A1(G140), .A2(n876), .ZN(n756) );
  NAND2_X1 U845 ( .A1(G104), .A2(n877), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U847 ( .A(KEYINPUT34), .B(n757), .ZN(n763) );
  NAND2_X1 U848 ( .A1(G128), .A2(n872), .ZN(n759) );
  NAND2_X1 U849 ( .A1(G116), .A2(n873), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U851 ( .A(KEYINPUT85), .B(n760), .ZN(n761) );
  XNOR2_X1 U852 ( .A(KEYINPUT35), .B(n761), .ZN(n762) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U854 ( .A(KEYINPUT36), .B(n764), .ZN(n895) );
  NOR2_X1 U855 ( .A1(n795), .A2(n895), .ZN(n765) );
  XNOR2_X1 U856 ( .A(n765), .B(KEYINPUT86), .ZN(n986) );
  NAND2_X1 U857 ( .A1(n799), .A2(n986), .ZN(n793) );
  XOR2_X1 U858 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n767) );
  NAND2_X1 U859 ( .A1(G105), .A2(n877), .ZN(n766) );
  XNOR2_X1 U860 ( .A(n767), .B(n766), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G129), .A2(n872), .ZN(n769) );
  NAND2_X1 U862 ( .A1(G117), .A2(n873), .ZN(n768) );
  NAND2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U864 ( .A(KEYINPUT89), .B(n770), .Z(n771) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n876), .A2(G141), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n888) );
  AND2_X1 U868 ( .A1(n888), .A2(G1996), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G95), .A2(n877), .ZN(n775) );
  XNOR2_X1 U870 ( .A(n775), .B(KEYINPUT88), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G119), .A2(n872), .ZN(n777) );
  NAND2_X1 U872 ( .A1(G131), .A2(n876), .ZN(n776) );
  NAND2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U874 ( .A1(G107), .A2(n873), .ZN(n778) );
  XNOR2_X1 U875 ( .A(KEYINPUT87), .B(n778), .ZN(n779) );
  NOR2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n884) );
  AND2_X1 U878 ( .A1(n884), .A2(G1991), .ZN(n783) );
  NOR2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n979) );
  NOR2_X1 U880 ( .A1(n979), .A2(n785), .ZN(n790) );
  INV_X1 U881 ( .A(n790), .ZN(n786) );
  AND2_X1 U882 ( .A1(n793), .A2(n786), .ZN(n818) );
  AND2_X1 U883 ( .A1(n942), .A2(n818), .ZN(n801) );
  NOR2_X1 U884 ( .A1(G1996), .A2(n888), .ZN(n983) );
  NOR2_X1 U885 ( .A1(n884), .A2(G1991), .ZN(n787) );
  XNOR2_X1 U886 ( .A(n787), .B(KEYINPUT102), .ZN(n976) );
  NOR2_X1 U887 ( .A1(G1986), .A2(G290), .ZN(n788) );
  NOR2_X1 U888 ( .A1(n976), .A2(n788), .ZN(n789) );
  NOR2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n983), .A2(n791), .ZN(n792) );
  XNOR2_X1 U891 ( .A(KEYINPUT39), .B(n792), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n895), .A2(n795), .ZN(n990) );
  NAND2_X1 U894 ( .A1(n796), .A2(n990), .ZN(n797) );
  AND2_X1 U895 ( .A1(n797), .A2(n799), .ZN(n819) );
  XNOR2_X1 U896 ( .A(G1986), .B(KEYINPUT84), .ZN(n798) );
  XNOR2_X1 U897 ( .A(n798), .B(G290), .ZN(n935) );
  NAND2_X1 U898 ( .A1(n935), .A2(n799), .ZN(n800) );
  OR2_X1 U899 ( .A1(n819), .A2(n800), .ZN(n822) );
  NAND2_X1 U900 ( .A1(n801), .A2(n822), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n824) );
  INV_X1 U903 ( .A(n806), .ZN(n809) );
  NOR2_X1 U904 ( .A1(G2090), .A2(G303), .ZN(n807) );
  NAND2_X1 U905 ( .A1(G8), .A2(n807), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n810), .A2(n814), .ZN(n816) );
  NOR2_X1 U908 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n811), .B(KEYINPUT24), .ZN(n812) );
  XNOR2_X1 U910 ( .A(KEYINPUT91), .B(n812), .ZN(n813) );
  OR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  AND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n820) );
  OR2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n825) );
  XNOR2_X1 U918 ( .A(n826), .B(n825), .ZN(G329) );
  NAND2_X1 U919 ( .A1(n828), .A2(G2106), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n827), .B(KEYINPUT106), .ZN(G217) );
  INV_X1 U921 ( .A(n828), .ZN(G223) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U932 ( .A(G1996), .B(KEYINPUT41), .ZN(n844) );
  XOR2_X1 U933 ( .A(G1981), .B(G1961), .Z(n835) );
  XNOR2_X1 U934 ( .A(G1991), .B(G1966), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n840) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n838) );
  XOR2_X1 U937 ( .A(G1986), .B(n836), .Z(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U940 ( .A(KEYINPUT108), .B(G2474), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2084), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2078), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n850) );
  XNOR2_X1 U947 ( .A(G2072), .B(G2090), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT43), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2678), .B(KEYINPUT107), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n854), .B(n853), .Z(G227) );
  INV_X1 U953 ( .A(n855), .ZN(G319) );
  NAND2_X1 U954 ( .A1(G124), .A2(n872), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n856), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G136), .A2(n876), .ZN(n857) );
  XOR2_X1 U957 ( .A(KEYINPUT109), .B(n857), .Z(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G112), .A2(n873), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G100), .A2(n877), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U963 ( .A1(G139), .A2(n876), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G103), .A2(n877), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(n866), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G127), .A2(n872), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G115), .A2(n873), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n993) );
  NAND2_X1 U972 ( .A1(G130), .A2(n872), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G118), .A2(n873), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U975 ( .A1(G142), .A2(n876), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n880), .Z(n881) );
  NOR2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n993), .B(n883), .ZN(n894) );
  XOR2_X1 U981 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n886) );
  XOR2_X1 U982 ( .A(n884), .B(KEYINPUT48), .Z(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U984 ( .A(G160), .B(n887), .ZN(n892) );
  XOR2_X1 U985 ( .A(n977), .B(G162), .Z(n890) );
  XOR2_X1 U986 ( .A(G164), .B(n888), .Z(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U990 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n922), .B(G286), .ZN(n899) );
  XOR2_X1 U993 ( .A(G301), .B(n921), .Z(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n917) );
  XNOR2_X1 U1000 ( .A(G2427), .B(KEYINPUT105), .ZN(n914) );
  XOR2_X1 U1001 ( .A(G2443), .B(G2438), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2430), .B(G2454), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1004 ( .A(KEYINPUT104), .B(G2435), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2446), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n915), .A2(G14), .ZN(n920) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n920), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(KEYINPUT56), .B(G16), .ZN(n948) );
  XOR2_X1 U1020 ( .A(G301), .B(G1961), .Z(n926) );
  XOR2_X1 U1021 ( .A(G1348), .B(n921), .Z(n924) );
  XNOR2_X1 U1022 ( .A(n922), .B(G1341), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n940) );
  XOR2_X1 U1025 ( .A(G1956), .B(n927), .Z(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT119), .ZN(n937) );
  AND2_X1 U1027 ( .A1(G303), .A2(G1971), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT120), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT121), .B(n938), .Z(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(KEYINPUT122), .B(n941), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(KEYINPUT57), .B(n944), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n1006) );
  XOR2_X1 U1041 ( .A(KEYINPUT124), .B(G4), .Z(n950) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n950), .B(n949), .ZN(n957) );
  XOR2_X1 U1044 ( .A(G1341), .B(G19), .Z(n952) );
  XOR2_X1 U1045 ( .A(G1956), .B(G20), .Z(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G6), .B(G1981), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(n955), .B(KEYINPUT123), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n958), .B(KEYINPUT125), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n959), .B(KEYINPUT60), .ZN(n966) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n963) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1060 ( .A(G1966), .B(KEYINPUT126), .Z(n967) );
  XNOR2_X1 U1061 ( .A(G21), .B(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G5), .B(G1961), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1065 ( .A(KEYINPUT61), .B(n972), .Z(n973) );
  NOR2_X1 U1066 ( .A1(G16), .A2(n973), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(KEYINPUT127), .B(n974), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n975), .A2(G11), .ZN(n1004) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n981) );
  XOR2_X1 U1071 ( .A(G160), .B(G2084), .Z(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n988) );
  XOR2_X1 U1073 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT51), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n989), .B(KEYINPUT113), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(KEYINPUT114), .B(n992), .ZN(n998) );
  XOR2_X1 U1081 ( .A(G2072), .B(n993), .Z(n995) );
  XOR2_X1 U1082 ( .A(G164), .B(G2078), .Z(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1084 ( .A(KEYINPUT50), .B(n996), .Z(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(n999), .B(KEYINPUT52), .ZN(n1000) );
  INV_X1 U1087 ( .A(KEYINPUT55), .ZN(n1028) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n1028), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(G29), .A2(n1001), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT115), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1031) );
  XNOR2_X1 U1093 ( .A(G2084), .B(G34), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(KEYINPUT54), .ZN(n1026) );
  XNOR2_X1 U1095 ( .A(G2090), .B(G35), .ZN(n1023) );
  XOR2_X1 U1096 ( .A(G1991), .B(G25), .Z(n1008) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(G28), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT116), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(n1010), .B(G27), .Z(n1013) );
  XNOR2_X1 U1100 ( .A(G32), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(G2067), .B(G26), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G33), .B(G2072), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(n1020), .B(KEYINPUT117), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT53), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT118), .B(n1024), .Z(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1028), .B(n1027), .ZN(n1029) );
  NOR2_X1 U1113 ( .A1(G29), .A2(n1029), .ZN(n1030) );
  NOR2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(n1032), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
  INV_X1 U1117 ( .A(G303), .ZN(G166) );
endmodule

