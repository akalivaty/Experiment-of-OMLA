

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U558 ( .A1(n779), .A2(n615), .ZN(n616) );
  NAND2_X1 U559 ( .A1(n891), .A2(G101), .ZN(n561) );
  XNOR2_X2 U560 ( .A(n556), .B(KEYINPUT67), .ZN(n690) );
  NAND2_X1 U561 ( .A1(n735), .A2(n753), .ZN(n526) );
  XOR2_X1 U562 ( .A(KEYINPUT26), .B(n613), .Z(n527) );
  OR2_X1 U563 ( .A1(KEYINPUT33), .A2(n686), .ZN(n528) );
  AND2_X1 U564 ( .A1(n632), .A2(G1996), .ZN(n613) );
  XNOR2_X1 U565 ( .A(n654), .B(KEYINPUT30), .ZN(n655) );
  INV_X1 U566 ( .A(KEYINPUT99), .ZN(n662) );
  INV_X1 U567 ( .A(G2104), .ZN(n555) );
  NOR2_X1 U568 ( .A1(n526), .A2(n737), .ZN(n738) );
  NOR2_X1 U569 ( .A1(G651), .A2(n544), .ZN(n792) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n552), .Z(n888) );
  XNOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .ZN(n529) );
  XNOR2_X1 U572 ( .A(n529), .B(KEYINPUT69), .ZN(n544) );
  NAND2_X1 U573 ( .A1(G87), .A2(n544), .ZN(n530) );
  XNOR2_X1 U574 ( .A(n530), .B(KEYINPUT82), .ZN(n537) );
  INV_X1 U575 ( .A(G651), .ZN(n543) );
  NOR2_X1 U576 ( .A1(G543), .A2(n543), .ZN(n531) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n531), .Z(n532) );
  XNOR2_X1 U578 ( .A(KEYINPUT70), .B(n532), .ZN(n785) );
  NAND2_X1 U579 ( .A1(G49), .A2(n792), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G74), .A2(G651), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U582 ( .A1(n785), .A2(n535), .ZN(n536) );
  NAND2_X1 U583 ( .A1(n537), .A2(n536), .ZN(G288) );
  NAND2_X1 U584 ( .A1(n792), .A2(G51), .ZN(n539) );
  NAND2_X1 U585 ( .A1(G63), .A2(n785), .ZN(n538) );
  NAND2_X1 U586 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n540), .B(KEYINPUT75), .ZN(n541) );
  XNOR2_X1 U588 ( .A(n541), .B(KEYINPUT6), .ZN(n550) );
  XNOR2_X1 U589 ( .A(KEYINPUT5), .B(KEYINPUT74), .ZN(n548) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n788) );
  NAND2_X1 U591 ( .A1(n788), .A2(G89), .ZN(n542) );
  XNOR2_X1 U592 ( .A(n542), .B(KEYINPUT4), .ZN(n546) );
  NOR2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n784) );
  NAND2_X1 U594 ( .A1(G76), .A2(n784), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U596 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U597 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U598 ( .A(KEYINPUT7), .B(n551), .ZN(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U600 ( .A1(G2105), .A2(G2104), .ZN(n552) );
  NAND2_X1 U601 ( .A1(G138), .A2(n888), .ZN(n554) );
  NOR2_X4 U602 ( .A1(G2105), .A2(n555), .ZN(n891) );
  NAND2_X1 U603 ( .A1(G102), .A2(n891), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n554), .A2(n553), .ZN(n560) );
  AND2_X1 U605 ( .A1(n555), .A2(G2105), .ZN(n884) );
  NAND2_X1 U606 ( .A1(G126), .A2(n884), .ZN(n558) );
  NAND2_X1 U607 ( .A1(G2104), .A2(G2105), .ZN(n556) );
  NAND2_X1 U608 ( .A1(G114), .A2(n690), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U610 ( .A1(n560), .A2(n559), .ZN(G164) );
  XOR2_X1 U611 ( .A(n561), .B(KEYINPUT23), .Z(n563) );
  NAND2_X1 U612 ( .A1(n884), .A2(G125), .ZN(n562) );
  NAND2_X1 U613 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U614 ( .A(n564), .B(KEYINPUT66), .ZN(n569) );
  NAND2_X1 U615 ( .A1(G113), .A2(n690), .ZN(n565) );
  XNOR2_X1 U616 ( .A(n565), .B(KEYINPUT68), .ZN(n567) );
  NAND2_X1 U617 ( .A1(n888), .A2(G137), .ZN(n566) );
  NAND2_X1 U618 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U619 ( .A1(n569), .A2(n568), .ZN(G160) );
  NAND2_X1 U620 ( .A1(n792), .A2(G52), .ZN(n571) );
  NAND2_X1 U621 ( .A1(G64), .A2(n785), .ZN(n570) );
  NAND2_X1 U622 ( .A1(n571), .A2(n570), .ZN(n577) );
  NAND2_X1 U623 ( .A1(G90), .A2(n788), .ZN(n573) );
  NAND2_X1 U624 ( .A1(G77), .A2(n784), .ZN(n572) );
  NAND2_X1 U625 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  XNOR2_X1 U627 ( .A(KEYINPUT72), .B(n575), .ZN(n576) );
  NOR2_X1 U628 ( .A1(n577), .A2(n576), .ZN(G171) );
  NAND2_X1 U629 ( .A1(G75), .A2(n784), .ZN(n579) );
  NAND2_X1 U630 ( .A1(G50), .A2(n792), .ZN(n578) );
  NAND2_X1 U631 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U632 ( .A1(n788), .A2(G88), .ZN(n581) );
  NAND2_X1 U633 ( .A1(G62), .A2(n785), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U635 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U636 ( .A(n584), .B(KEYINPUT85), .Z(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(n784), .A2(G73), .ZN(n586) );
  XNOR2_X1 U639 ( .A(KEYINPUT84), .B(KEYINPUT2), .ZN(n585) );
  XNOR2_X1 U640 ( .A(n586), .B(n585), .ZN(n593) );
  NAND2_X1 U641 ( .A1(G86), .A2(n788), .ZN(n588) );
  NAND2_X1 U642 ( .A1(G48), .A2(n792), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U644 ( .A1(G61), .A2(n785), .ZN(n589) );
  XNOR2_X1 U645 ( .A(KEYINPUT83), .B(n589), .ZN(n590) );
  NOR2_X1 U646 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U647 ( .A1(n593), .A2(n592), .ZN(G305) );
  NAND2_X1 U648 ( .A1(G85), .A2(n788), .ZN(n595) );
  NAND2_X1 U649 ( .A1(G72), .A2(n784), .ZN(n594) );
  NAND2_X1 U650 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U651 ( .A1(n792), .A2(G47), .ZN(n597) );
  NAND2_X1 U652 ( .A1(G60), .A2(n785), .ZN(n596) );
  NAND2_X1 U653 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U654 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U655 ( .A(KEYINPUT71), .B(n600), .ZN(G290) );
  NAND2_X1 U656 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  NOR2_X2 U657 ( .A1(G164), .A2(G1384), .ZN(n687) );
  INV_X1 U658 ( .A(n687), .ZN(n601) );
  NAND2_X1 U659 ( .A1(G160), .A2(G40), .ZN(n688) );
  NOR2_X4 U660 ( .A1(n601), .A2(n688), .ZN(n632) );
  INV_X1 U661 ( .A(n632), .ZN(n664) );
  INV_X1 U662 ( .A(G1961), .ZN(n997) );
  NAND2_X1 U663 ( .A1(n664), .A2(n997), .ZN(n603) );
  XNOR2_X1 U664 ( .A(G2078), .B(KEYINPUT25), .ZN(n951) );
  NAND2_X1 U665 ( .A1(n632), .A2(n951), .ZN(n602) );
  NAND2_X1 U666 ( .A1(n603), .A2(n602), .ZN(n656) );
  NAND2_X1 U667 ( .A1(n656), .A2(G171), .ZN(n652) );
  NAND2_X1 U668 ( .A1(n785), .A2(G56), .ZN(n604) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n604), .Z(n610) );
  NAND2_X1 U670 ( .A1(n788), .A2(G81), .ZN(n605) );
  XNOR2_X1 U671 ( .A(n605), .B(KEYINPUT12), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G68), .A2(n784), .ZN(n606) );
  NAND2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U674 ( .A(KEYINPUT13), .B(n608), .Z(n609) );
  NOR2_X1 U675 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U676 ( .A1(n792), .A2(G43), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n612), .A2(n611), .ZN(n779) );
  NAND2_X1 U678 ( .A1(n664), .A2(G1341), .ZN(n614) );
  NAND2_X1 U679 ( .A1(n527), .A2(n614), .ZN(n615) );
  XNOR2_X1 U680 ( .A(n616), .B(KEYINPUT65), .ZN(n627) );
  NAND2_X1 U681 ( .A1(n788), .A2(G92), .ZN(n618) );
  NAND2_X1 U682 ( .A1(G66), .A2(n785), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U684 ( .A1(G79), .A2(n784), .ZN(n620) );
  NAND2_X1 U685 ( .A1(G54), .A2(n792), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U687 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U688 ( .A(KEYINPUT15), .B(n623), .ZN(n769) );
  INV_X1 U689 ( .A(n769), .ZN(n1006) );
  AND2_X1 U690 ( .A1(n664), .A2(G1348), .ZN(n625) );
  AND2_X1 U691 ( .A1(n632), .A2(G2067), .ZN(n624) );
  NOR2_X1 U692 ( .A1(n625), .A2(n624), .ZN(n628) );
  NOR2_X1 U693 ( .A1(n1006), .A2(n628), .ZN(n626) );
  OR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n644) );
  AND2_X1 U695 ( .A1(n628), .A2(n1006), .ZN(n642) );
  NAND2_X1 U696 ( .A1(G2072), .A2(n632), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT97), .B(n629), .ZN(n631) );
  INV_X1 U698 ( .A(KEYINPUT27), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(n634) );
  INV_X1 U700 ( .A(G1956), .ZN(n842) );
  NOR2_X1 U701 ( .A1(n632), .A2(n842), .ZN(n633) );
  NOR2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n645) );
  NAND2_X1 U703 ( .A1(n792), .A2(G53), .ZN(n636) );
  NAND2_X1 U704 ( .A1(G65), .A2(n785), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U706 ( .A1(G91), .A2(n788), .ZN(n638) );
  NAND2_X1 U707 ( .A1(G78), .A2(n784), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n1007) );
  AND2_X1 U710 ( .A1(n645), .A2(n1007), .ZN(n641) );
  NOR2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U713 ( .A1(n645), .A2(n1007), .ZN(n646) );
  XOR2_X1 U714 ( .A(n646), .B(KEYINPUT28), .Z(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n650) );
  XOR2_X1 U716 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n649) );
  XNOR2_X1 U717 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n661) );
  NAND2_X1 U719 ( .A1(G8), .A2(n664), .ZN(n745) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n745), .ZN(n675) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n664), .ZN(n672) );
  NOR2_X1 U722 ( .A1(n675), .A2(n672), .ZN(n653) );
  NAND2_X1 U723 ( .A1(G8), .A2(n653), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n655), .A2(G168), .ZN(n658) );
  NOR2_X1 U725 ( .A1(G171), .A2(n656), .ZN(n657) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT31), .B(n659), .Z(n660) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n673) );
  NAND2_X1 U729 ( .A1(G286), .A2(n673), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n669) );
  NOR2_X1 U731 ( .A1(G1971), .A2(n745), .ZN(n666) );
  NOR2_X1 U732 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U734 ( .A1(G303), .A2(n667), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n670), .A2(G8), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U738 ( .A1(G8), .A2(n672), .ZN(n677) );
  INV_X1 U739 ( .A(n673), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n739) );
  NOR2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NOR2_X1 U744 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n1000), .A2(n680), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n739), .A2(n681), .ZN(n682) );
  NAND2_X1 U747 ( .A1(n1001), .A2(n682), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT100), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n684), .A2(n745), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(KEYINPUT64), .ZN(n686) );
  XOR2_X1 U751 ( .A(G1981), .B(G305), .Z(n1017) );
  XNOR2_X1 U752 ( .A(G1986), .B(G290), .ZN(n999) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U754 ( .A(n689), .B(KEYINPUT92), .Z(n701) );
  INV_X1 U755 ( .A(n701), .ZN(n730) );
  NAND2_X1 U756 ( .A1(n999), .A2(n730), .ZN(n749) );
  AND2_X1 U757 ( .A1(n1017), .A2(n749), .ZN(n735) );
  NAND2_X1 U758 ( .A1(n690), .A2(G116), .ZN(n691) );
  XOR2_X1 U759 ( .A(KEYINPUT93), .B(n691), .Z(n693) );
  NAND2_X1 U760 ( .A1(n884), .A2(G128), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(KEYINPUT35), .ZN(n699) );
  NAND2_X1 U763 ( .A1(G140), .A2(n888), .ZN(n696) );
  NAND2_X1 U764 ( .A1(G104), .A2(n891), .ZN(n695) );
  NAND2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U766 ( .A(KEYINPUT34), .B(n697), .Z(n698) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U768 ( .A(n700), .B(KEYINPUT36), .Z(n876) );
  XNOR2_X1 U769 ( .A(KEYINPUT37), .B(G2067), .ZN(n728) );
  OR2_X1 U770 ( .A1(n876), .A2(n728), .ZN(n973) );
  NOR2_X1 U771 ( .A1(n701), .A2(n973), .ZN(n733) );
  NAND2_X1 U772 ( .A1(G129), .A2(n884), .ZN(n703) );
  NAND2_X1 U773 ( .A1(G117), .A2(n690), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U775 ( .A(KEYINPUT94), .B(n704), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n891), .A2(G105), .ZN(n705) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n705), .Z(n706) );
  NOR2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n888), .A2(G141), .ZN(n708) );
  NAND2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n881) );
  NOR2_X1 U781 ( .A1(G1996), .A2(n881), .ZN(n985) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n881), .ZN(n710) );
  XNOR2_X1 U783 ( .A(n710), .B(KEYINPUT95), .ZN(n718) );
  NAND2_X1 U784 ( .A1(G131), .A2(n888), .ZN(n712) );
  NAND2_X1 U785 ( .A1(G95), .A2(n891), .ZN(n711) );
  NAND2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U787 ( .A1(G119), .A2(n884), .ZN(n714) );
  NAND2_X1 U788 ( .A1(G107), .A2(n690), .ZN(n713) );
  NAND2_X1 U789 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U790 ( .A1(n716), .A2(n715), .ZN(n880) );
  AND2_X1 U791 ( .A1(G1991), .A2(n880), .ZN(n717) );
  NOR2_X1 U792 ( .A1(n718), .A2(n717), .ZN(n974) );
  XOR2_X1 U793 ( .A(KEYINPUT96), .B(n730), .Z(n719) );
  NOR2_X1 U794 ( .A1(n974), .A2(n719), .ZN(n732) );
  NOR2_X1 U795 ( .A1(G1991), .A2(n880), .ZN(n720) );
  XOR2_X1 U796 ( .A(KEYINPUT101), .B(n720), .Z(n978) );
  NOR2_X1 U797 ( .A1(G1986), .A2(G290), .ZN(n721) );
  NOR2_X1 U798 ( .A1(n978), .A2(n721), .ZN(n722) );
  NOR2_X1 U799 ( .A1(n732), .A2(n722), .ZN(n723) );
  XNOR2_X1 U800 ( .A(n723), .B(KEYINPUT102), .ZN(n724) );
  NOR2_X1 U801 ( .A1(n985), .A2(n724), .ZN(n725) );
  XOR2_X1 U802 ( .A(KEYINPUT39), .B(n725), .Z(n726) );
  NOR2_X1 U803 ( .A1(n733), .A2(n726), .ZN(n727) );
  XNOR2_X1 U804 ( .A(n727), .B(KEYINPUT103), .ZN(n729) );
  NAND2_X1 U805 ( .A1(n876), .A2(n728), .ZN(n989) );
  NAND2_X1 U806 ( .A1(n729), .A2(n989), .ZN(n731) );
  AND2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n750) );
  NOR2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U809 ( .A1(n750), .A2(n734), .ZN(n753) );
  NAND2_X1 U810 ( .A1(n1000), .A2(KEYINPUT33), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n736), .A2(n745), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n528), .A2(n738), .ZN(n755) );
  NOR2_X1 U813 ( .A1(G2090), .A2(G303), .ZN(n740) );
  NAND2_X1 U814 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n739), .A2(n741), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n742), .A2(n745), .ZN(n747) );
  NOR2_X1 U817 ( .A1(G1981), .A2(G305), .ZN(n743) );
  XOR2_X1 U818 ( .A(n743), .B(KEYINPUT24), .Z(n744) );
  OR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n751) );
  OR2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U823 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U825 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U826 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U828 ( .A1(n884), .A2(G123), .ZN(n757) );
  XNOR2_X1 U829 ( .A(n757), .B(KEYINPUT18), .ZN(n759) );
  NAND2_X1 U830 ( .A1(G111), .A2(n690), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U832 ( .A1(G135), .A2(n888), .ZN(n761) );
  NAND2_X1 U833 ( .A1(G99), .A2(n891), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U835 ( .A1(n763), .A2(n762), .ZN(n977) );
  XNOR2_X1 U836 ( .A(n977), .B(G2096), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n764), .B(KEYINPUT79), .ZN(n765) );
  OR2_X1 U838 ( .A1(G2100), .A2(n765), .ZN(G156) );
  INV_X1 U839 ( .A(G132), .ZN(G219) );
  INV_X1 U840 ( .A(G82), .ZN(G220) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  INV_X1 U842 ( .A(G171), .ZN(G301) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n766) );
  XOR2_X1 U844 ( .A(n766), .B(KEYINPUT10), .Z(n919) );
  NAND2_X1 U845 ( .A1(n919), .A2(G567), .ZN(n767) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  INV_X1 U847 ( .A(n779), .ZN(n1003) );
  NAND2_X1 U848 ( .A1(n1003), .A2(G860), .ZN(n768) );
  XOR2_X1 U849 ( .A(KEYINPUT73), .B(n768), .Z(G153) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U851 ( .A(G868), .ZN(n809) );
  NAND2_X1 U852 ( .A1(n769), .A2(n809), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n771), .A2(n770), .ZN(G284) );
  INV_X1 U854 ( .A(n1007), .ZN(G299) );
  NOR2_X1 U855 ( .A1(G286), .A2(n809), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G868), .A2(G299), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U858 ( .A(KEYINPUT76), .B(n774), .ZN(G297) );
  INV_X1 U859 ( .A(G559), .ZN(n775) );
  NOR2_X1 U860 ( .A1(G860), .A2(n775), .ZN(n776) );
  XNOR2_X1 U861 ( .A(KEYINPUT77), .B(n776), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n777), .A2(n1006), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U864 ( .A1(G868), .A2(n779), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G868), .A2(n1006), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U868 ( .A(KEYINPUT78), .B(n783), .ZN(G282) );
  NAND2_X1 U869 ( .A1(n784), .A2(G80), .ZN(n787) );
  NAND2_X1 U870 ( .A1(G67), .A2(n785), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U872 ( .A1(G93), .A2(n788), .ZN(n789) );
  XNOR2_X1 U873 ( .A(KEYINPUT81), .B(n789), .ZN(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U875 ( .A1(n792), .A2(G55), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n794), .A2(n793), .ZN(n808) );
  XOR2_X1 U877 ( .A(n1003), .B(KEYINPUT80), .Z(n796) );
  NAND2_X1 U878 ( .A1(n1006), .A2(G559), .ZN(n795) );
  XNOR2_X1 U879 ( .A(n796), .B(n795), .ZN(n806) );
  NOR2_X1 U880 ( .A1(n806), .A2(G860), .ZN(n797) );
  XOR2_X1 U881 ( .A(n808), .B(n797), .Z(G145) );
  XOR2_X1 U882 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n799) );
  XNOR2_X1 U883 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U885 ( .A(G305), .B(n800), .ZN(n802) );
  XOR2_X1 U886 ( .A(G299), .B(G166), .Z(n801) );
  XNOR2_X1 U887 ( .A(n802), .B(n801), .ZN(n803) );
  XOR2_X1 U888 ( .A(n803), .B(G288), .Z(n804) );
  XNOR2_X1 U889 ( .A(n808), .B(n804), .ZN(n805) );
  XNOR2_X1 U890 ( .A(G290), .B(n805), .ZN(n900) );
  XNOR2_X1 U891 ( .A(n900), .B(n806), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n807), .A2(G868), .ZN(n811) );
  NAND2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U895 ( .A(KEYINPUT89), .B(n812), .Z(G295) );
  XOR2_X1 U896 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n814) );
  NAND2_X1 U897 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n815), .ZN(n816) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n816), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n817), .A2(G2072), .ZN(G158) );
  NAND2_X1 U902 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U903 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G108), .A2(n819), .ZN(n831) );
  NAND2_X1 U905 ( .A1(G567), .A2(n831), .ZN(n820) );
  XNOR2_X1 U906 ( .A(n820), .B(KEYINPUT91), .ZN(n825) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n821) );
  XNOR2_X1 U908 ( .A(KEYINPUT22), .B(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n822), .A2(G96), .ZN(n823) );
  OR2_X1 U910 ( .A1(G218), .A2(n823), .ZN(n832) );
  AND2_X1 U911 ( .A1(G2106), .A2(n832), .ZN(n824) );
  NOR2_X1 U912 ( .A1(n825), .A2(n824), .ZN(G319) );
  INV_X1 U913 ( .A(G319), .ZN(n827) );
  NAND2_X1 U914 ( .A1(G661), .A2(G483), .ZN(n826) );
  NOR2_X1 U915 ( .A1(n827), .A2(n826), .ZN(n830) );
  NAND2_X1 U916 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n919), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(G2084), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2078), .B(G2072), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U931 ( .A(n835), .B(G2100), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U934 ( .A(G2096), .B(G2678), .Z(n839) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U937 ( .A(n841), .B(n840), .Z(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT107), .B(G1976), .Z(n844) );
  XOR2_X1 U939 ( .A(n842), .B(G1981), .Z(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U941 ( .A(n845), .B(KEYINPUT41), .Z(n848) );
  INV_X1 U942 ( .A(G1996), .ZN(n846) );
  XOR2_X1 U943 ( .A(n846), .B(G1991), .Z(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n852) );
  XNOR2_X1 U945 ( .A(G1971), .B(n997), .ZN(n850) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U948 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U949 ( .A(G2474), .B(KEYINPUT106), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G124), .A2(n884), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n855), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G136), .A2(n888), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n856), .B(KEYINPUT108), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U956 ( .A1(G100), .A2(n891), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G112), .A2(n690), .ZN(n859) );
  NAND2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U959 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n874) );
  NAND2_X1 U963 ( .A1(G130), .A2(n884), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G118), .A2(n690), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U966 ( .A1(n891), .A2(G106), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT109), .B(n867), .Z(n869) );
  NAND2_X1 U968 ( .A1(n888), .A2(G142), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n870), .B(KEYINPUT45), .Z(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n875) );
  XOR2_X1 U973 ( .A(n875), .B(G162), .Z(n878) );
  XOR2_X1 U974 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n977), .B(n879), .ZN(n883) );
  XOR2_X1 U977 ( .A(n881), .B(n880), .Z(n882) );
  XNOR2_X1 U978 ( .A(n883), .B(n882), .ZN(n896) );
  NAND2_X1 U979 ( .A1(G127), .A2(n884), .ZN(n886) );
  NAND2_X1 U980 ( .A1(G115), .A2(n690), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n887), .B(KEYINPUT47), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G139), .A2(n888), .ZN(n889) );
  NAND2_X1 U984 ( .A1(n890), .A2(n889), .ZN(n894) );
  NAND2_X1 U985 ( .A1(G103), .A2(n891), .ZN(n892) );
  XNOR2_X1 U986 ( .A(KEYINPUT111), .B(n892), .ZN(n893) );
  NOR2_X1 U987 ( .A1(n894), .A2(n893), .ZN(n968) );
  XOR2_X1 U988 ( .A(G160), .B(n968), .Z(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U991 ( .A(n1003), .B(G286), .Z(n899) );
  XOR2_X1 U992 ( .A(G301), .B(n1006), .Z(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U994 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U995 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2438), .B(KEYINPUT104), .Z(n904) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2430), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(n905), .B(G2435), .Z(n907) );
  XNOR2_X1 U1000 ( .A(G1348), .B(G1341), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2427), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2446), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n918), .ZN(G401) );
  INV_X1 U1016 ( .A(n919), .ZN(G223) );
  XOR2_X1 U1017 ( .A(G5), .B(G1961), .Z(n940) );
  XOR2_X1 U1018 ( .A(G4), .B(KEYINPUT124), .Z(n921) );
  XNOR2_X1 U1019 ( .A(G1348), .B(KEYINPUT59), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n921), .B(n920), .ZN(n928) );
  XOR2_X1 U1021 ( .A(G1341), .B(G19), .Z(n923) );
  XOR2_X1 U1022 ( .A(G1956), .B(G20), .Z(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G6), .B(G1981), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT123), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n929), .B(KEYINPUT60), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT125), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(G1986), .B(G24), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1033 ( .A(G1976), .B(KEYINPUT126), .Z(n933) );
  XNOR2_X1 U1034 ( .A(G23), .B(n933), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT58), .B(n936), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(G21), .B(G1966), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(KEYINPUT61), .B(n943), .ZN(n944) );
  INV_X1 U1042 ( .A(G16), .ZN(n1024) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n1024), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n945), .A2(G11), .ZN(n996) );
  XNOR2_X1 U1045 ( .A(KEYINPUT54), .B(G34), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(n946), .B(KEYINPUT118), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G2084), .B(n947), .ZN(n965) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(KEYINPUT116), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(KEYINPUT115), .B(G2067), .ZN(n948) );
  XNOR2_X1 U1050 ( .A(n948), .B(G26), .ZN(n955) );
  XOR2_X1 U1051 ( .A(G1991), .B(G25), .Z(n950) );
  XOR2_X1 U1052 ( .A(G1996), .B(G32), .Z(n949) );
  NAND2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1054 ( .A(G27), .B(n951), .Z(n952) );
  NOR2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1057 ( .A(G2072), .B(G33), .Z(n956) );
  NAND2_X1 U1058 ( .A1(G28), .A2(n956), .ZN(n957) );
  NOR2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1060 ( .A(n960), .B(n959), .ZN(n962) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1063 ( .A(KEYINPUT117), .B(n963), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(G29), .A2(n966), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(n967), .B(KEYINPUT55), .ZN(n994) );
  XOR2_X1 U1067 ( .A(G2072), .B(n968), .Z(n970) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n969) );
  NOR2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1070 ( .A(KEYINPUT114), .B(n971), .ZN(n972) );
  XNOR2_X1 U1071 ( .A(n972), .B(KEYINPUT50), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1073 ( .A(G160), .B(G2084), .Z(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(KEYINPUT113), .B(n981), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n988) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(KEYINPUT51), .B(n986), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT52), .B(n991), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(G29), .A2(n992), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1029) );
  XOR2_X1 U1088 ( .A(n997), .B(G301), .Z(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1016) );
  INV_X1 U1090 ( .A(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1092 ( .A(G1341), .B(n1003), .Z(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(n1006), .B(G1348), .Z(n1009) );
  XOR2_X1 U1095 ( .A(n1007), .B(G1956), .Z(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G166), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT121), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G168), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(n1019), .B(KEYINPUT57), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1024), .B(KEYINPUT56), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT122), .B(n1027), .Z(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(n1030), .B(KEYINPUT62), .ZN(n1031) );
  XOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1031), .Z(G150) );
  INV_X1 U1114 ( .A(G150), .ZN(G311) );
endmodule

