//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT0), .A4(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT0), .A4(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(new_n200), .B2(G146), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n198), .A2(KEYINPUT64), .A3(G143), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n199), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT65), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n200), .A2(G146), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n198), .B2(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n200), .A3(G146), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n218), .A2(new_n219), .A3(new_n212), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n197), .B(new_n207), .C1(new_n214), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n227), .B2(G119), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT68), .A3(G116), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n228), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n228), .A3(new_n232), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT69), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n230), .A2(new_n232), .A3(new_n237), .A4(new_n228), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n226), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n191), .A2(G134), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n188), .A2(G137), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n196), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n199), .A2(new_n201), .A3(new_n246), .A4(G128), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n218), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n221), .A2(new_n241), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT28), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n245), .A2(new_n250), .A3(KEYINPUT70), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT70), .B1(new_n245), .B2(new_n250), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n221), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n241), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n254), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n241), .A3(new_n221), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n253), .B1(new_n264), .B2(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G210), .ZN(new_n268));
  INV_X1    g082(.A(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(KEYINPUT29), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n263), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n257), .A2(KEYINPUT30), .ZN(new_n277));
  AND4_X1   g091(.A1(new_n246), .A2(new_n199), .A3(new_n201), .A4(G128), .ZN(new_n278));
  INV_X1    g092(.A(new_n249), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n211), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n196), .A2(new_n244), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT67), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n245), .A2(new_n250), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n221), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(KEYINPUT30), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n276), .B1(new_n286), .B2(new_n258), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n287), .B2(new_n272), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(KEYINPUT71), .A3(new_n258), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n263), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT71), .B1(new_n285), .B2(new_n258), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n253), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT73), .A4(new_n272), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT30), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n262), .B2(new_n221), .ZN(new_n296));
  AND4_X1   g110(.A1(new_n295), .A2(new_n221), .A3(new_n282), .A4(new_n284), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n258), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n263), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n300));
  INV_X1    g114(.A(new_n272), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n288), .A2(new_n294), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n292), .A2(new_n293), .A3(new_n272), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n275), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G472), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT75), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n298), .A2(new_n263), .A3(new_n272), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n298), .A2(KEYINPUT31), .A3(new_n263), .A4(new_n272), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n292), .A2(new_n293), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(new_n301), .ZN(new_n315));
  NOR2_X1   g129(.A1(G472), .A2(G902), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT72), .ZN(new_n317));
  OR3_X1    g131(.A1(new_n315), .A2(KEYINPUT32), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT32), .B1(new_n315), .B2(new_n317), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n304), .A2(new_n305), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n288), .A2(new_n294), .A3(new_n302), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n321), .B(G472), .C1(new_n326), .C2(new_n275), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n309), .A2(new_n320), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n231), .A2(G128), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n329), .A2(KEYINPUT23), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n248), .A2(G119), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(KEYINPUT23), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n331), .A2(new_n329), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT24), .B(G110), .Z(new_n336));
  OAI22_X1  g150(.A1(new_n334), .A2(G110), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n338), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  XNOR2_X1  g153(.A(G125), .B(G140), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G146), .ZN(new_n342));
  INV_X1    g156(.A(new_n340), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n337), .B(new_n342), .C1(G146), .C2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n341), .B(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n334), .A2(G110), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n335), .A2(new_n336), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT76), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n352), .B2(new_n349), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT25), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n356), .A2(KEYINPUT25), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n355), .A2(new_n274), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G217), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(G234), .B2(new_n274), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n349), .A2(new_n352), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n349), .B2(new_n353), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n356), .B(KEYINPUT25), .C1(new_n363), .C2(G902), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n361), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n355), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT78), .Z(new_n369));
  NAND2_X1  g183(.A1(new_n328), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(G110), .B(G140), .ZN(new_n371));
  INV_X1    g185(.A(G227), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G953), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n371), .B(new_n373), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT80), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n382), .A2(new_n386), .A3(new_n383), .A4(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(G101), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n377), .A2(new_n380), .A3(new_n269), .A4(new_n381), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT4), .A4(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT79), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n388), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n211), .A2(KEYINPUT65), .A3(new_n213), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n219), .B1(new_n218), .B2(new_n212), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n396), .A2(new_n397), .B1(new_n203), .B2(new_n206), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n379), .A2(G104), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n376), .A2(G107), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n391), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n391), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n250), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT10), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n407), .A2(G128), .B1(new_n199), .B2(new_n201), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n391), .B(new_n401), .C1(new_n278), .C2(new_n408), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(KEYINPUT10), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n395), .A2(new_n398), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n197), .B(KEYINPUT82), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n375), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n197), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n391), .A2(new_n401), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n247), .B1(new_n249), .B2(new_n204), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n280), .A2(new_n416), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n414), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n280), .A2(new_n415), .A3(new_n416), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT12), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n409), .B(KEYINPUT83), .C1(new_n250), .C2(new_n417), .ZN(new_n424));
  AND4_X1   g238(.A1(KEYINPUT12), .A2(new_n424), .A3(new_n197), .A4(new_n422), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT84), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n197), .A3(new_n422), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n421), .A2(KEYINPUT12), .A3(new_n422), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n413), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT85), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n411), .A2(new_n412), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n414), .B2(new_n411), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n375), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n413), .A2(new_n426), .A3(new_n438), .A4(new_n432), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n274), .ZN(new_n442));
  NAND2_X1  g256(.A1(G469), .A2(G902), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n413), .B1(new_n414), .B2(new_n411), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n411), .A2(new_n412), .B1(new_n429), .B2(new_n430), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n374), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n442), .B(new_n443), .C1(new_n441), .C2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT9), .B(G234), .ZN(new_n448));
  OAI21_X1  g262(.A(G221), .B1(new_n448), .B2(G902), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT86), .B1(new_n398), .B2(new_n338), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n207), .B1(new_n214), .B2(new_n220), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(G125), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n280), .A2(KEYINPUT87), .A3(new_n338), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n250), .B2(G125), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n453), .A2(new_n456), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G224), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(new_n461), .B2(G953), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT8), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n236), .A2(KEYINPUT5), .A3(new_n238), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n227), .A2(G119), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n222), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n234), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n417), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT5), .A4(new_n228), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n233), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT88), .B1(new_n474), .B2(new_n416), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n417), .A2(new_n476), .A3(new_n233), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n465), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n395), .A2(new_n258), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n470), .B1(new_n404), .B2(new_n403), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n464), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT89), .B(new_n465), .C1(new_n471), .C2(new_n478), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n463), .A2(new_n481), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n460), .A2(new_n462), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n274), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT90), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n482), .A2(new_n483), .ZN(new_n490));
  INV_X1    g304(.A(new_n464), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n461), .A2(G953), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n460), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n496), .A3(new_n491), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n274), .C1(new_n486), .C2(new_n487), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n489), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n489), .A2(new_n502), .A3(new_n498), .A4(new_n500), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n452), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT94), .B(G122), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n227), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n508), .A2(G107), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n508), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n509), .B2(G116), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n227), .A3(G122), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT96), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n515), .A2(KEYINPUT96), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n512), .A2(new_n513), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n511), .B1(new_n518), .B2(G107), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n248), .A2(G143), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(G128), .B2(new_n200), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n248), .A2(KEYINPUT95), .A3(G143), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(G134), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n508), .A2(G107), .A3(new_n510), .ZN(new_n526));
  OAI21_X1  g340(.A(G107), .B1(new_n508), .B2(new_n510), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n200), .A2(G128), .ZN(new_n529));
  OAI21_X1  g343(.A(G134), .B1(new_n529), .B2(KEYINPUT13), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n524), .B(new_n530), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n519), .A2(new_n525), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n448), .A2(new_n360), .A3(G953), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT97), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n517), .A2(new_n516), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n513), .B1(new_n507), .B2(new_n227), .ZN(new_n538));
  OAI21_X1  g352(.A(G107), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n525), .A2(new_n526), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n542));
  INV_X1    g356(.A(new_n533), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n534), .A2(new_n535), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n274), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n546), .B(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G113), .B(G122), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n376), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n266), .A2(new_n267), .A3(G214), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(new_n200), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n200), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n195), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n195), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT92), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT19), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n343), .A2(KEYINPUT93), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT93), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n560), .A2(KEYINPUT93), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n340), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n198), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n553), .B(new_n200), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G131), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n556), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n559), .A2(new_n342), .A3(new_n566), .A4(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT18), .A3(G131), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n567), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n340), .B(new_n198), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n552), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n568), .A2(new_n578), .A3(new_n556), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n341), .B(new_n198), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n558), .A2(KEYINPUT17), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n576), .A2(new_n582), .A3(new_n552), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G475), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n585), .A4(new_n274), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n552), .B1(new_n576), .B2(new_n582), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n274), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G475), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n585), .B(new_n274), .C1(new_n577), .C2(new_n583), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n267), .A2(G952), .ZN(new_n594));
  NAND2_X1  g408(.A1(G234), .A2(G237), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT21), .B(G898), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(G902), .A3(G953), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n550), .A2(new_n593), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n450), .A2(new_n506), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n370), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(new_n269), .ZN(G3));
  NAND2_X1  g420(.A1(new_n312), .A2(new_n313), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n314), .A2(new_n301), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n308), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n315), .A2(new_n317), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n369), .A2(new_n450), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n504), .A2(new_n505), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n451), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n534), .A2(new_n616), .A3(new_n535), .A4(new_n544), .ZN(new_n617));
  AOI211_X1 g431(.A(KEYINPUT98), .B(new_n533), .C1(new_n536), .C2(new_n540), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n541), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT33), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(G478), .A3(new_n274), .ZN(new_n623));
  AOI21_X1  g437(.A(G478), .B1(new_n545), .B2(new_n274), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n593), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n602), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n615), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NOR2_X1   g449(.A1(new_n549), .A2(new_n593), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n630), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT99), .Z(new_n638));
  NAND3_X1  g452(.A1(new_n613), .A2(new_n506), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NAND4_X1  g455(.A1(new_n450), .A2(new_n506), .A3(new_n603), .A4(new_n612), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n353), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n349), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n366), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n365), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT100), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n652));
  INV_X1    g466(.A(new_n648), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n328), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n596), .B1(new_n600), .B2(G900), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n549), .A2(new_n593), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n450), .A2(new_n506), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n652), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n449), .A2(new_n506), .A3(new_n447), .A4(new_n657), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(KEYINPUT101), .A3(new_n328), .A4(new_n653), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(new_n655), .B(KEYINPUT39), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n450), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n647), .B1(new_n665), .B2(KEYINPUT40), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n287), .A2(new_n301), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n274), .B1(new_n264), .B2(new_n272), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n320), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n550), .A2(new_n593), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n671), .A2(new_n452), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n614), .B(KEYINPUT38), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n666), .A2(new_n667), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  AND4_X1   g490(.A1(new_n449), .A2(new_n614), .A3(new_n447), .A4(new_n451), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n547), .B(G902), .C1(new_n617), .C2(new_n621), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n593), .B(new_n655), .C1(new_n678), .C2(new_n624), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n677), .A2(new_n328), .A3(new_n680), .A4(new_n653), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  AND3_X1   g496(.A1(new_n440), .A2(new_n441), .A3(new_n274), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n441), .B1(new_n440), .B2(new_n274), .ZN(new_n684));
  INV_X1    g498(.A(new_n449), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n506), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n631), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n328), .A3(new_n369), .A4(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  AND3_X1   g507(.A1(new_n687), .A2(new_n328), .A3(new_n369), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n638), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n506), .A2(new_n686), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n506), .B2(new_n686), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n654), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n603), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND4_X1  g517(.A1(new_n506), .A2(new_n686), .A3(new_n593), .A4(new_n550), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n609), .B2(new_n308), .ZN(new_n706));
  OAI211_X1 g520(.A(KEYINPUT104), .B(G472), .C1(new_n315), .C2(G902), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n607), .B1(new_n272), .B2(new_n265), .ZN(new_n709));
  INV_X1    g523(.A(new_n317), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n368), .A3(new_n630), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  OR3_X1    g527(.A1(new_n704), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n713), .B1(new_n704), .B2(new_n712), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n679), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n626), .A2(KEYINPUT106), .A3(new_n593), .A4(new_n655), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n647), .A2(new_n708), .A3(new_n711), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n698), .B2(new_n699), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  AND2_X1   g538(.A1(new_n328), .A2(new_n369), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT108), .B1(new_n614), .B2(new_n452), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n504), .A2(new_n727), .A3(new_n451), .A4(new_n505), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n442), .A2(new_n443), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  OR3_X1    g544(.A1(new_n445), .A2(new_n730), .A3(new_n374), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n445), .B2(new_n374), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n444), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(new_n441), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n685), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n726), .A2(new_n728), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT42), .B1(new_n719), .B2(new_n720), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n725), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n328), .A2(new_n368), .A3(new_n721), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n726), .A2(new_n728), .A3(new_n735), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT42), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND3_X1  g557(.A1(new_n725), .A2(new_n736), .A3(new_n657), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  NOR2_X1   g559(.A1(new_n627), .A2(new_n593), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT43), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n747), .B(new_n647), .C1(new_n611), .C2(new_n610), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT44), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n726), .A2(new_n728), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n446), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(G469), .B(new_n752), .C1(new_n733), .C2(new_n751), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(new_n443), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n442), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(new_n449), .A3(new_n664), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n749), .A2(new_n750), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT109), .B(G137), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G39));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n449), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT110), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n757), .A2(new_n764), .A3(new_n449), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n763), .A2(new_n765), .B1(KEYINPUT111), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n328), .A2(new_n369), .A3(new_n679), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n750), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  NOR2_X1   g588(.A1(new_n683), .A2(new_n684), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n671), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n746), .A2(new_n368), .A3(new_n449), .A4(new_n451), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n775), .B1(KEYINPUT112), .B2(new_n780), .ZN(new_n781));
  OR4_X1    g595(.A1(new_n674), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n783));
  AND2_X1   g597(.A1(new_n750), .A2(new_n686), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n369), .A2(new_n784), .A3(new_n597), .A4(new_n671), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n628), .A3(new_n627), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT120), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT120), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n747), .A2(new_n597), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n708), .A2(new_n711), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n368), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n674), .A2(new_n451), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n686), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n789), .A2(new_n790), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n787), .A2(new_n788), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n784), .A2(new_n647), .A3(new_n793), .A4(new_n792), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n775), .A2(new_n685), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n768), .B2(new_n770), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n794), .A2(new_n750), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n783), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n785), .A2(new_n629), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n368), .A2(new_n784), .A3(new_n328), .A4(new_n792), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n807), .B(new_n594), .C1(KEYINPUT48), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(KEYINPUT48), .B2(new_n808), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n803), .A2(KEYINPUT121), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n803), .A2(KEYINPUT121), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n804), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT51), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n806), .B(new_n810), .C1(new_n801), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n370), .A2(new_n604), .B1(new_n642), .B2(new_n648), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n632), .A2(KEYINPUT113), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n615), .B2(new_n631), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n818), .B(new_n820), .C1(new_n615), .C2(new_n637), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n821), .B2(new_n613), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n714), .A2(new_n715), .B1(new_n694), .B2(new_n638), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n691), .A3(new_n702), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n593), .A2(new_n656), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n750), .A2(KEYINPUT114), .A3(new_n549), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n726), .A2(new_n549), .A3(new_n825), .A4(new_n728), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n450), .A3(new_n701), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n736), .A2(new_n722), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n742), .A2(new_n830), .A3(new_n744), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n723), .A2(new_n681), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n671), .A2(new_n647), .A3(new_n656), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n615), .A2(new_n672), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n735), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n662), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n835), .A2(new_n662), .A3(KEYINPUT52), .A4(new_n838), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n839), .A2(KEYINPUT115), .A3(new_n840), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n833), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n841), .A2(new_n849), .A3(new_n843), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n841), .B2(new_n843), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n848), .B(new_n833), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n833), .A2(new_n844), .A3(new_n848), .A4(new_n845), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n691), .A2(new_n823), .A3(new_n702), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n738), .A2(new_n744), .A3(new_n741), .A4(new_n831), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n829), .A2(new_n701), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n450), .B1(new_n827), .B2(new_n828), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n862), .A3(new_n822), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n834), .B1(new_n659), .B2(new_n661), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n864), .B2(new_n838), .ZN(new_n865));
  AND4_X1   g679(.A1(KEYINPUT52), .A2(new_n835), .A3(new_n662), .A4(new_n838), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT116), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n841), .A2(new_n849), .A3(new_n843), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(KEYINPUT54), .B(new_n856), .C1(new_n869), .C2(new_n848), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n816), .B1(new_n855), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n816), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n794), .A2(new_n700), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n815), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(G952), .A2(G953), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n782), .B1(new_n875), .B2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n853), .A2(new_n274), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n493), .A2(new_n497), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n495), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n882), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n267), .A2(G952), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G51));
  AND2_X1   g700(.A1(new_n847), .A2(new_n852), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n855), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n443), .B(KEYINPUT57), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n440), .B(KEYINPUT122), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n853), .A2(new_n274), .A3(new_n753), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(G54));
  NAND3_X1  g709(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(new_n584), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n885), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n889), .A2(new_n622), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n885), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n905));
  INV_X1    g719(.A(new_n870), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n847), .B2(new_n852), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT117), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n900), .B1(new_n908), .B2(new_n872), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n622), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n901), .B1(new_n871), .B2(new_n873), .ZN(new_n911));
  INV_X1    g725(.A(new_n622), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(KEYINPUT123), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n910), .B2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT60), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n887), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n885), .B1(new_n917), .B2(new_n363), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n887), .A2(new_n645), .A3(new_n916), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n919), .B(new_n920), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n917), .A2(new_n363), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n917), .A2(KEYINPUT125), .A3(new_n363), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n926), .A2(new_n903), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n925), .A2(new_n931), .ZN(G66));
  OAI21_X1  g746(.A(G953), .B1(new_n599), .B2(new_n461), .ZN(new_n933));
  INV_X1    g747(.A(new_n824), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n880), .B1(G898), .B2(new_n267), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(G69));
  XOR2_X1   g751(.A(new_n286), .B(new_n565), .Z(new_n938));
  AND2_X1   g752(.A1(new_n773), .A2(new_n759), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n758), .A2(new_n368), .A3(new_n328), .A4(new_n837), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n742), .A2(new_n744), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT126), .Z(new_n942));
  NAND4_X1  g756(.A1(new_n939), .A2(new_n864), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n943), .B2(new_n267), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n372), .A2(G900), .A3(G953), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n864), .A2(new_n675), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  AND3_X1   g763(.A1(new_n750), .A2(new_n450), .A3(new_n664), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(new_n725), .C1(new_n629), .C2(new_n636), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n939), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n947), .B(new_n938), .C1(new_n952), .C2(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n946), .A2(new_n953), .ZN(G72));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n952), .B2(new_n824), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n885), .B1(new_n957), .B2(new_n668), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n943), .B2(new_n824), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n301), .A3(new_n287), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n288), .A2(new_n310), .A3(new_n302), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(new_n956), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n856), .B(new_n962), .C1(new_n869), .C2(new_n848), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n958), .A2(new_n960), .A3(new_n963), .ZN(G57));
endmodule


