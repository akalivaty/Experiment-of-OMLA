

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  NOR2_X2 U321 ( .A1(n457), .A2(n456), .ZN(n561) );
  XOR2_X1 U322 ( .A(n432), .B(n431), .Z(n522) );
  XNOR2_X1 U323 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U324 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U325 ( .A(n367), .B(n366), .Z(n572) );
  XNOR2_X1 U326 ( .A(n572), .B(KEYINPUT41), .ZN(n550) );
  XOR2_X1 U327 ( .A(n308), .B(n307), .Z(n531) );
  XNOR2_X1 U328 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U329 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n290) );
  XNOR2_X1 U331 ( .A(KEYINPUT89), .B(KEYINPUT20), .ZN(n289) );
  XNOR2_X1 U332 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U333 ( .A(n291), .B(G176GAT), .Z(n293) );
  XOR2_X1 U334 ( .A(G15GAT), .B(G127GAT), .Z(n376) );
  XNOR2_X1 U335 ( .A(n376), .B(KEYINPUT87), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n298) );
  XNOR2_X1 U337 ( .A(G99GAT), .B(G71GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n294), .B(G120GAT), .ZN(n363) );
  XOR2_X1 U339 ( .A(G43GAT), .B(G134GAT), .Z(n399) );
  XOR2_X1 U340 ( .A(n363), .B(n399), .Z(n296) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U343 ( .A(n298), .B(n297), .Z(n308) );
  XOR2_X1 U344 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n300) );
  XNOR2_X1 U345 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U347 ( .A(G113GAT), .B(n301), .Z(n317) );
  XOR2_X1 U348 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n303) );
  XNOR2_X1 U349 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U351 ( .A(n304), .B(KEYINPUT19), .Z(n306) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n432) );
  XNOR2_X1 U354 ( .A(n317), .B(n432), .ZN(n307) );
  INV_X1 U355 ( .A(n531), .ZN(n457) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U357 ( .A(KEYINPUT78), .B(G85GAT), .Z(n310) );
  XNOR2_X1 U358 ( .A(G162GAT), .B(G155GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n312) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G134GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n329) );
  XOR2_X1 U363 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n319) );
  XOR2_X1 U364 ( .A(KEYINPUT3), .B(KEYINPUT95), .Z(n316) );
  XNOR2_X1 U365 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n443) );
  XNOR2_X1 U367 ( .A(n317), .B(n443), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n327) );
  XOR2_X1 U369 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n321) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U372 ( .A(G57GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U373 ( .A(G120GAT), .B(G127GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U375 ( .A(n325), .B(n324), .Z(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U377 ( .A(n329), .B(n328), .Z(n473) );
  INV_X1 U378 ( .A(n473), .ZN(n519) );
  INV_X1 U379 ( .A(KEYINPUT54), .ZN(n434) );
  XOR2_X1 U380 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n369) );
  XOR2_X1 U381 ( .A(G113GAT), .B(G197GAT), .Z(n331) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(G141GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(n332), .B(G50GAT), .Z(n334) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G8GAT), .Z(n421) );
  XNOR2_X1 U386 ( .A(n421), .B(G43GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n339) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n335), .B(KEYINPUT7), .ZN(n404) );
  XOR2_X1 U390 ( .A(n404), .B(KEYINPUT67), .Z(n337) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U393 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U394 ( .A(KEYINPUT66), .B(KEYINPUT69), .Z(n341) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G15GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U397 ( .A(G1GAT), .B(KEYINPUT68), .Z(n343) );
  XNOR2_X1 U398 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U401 ( .A(n347), .B(n346), .Z(n507) );
  INV_X1 U402 ( .A(n507), .ZN(n569) );
  XNOR2_X1 U403 ( .A(G85GAT), .B(G92GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n348), .B(KEYINPUT73), .ZN(n400) );
  XOR2_X1 U405 ( .A(KEYINPUT71), .B(n400), .Z(n350) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n367) );
  XOR2_X1 U408 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n352) );
  XNOR2_X1 U409 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n354) );
  INV_X1 U411 ( .A(KEYINPUT76), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U413 ( .A(G176GAT), .B(G64GAT), .Z(n422) );
  XNOR2_X1 U414 ( .A(n422), .B(KEYINPUT31), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n358) );
  XNOR2_X1 U416 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n357), .B(KEYINPUT13), .ZN(n379) );
  XNOR2_X1 U418 ( .A(n358), .B(n379), .ZN(n365) );
  INV_X1 U419 ( .A(KEYINPUT72), .ZN(n362) );
  XOR2_X1 U420 ( .A(G148GAT), .B(G106GAT), .Z(n360) );
  XNOR2_X1 U421 ( .A(G204GAT), .B(G78GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n449) );
  XOR2_X1 U424 ( .A(n363), .B(n449), .Z(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  NAND2_X1 U426 ( .A1(n569), .A2(n550), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n388) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U429 ( .A(G1GAT), .B(G8GAT), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n373) );
  XNOR2_X1 U432 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n387) );
  XOR2_X1 U435 ( .A(G22GAT), .B(G155GAT), .Z(n439) );
  XOR2_X1 U436 ( .A(n439), .B(G211GAT), .Z(n378) );
  XNOR2_X1 U437 ( .A(n376), .B(G78GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U439 ( .A(n379), .B(KEYINPUT12), .Z(n381) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U442 ( .A(n383), .B(n382), .Z(n385) );
  XNOR2_X1 U443 ( .A(G183GAT), .B(G71GAT), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U445 ( .A(n387), .B(n386), .Z(n490) );
  INV_X1 U446 ( .A(n490), .ZN(n575) );
  NOR2_X1 U447 ( .A1(n388), .A2(n575), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n389), .B(KEYINPUT115), .ZN(n409) );
  XOR2_X1 U449 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n391) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(G190GAT), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n393) );
  XNOR2_X1 U453 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U455 ( .A(G50GAT), .B(G162GAT), .Z(n442) );
  XOR2_X1 U456 ( .A(n394), .B(n442), .Z(n396) );
  XNOR2_X1 U457 ( .A(G99GAT), .B(G106GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n408) );
  XOR2_X1 U460 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U463 ( .A(n403), .B(KEYINPUT10), .Z(n406) );
  XNOR2_X1 U464 ( .A(n404), .B(KEYINPUT9), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n560) );
  NOR2_X1 U467 ( .A1(n409), .A2(n560), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n410), .B(KEYINPUT47), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n560), .B(KEYINPUT105), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n411), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U471 ( .A1(n580), .A2(n490), .ZN(n412) );
  XOR2_X1 U472 ( .A(KEYINPUT45), .B(n412), .Z(n413) );
  NOR2_X1 U473 ( .A1(n569), .A2(n413), .ZN(n414) );
  NAND2_X1 U474 ( .A1(n414), .A2(n572), .ZN(n415) );
  NAND2_X1 U475 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U476 ( .A(KEYINPUT48), .B(n417), .ZN(n530) );
  XOR2_X1 U477 ( .A(KEYINPUT98), .B(KEYINPUT79), .Z(n419) );
  NAND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n430) );
  XOR2_X1 U481 ( .A(n422), .B(G92GAT), .Z(n428) );
  XNOR2_X1 U482 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n423), .B(KEYINPUT93), .ZN(n424) );
  XOR2_X1 U484 ( .A(n424), .B(KEYINPUT94), .Z(n426) );
  XNOR2_X1 U485 ( .A(G197GAT), .B(G218GAT), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n448) );
  XNOR2_X1 U487 ( .A(G204GAT), .B(n448), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  AND2_X1 U490 ( .A1(n530), .A2(n522), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  NOR2_X1 U492 ( .A1(n519), .A2(n435), .ZN(n566) );
  XOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n437) );
  XNOR2_X1 U494 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U496 ( .A(n438), .B(KEYINPUT96), .Z(n441) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT92), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U500 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n469) );
  NAND2_X1 U505 ( .A1(n566), .A2(n469), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n453) );
  INV_X1 U507 ( .A(KEYINPUT55), .ZN(n452) );
  NAND2_X1 U508 ( .A1(n561), .A2(n550), .ZN(n461) );
  XOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n459) );
  XOR2_X1 U510 ( .A(G176GAT), .B(KEYINPUT123), .Z(n458) );
  NAND2_X1 U511 ( .A1(n569), .A2(n572), .ZN(n494) );
  NOR2_X1 U512 ( .A1(n560), .A2(n490), .ZN(n462) );
  XNOR2_X1 U513 ( .A(n462), .B(KEYINPUT16), .ZN(n477) );
  XOR2_X1 U514 ( .A(KEYINPUT90), .B(n531), .Z(n464) );
  XOR2_X1 U515 ( .A(n469), .B(KEYINPUT28), .Z(n525) );
  XNOR2_X1 U516 ( .A(KEYINPUT27), .B(KEYINPUT99), .ZN(n463) );
  XOR2_X1 U517 ( .A(n463), .B(n522), .Z(n467) );
  NAND2_X1 U518 ( .A1(n519), .A2(n467), .ZN(n547) );
  NOR2_X1 U519 ( .A1(n525), .A2(n547), .ZN(n532) );
  NAND2_X1 U520 ( .A1(n464), .A2(n532), .ZN(n476) );
  NOR2_X1 U521 ( .A1(n469), .A2(n531), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n567) );
  NAND2_X1 U524 ( .A1(n467), .A2(n567), .ZN(n472) );
  NAND2_X1 U525 ( .A1(n522), .A2(n531), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n470), .Z(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n489) );
  NAND2_X1 U531 ( .A1(n477), .A2(n489), .ZN(n508) );
  NOR2_X1 U532 ( .A1(n494), .A2(n508), .ZN(n487) );
  NAND2_X1 U533 ( .A1(n519), .A2(n487), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  XOR2_X1 U536 ( .A(G8GAT), .B(KEYINPUT101), .Z(n481) );
  NAND2_X1 U537 ( .A1(n487), .A2(n522), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n483) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT102), .B(n484), .Z(n486) );
  NAND2_X1 U543 ( .A1(n487), .A2(n531), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n487), .A2(n525), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U547 ( .A1(n490), .A2(n489), .ZN(n491) );
  NOR2_X1 U548 ( .A1(n580), .A2(n491), .ZN(n493) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(n518) );
  NOR2_X1 U551 ( .A1(n494), .A2(n518), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n495), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U553 ( .A1(n504), .A2(n519), .ZN(n498) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n504), .A2(n522), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n502) );
  NAND2_X1 U561 ( .A1(n504), .A2(n531), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n525), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  NAND2_X1 U568 ( .A1(n507), .A2(n550), .ZN(n517) );
  NOR2_X1 U569 ( .A1(n517), .A2(n508), .ZN(n513) );
  NAND2_X1 U570 ( .A1(n513), .A2(n519), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n513), .A2(n522), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n531), .A2(n513), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U577 ( .A1(n513), .A2(n525), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n526), .A2(n519), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n531), .A2(n526), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n528) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  INV_X1 U592 ( .A(n530), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U594 ( .A1(n545), .A2(n533), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n541), .A2(n569), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U599 ( .A1(n541), .A2(n550), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U602 ( .A1(n541), .A2(n575), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U606 ( .A1(n541), .A2(n560), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U610 ( .A1(n530), .A2(n567), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n556), .A2(n569), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n554) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U616 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n556), .A2(n575), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n560), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n561), .A2(n569), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n575), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n565) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT124), .B(n568), .ZN(n579) );
  INV_X1 U635 ( .A(n579), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n576), .A2(n569), .ZN(n570) );
  XOR2_X1 U637 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  OR2_X1 U639 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

