//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G119), .B(G128), .ZN(new_n194));
  INV_X1    g008(.A(G110), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT24), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G110), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n205), .A2(G146), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(G146), .B1(new_n205), .B2(new_n206), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n200), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n200), .B(KEYINPUT73), .C1(new_n207), .C2(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT74), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n205), .A2(new_n206), .A3(new_n216), .A4(G146), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(new_n204), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n190), .A2(G119), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n192), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n196), .A3(new_n198), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(KEYINPUT75), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n215), .A3(new_n217), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n213), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G137), .ZN(new_n231));
  INV_X1    g045(.A(G221), .ZN(new_n232));
  INV_X1    g046(.A(G234), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n232), .A2(new_n233), .A3(G953), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n231), .B(new_n234), .Z(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n213), .A2(new_n226), .A3(new_n229), .A4(new_n235), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT76), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT25), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n237), .A2(new_n238), .A3(new_n239), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(G217), .B1(new_n233), .B2(G902), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT72), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n237), .A2(new_n239), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n233), .B2(G217), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n246), .A2(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n256), .C2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT65), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n255), .A3(new_n257), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT64), .B(G131), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(G137), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n266), .A2(new_n269), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n268), .A2(G137), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n270), .A2(G134), .ZN(new_n275));
  OAI21_X1  g089(.A(G131), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n265), .A2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n280));
  OAI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(KEYINPUT2), .B2(G113), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n188), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G119), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n282), .B2(new_n284), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n286), .B1(new_n291), .B2(new_n281), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n273), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT0), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n190), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n258), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G143), .B(G146), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n296), .B2(new_n190), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  AND4_X1   g117(.A1(new_n253), .A2(new_n278), .A3(new_n292), .A4(new_n303), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n265), .A2(new_n277), .B1(new_n295), .B2(new_n302), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n253), .B1(new_n305), .B2(new_n292), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n281), .A2(new_n285), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n281), .A3(new_n288), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n278), .A2(new_n312), .A3(new_n303), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n278), .B2(new_n303), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G237), .ZN(new_n316));
  INV_X1    g130(.A(G953), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G210), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT27), .Z(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(KEYINPUT31), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n307), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n322), .A2(KEYINPUT31), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n325), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n307), .A2(new_n315), .A3(new_n323), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n278), .A2(new_n292), .A3(new_n303), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n278), .A2(new_n303), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n311), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n305), .A2(new_n253), .A3(new_n292), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT28), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n321), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n342));
  NOR2_X1   g156(.A1(G472), .A2(G902), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n326), .A2(new_n328), .B1(new_n339), .B2(new_n321), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT32), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n330), .A2(KEYINPUT70), .A3(new_n337), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT70), .B1(new_n330), .B2(new_n337), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n321), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(KEYINPUT29), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n336), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n238), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT71), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(KEYINPUT71), .A3(new_n238), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n307), .A2(new_n315), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n359), .B2(new_n321), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n339), .B2(new_n321), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G472), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n252), .B1(new_n348), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n316), .A2(new_n317), .A3(G143), .A4(G214), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n316), .A2(new_n317), .A3(G214), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT82), .A4(G214), .ZN(new_n371));
  AND4_X1   g185(.A1(KEYINPUT83), .A2(new_n370), .A3(new_n256), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(G143), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT83), .B1(new_n373), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n367), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT18), .A3(G131), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n367), .C1(new_n372), .C2(new_n374), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n219), .B(G146), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n266), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n207), .A2(new_n208), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(KEYINPUT85), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n381), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT17), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n367), .B(new_n266), .C1(new_n372), .C2(new_n374), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT85), .B1(new_n382), .B2(new_n383), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n380), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT86), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n380), .B(new_n395), .C1(new_n389), .C2(new_n390), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n238), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G475), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n391), .A2(new_n394), .ZN(new_n402));
  INV_X1    g216(.A(new_n394), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n380), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n385), .A2(new_n387), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n219), .B(KEYINPUT19), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n405), .B(new_n218), .C1(G146), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(G475), .A2(G902), .ZN(new_n409));
  AND4_X1   g223(.A1(new_n401), .A2(new_n402), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n391), .A2(new_n394), .B1(new_n407), .B2(new_n404), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n401), .B1(new_n411), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n400), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(KEYINPUT91), .A2(G952), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT91), .A2(G952), .ZN(new_n416));
  AOI21_X1  g230(.A(G953), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n233), .B2(new_n316), .ZN(new_n418));
  AOI211_X1 g232(.A(new_n238), .B(new_n317), .C1(G234), .C2(G237), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(G898), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n424));
  INV_X1    g238(.A(G122), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT87), .B1(new_n425), .B2(G116), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n283), .A3(G122), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G107), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(G116), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n190), .A2(G143), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n256), .A2(G128), .ZN(new_n436));
  AND2_X1   g250(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n437));
  OAI22_X1  g251(.A1(new_n256), .A2(G128), .B1(KEYINPUT88), .B2(KEYINPUT13), .ZN(new_n438));
  OAI221_X1 g252(.A(G134), .B1(new_n435), .B2(new_n436), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G134), .B1(new_n438), .B2(new_n437), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n435), .A2(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n429), .A2(KEYINPUT14), .B1(G116), .B2(new_n425), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n426), .A2(new_n428), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n430), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n441), .A2(G134), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n268), .B1(new_n435), .B2(new_n436), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n445), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n448), .A3(new_n431), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G107), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT89), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n444), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(G217), .A3(new_n317), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n424), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n459), .ZN(new_n466));
  INV_X1    g280(.A(new_n444), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n464), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n472), .A3(new_n238), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n470), .A2(new_n472), .A3(new_n238), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n413), .A2(new_n423), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n430), .A3(G104), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n393), .A2(G107), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G101), .ZN(new_n488));
  INV_X1    g302(.A(G101), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n485), .A3(new_n489), .A4(new_n486), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n487), .A2(new_n492), .A3(G101), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n311), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n430), .A2(G104), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n393), .A2(G107), .ZN(new_n496));
  OAI21_X1  g310(.A(G101), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT5), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n309), .B2(new_n288), .ZN(new_n500));
  OAI21_X1  g314(.A(G113), .B1(new_n282), .B2(KEYINPUT5), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n498), .B(new_n308), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G122), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n494), .A2(new_n502), .A3(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(KEYINPUT6), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n265), .A2(new_n203), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n302), .A2(G125), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G224), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(G953), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n515), .A3(new_n510), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n503), .A2(new_n518), .A3(new_n505), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n508), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n504), .B(KEYINPUT8), .Z(new_n525));
  NOR2_X1   g339(.A1(new_n285), .A2(new_n499), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n308), .B1(new_n501), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n525), .B1(new_n527), .B2(new_n498), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n308), .B1(new_n500), .B2(new_n501), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n498), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n509), .A2(new_n521), .A3(new_n515), .A4(new_n510), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n507), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n238), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n482), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n530), .A2(new_n507), .A3(new_n531), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n535), .B2(new_n523), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n508), .A2(new_n517), .A3(new_n519), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n481), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n538), .A3(KEYINPUT81), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(new_n482), .C1(new_n520), .C2(new_n533), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n264), .A2(KEYINPUT77), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT1), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(G143), .B2(new_n254), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n258), .B1(new_n546), .B2(new_n190), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n300), .A2(new_n548), .A3(new_n263), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n498), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n491), .A2(new_n302), .A3(new_n493), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n294), .A2(new_n273), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n490), .A2(new_n497), .A3(KEYINPUT10), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n265), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n490), .A2(new_n497), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n262), .A2(new_n559), .A3(new_n264), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT12), .B1(new_n561), .B2(new_n295), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n563), .B(new_n555), .C1(new_n551), .C2(new_n560), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n558), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n317), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n558), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n295), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G469), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT79), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n565), .A2(new_n568), .B1(new_n571), .B2(new_n573), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(G469), .C1(new_n579), .C2(G902), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n562), .A2(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n558), .A2(new_n570), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n570), .B1(new_n573), .B2(new_n558), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n576), .B(new_n238), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n587));
  INV_X1    g401(.A(new_n558), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n551), .A2(new_n552), .B1(new_n556), .B2(new_n265), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n555), .B1(new_n589), .B2(new_n554), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n568), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n558), .B(new_n570), .C1(new_n562), .C2(new_n564), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n587), .B1(new_n593), .B2(new_n576), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n577), .B(new_n580), .C1(new_n586), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n232), .B1(new_n462), .B2(new_n238), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n364), .A2(new_n480), .A3(new_n543), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NOR2_X1   g415(.A1(new_n474), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n468), .A2(KEYINPUT92), .A3(new_n463), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n466), .A2(new_n467), .A3(new_n464), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n460), .A2(new_n464), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(KEYINPUT92), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT33), .B1(new_n470), .B2(new_n472), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n602), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT93), .B(G478), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n473), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n413), .A2(KEYINPUT94), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT94), .B1(new_n413), .B2(new_n614), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G472), .B1(new_n345), .B2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n341), .A2(new_n343), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n251), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n598), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n540), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n534), .B2(new_n538), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n423), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n617), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  OAI211_X1 g442(.A(new_n479), .B(new_n400), .C1(new_n410), .C2(new_n412), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n624), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n422), .B(KEYINPUT95), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n621), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n246), .A2(new_n248), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n230), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n250), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n595), .A2(new_n597), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n618), .A2(new_n619), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n480), .A2(new_n640), .A3(new_n543), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G12));
  NAND2_X1  g459(.A1(new_n348), .A2(new_n363), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT20), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n411), .A2(new_n401), .A3(new_n409), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n648), .A2(new_n649), .B1(G475), .B2(new_n399), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n419), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n418), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n650), .A2(new_n479), .A3(new_n623), .A4(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n646), .B(new_n640), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n629), .A2(new_n653), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT97), .B1(new_n658), .B2(new_n623), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT98), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n595), .A2(new_n597), .A3(new_n639), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n348), .B2(new_n363), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n655), .A2(new_n656), .ZN(new_n663));
  INV_X1    g477(.A(new_n629), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(KEYINPUT97), .A3(new_n623), .A4(new_n654), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n662), .A2(new_n663), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  AND2_X1   g483(.A1(new_n539), .A2(new_n542), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT38), .ZN(new_n671));
  INV_X1    g485(.A(new_n639), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n479), .A2(new_n413), .A3(new_n672), .A4(new_n540), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n653), .B(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n595), .A2(new_n597), .A3(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n671), .B(new_n673), .C1(new_n674), .C2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n321), .B1(new_n307), .B2(new_n315), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n238), .B1(new_n335), .B2(new_n352), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n345), .A2(KEYINPUT32), .A3(new_n346), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n348), .A2(KEYINPUT99), .A3(new_n681), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n677), .A2(new_n674), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n678), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT102), .B(G143), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G45));
  NAND3_X1  g509(.A1(new_n413), .A2(new_n614), .A3(new_n654), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n413), .A2(new_n614), .A3(KEYINPUT103), .A4(new_n654), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n640), .A2(new_n646), .A3(new_n623), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  OAI21_X1  g518(.A(new_n625), .B1(new_n615), .B2(new_n616), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n593), .A2(new_n576), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n593), .A2(new_n587), .A3(new_n576), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n596), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n364), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT41), .B(G113), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n364), .A2(new_n630), .A3(new_n631), .A4(new_n711), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT104), .B(G116), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G18));
  NAND3_X1  g532(.A1(new_n709), .A2(new_n597), .A3(new_n623), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n480), .A2(new_n646), .A3(new_n639), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND4_X1  g536(.A1(new_n709), .A2(new_n623), .A3(new_n597), .A4(new_n631), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n326), .A2(new_n328), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n352), .B1(new_n336), .B2(new_n351), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n343), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n618), .A2(new_n726), .A3(new_n251), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n413), .A2(new_n479), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT105), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n425), .ZN(G24));
  NAND3_X1  g547(.A1(new_n618), .A2(new_n639), .A3(new_n726), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n719), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n698), .A2(new_n699), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n203), .ZN(G27));
  NAND2_X1  g551(.A1(new_n569), .A2(new_n574), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n576), .B1(new_n738), .B2(new_n238), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n707), .B2(new_n708), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT106), .B1(new_n740), .B2(new_n596), .ZN(new_n741));
  OAI21_X1  g555(.A(G469), .B1(new_n579), .B2(G902), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n586), .B2(new_n594), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n597), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n670), .A2(new_n622), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n364), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n701), .A2(new_n748), .A3(KEYINPUT42), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n364), .A2(new_n746), .A3(new_n747), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n700), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n364), .A2(new_n746), .A3(new_n658), .A4(new_n747), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  OAI21_X1  g570(.A(G469), .B1(new_n579), .B2(KEYINPUT45), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n569), .A2(new_n574), .A3(KEYINPUT45), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(G469), .A2(G902), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n707), .A2(new_n708), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n761), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n597), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(new_n676), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n641), .A2(new_n672), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT108), .Z(new_n770));
  NAND2_X1  g584(.A1(new_n470), .A2(new_n472), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n603), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n463), .B(new_n444), .C1(new_n454), .C2(new_n459), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT92), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n469), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT33), .B1(new_n775), .B2(new_n604), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n777), .A2(new_n602), .B1(new_n473), .B2(new_n612), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n413), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT107), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n770), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n747), .B(new_n768), .C1(new_n786), .C2(KEYINPUT44), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(KEYINPUT44), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n270), .ZN(G39));
  INV_X1    g604(.A(new_n747), .ZN(new_n791));
  OR4_X1    g605(.A1(new_n646), .A2(new_n700), .A3(new_n251), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n766), .B(new_n597), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(new_n767), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n201), .ZN(G42));
  AOI21_X1  g613(.A(new_n736), .B1(new_n660), .B2(new_n667), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n672), .A2(new_n597), .A3(new_n743), .A4(new_n654), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n686), .B2(new_n687), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n729), .A2(new_n623), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n701), .A2(new_n702), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n736), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT110), .B1(new_n668), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n808), .B(new_n736), .C1(new_n660), .C2(new_n667), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n805), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n716), .B(new_n721), .C1(new_n705), .C2(new_n712), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n732), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n753), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n629), .B1(new_n650), .B2(new_n778), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n621), .A2(new_n543), .A3(new_n817), .A4(new_n631), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n755), .A2(new_n818), .A3(new_n600), .A4(new_n642), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n734), .B1(new_n741), .B2(new_n745), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n698), .A3(new_n699), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n413), .A2(new_n479), .A3(new_n653), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n640), .A3(new_n646), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n791), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n819), .B2(new_n824), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n816), .A2(new_n827), .A3(KEYINPUT53), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n819), .A2(new_n824), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n815), .A3(new_n753), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n668), .A2(new_n804), .A3(new_n806), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n800), .A2(KEYINPUT52), .A3(new_n804), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n813), .A2(new_n829), .B1(new_n836), .B2(KEYINPUT53), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(KEYINPUT112), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n830), .A2(new_n815), .A3(new_n753), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n807), .A2(new_n809), .A3(new_n811), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n805), .ZN(new_n844));
  INV_X1    g658(.A(new_n835), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n845), .B2(new_n805), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n837), .B2(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n840), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n418), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n747), .A2(new_n711), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n784), .A2(new_n853), .A3(new_n364), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n418), .B1(new_n780), .B2(new_n782), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT48), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n364), .A4(new_n854), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n417), .ZN(new_n861));
  INV_X1    g675(.A(new_n688), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n853), .A2(new_n747), .A3(new_n251), .A4(new_n711), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(new_n864), .B2(new_n617), .ZN(new_n865));
  INV_X1    g679(.A(new_n727), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n720), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n860), .B(new_n865), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n711), .A2(new_n622), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n671), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n857), .A2(new_n872), .A3(new_n866), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n857), .A2(new_n866), .A3(new_n874), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n872), .B1(new_n878), .B2(KEYINPUT115), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n877), .A2(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n413), .A2(new_n614), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n862), .A2(new_n863), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT116), .A4(new_n882), .ZN(new_n886));
  INV_X1    g700(.A(new_n734), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n857), .A2(new_n887), .A3(new_n854), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT51), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n857), .A2(new_n866), .A3(new_n747), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n709), .A2(new_n596), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n797), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n871), .B1(new_n881), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n897));
  INV_X1    g711(.A(new_n795), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n796), .B1(new_n766), .B2(new_n597), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n891), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n797), .A2(new_n897), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n896), .B1(new_n903), .B2(new_n890), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n877), .A2(new_n878), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n879), .A2(new_n880), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n895), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n894), .A2(new_n908), .A3(KEYINPUT118), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT118), .B1(new_n894), .B2(new_n908), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n852), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n710), .A2(KEYINPUT49), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n710), .A2(KEYINPUT49), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n251), .A2(new_n540), .A3(new_n597), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n671), .A2(new_n913), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n862), .A3(new_n779), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n912), .A2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n317), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n846), .A2(new_n841), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n815), .A2(new_n753), .A3(KEYINPUT53), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n600), .A2(new_n755), .A3(new_n818), .A4(new_n642), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n821), .A2(new_n823), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n747), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT111), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n922), .A2(new_n926), .A3(new_n826), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n843), .B2(new_n805), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n238), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT56), .B1(new_n929), .B2(G210), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n508), .A2(new_n519), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT119), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT120), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(new_n517), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n920), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n837), .A2(G210), .A3(G902), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n935), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT121), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n919), .B1(new_n940), .B2(new_n935), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n930), .A2(new_n936), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(new_n946), .ZN(G51));
  XOR2_X1   g761(.A(new_n760), .B(KEYINPUT57), .Z(new_n948));
  NOR2_X1   g762(.A1(new_n838), .A2(new_n839), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n591), .A2(new_n592), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n929), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(new_n759), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n919), .B1(new_n953), .B2(new_n955), .ZN(G54));
  INV_X1    g770(.A(new_n411), .ZN(new_n957));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .A4(new_n411), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n920), .ZN(G60));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n777), .B1(new_n852), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n777), .B(new_n964), .C1(new_n949), .C2(new_n950), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n920), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n249), .B1(new_n837), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT123), .B1(new_n972), .B2(new_n919), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n921), .B2(new_n928), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n974), .B(new_n920), .C1(new_n975), .C2(new_n249), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n637), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n972), .A2(new_n919), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n420), .B2(new_n512), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  INV_X1    g799(.A(new_n815), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n818), .A2(new_n600), .A3(new_n642), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n989), .B2(G953), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n932), .B1(G898), .B2(new_n317), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  NOR2_X1   g807(.A1(new_n313), .A2(new_n314), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n406), .B(KEYINPUT126), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(G953), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n810), .A2(new_n693), .A3(new_n703), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n810), .A2(new_n693), .A3(KEYINPUT62), .A4(new_n703), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND4_X1   g816(.A1(new_n364), .A2(new_n677), .A3(new_n817), .A4(new_n747), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n798), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n787), .B2(new_n788), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT127), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  AOI211_X1 g822(.A(new_n1008), .B(new_n1005), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n997), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n810), .A2(new_n703), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n768), .A2(new_n364), .A3(new_n803), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1012), .A2(new_n755), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1013), .B(new_n753), .C1(new_n797), .C2(new_n792), .ZN(new_n1014));
  NOR4_X1   g828(.A1(new_n789), .A2(new_n1011), .A3(new_n1014), .A4(G953), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n651), .A2(new_n317), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n996), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G227), .A2(G900), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(G953), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1010), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(G953), .A3(new_n1018), .A4(new_n996), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1020), .A2(new_n1022), .ZN(G72));
  NOR2_X1   g837(.A1(new_n359), .A2(new_n352), .ZN(new_n1024));
  NOR4_X1   g838(.A1(new_n789), .A2(new_n1011), .A3(new_n1014), .A4(new_n988), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1024), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1024), .A2(new_n679), .A3(new_n1028), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n848), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1029), .A2(new_n920), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1007), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1002), .A2(new_n1006), .A3(KEYINPUT127), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1033), .A2(new_n989), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n1027), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1032), .B1(new_n1036), .B2(new_n679), .ZN(G57));
endmodule


