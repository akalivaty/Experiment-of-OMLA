//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT19), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT72), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT72), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n190), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT71), .B1(new_n194), .B2(G140), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n192), .A3(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT86), .B1(new_n193), .B2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT72), .A2(G125), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(G140), .A3(new_n189), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT86), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(new_n195), .A4(new_n197), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n188), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G125), .B(G140), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT19), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n187), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G237), .ZN(new_n208));
  INV_X1    g022(.A(G953), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G214), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(G237), .A2(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(G143), .A3(G214), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n217), .A3(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n201), .A2(KEYINPUT16), .A3(new_n195), .A4(new_n197), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n200), .A2(new_n189), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT16), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n192), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(G146), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n207), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n205), .A2(new_n187), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n199), .A2(new_n203), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n187), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n215), .A2(KEYINPUT18), .A3(G131), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n212), .B(new_n214), .C1(new_n231), .C2(new_n217), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(KEYINPUT87), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT87), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n207), .A2(new_n225), .B1(new_n229), .B2(new_n233), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(new_n238), .ZN(new_n243));
  MUX2_X1   g057(.A(new_n219), .B(new_n216), .S(KEYINPUT17), .Z(new_n244));
  AOI21_X1  g058(.A(G146), .B1(new_n220), .B2(new_n223), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n246), .A3(new_n224), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n234), .A3(new_n238), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(G475), .A2(G902), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT20), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT88), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n254), .A3(KEYINPUT20), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n249), .A2(new_n256), .A3(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n249), .A2(new_n259), .A3(new_n256), .A4(new_n250), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n255), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n247), .A2(new_n234), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n239), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n248), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G475), .ZN(new_n267));
  XNOR2_X1  g081(.A(G128), .B(G143), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G116), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT14), .A3(G122), .ZN(new_n272));
  XNOR2_X1  g086(.A(G116), .B(G122), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(G107), .B(new_n272), .C1(new_n274), .C2(KEYINPUT14), .ZN(new_n275));
  INV_X1    g089(.A(G107), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n270), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n273), .B(new_n276), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n268), .A2(KEYINPUT13), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  OR3_X1    g095(.A1(new_n281), .A2(KEYINPUT13), .A3(G143), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(G134), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n268), .A2(new_n269), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT9), .B(G234), .ZN(new_n287));
  INV_X1    g101(.A(G217), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n287), .A2(new_n288), .A3(G953), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT90), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n286), .A2(new_n290), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n265), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT15), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G478), .ZN(new_n298));
  INV_X1    g112(.A(G478), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n295), .B(new_n265), .C1(KEYINPUT15), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(G234), .A2(G237), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(G952), .A3(new_n209), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(G902), .A3(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT21), .B(G898), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n261), .A2(new_n267), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G221), .B1(new_n287), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT11), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n269), .B2(G137), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n269), .A2(G137), .ZN(new_n317));
  INV_X1    g131(.A(G137), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT11), .A3(G134), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G131), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n316), .A2(new_n319), .A3(new_n217), .A4(new_n317), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n276), .A2(G104), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n237), .A2(G107), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT79), .B1(new_n327), .B2(G101), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n329));
  INV_X1    g143(.A(G101), .ZN(new_n330));
  AOI211_X1 g144(.A(new_n329), .B(new_n330), .C1(new_n325), .C2(new_n326), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n187), .A2(G143), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n211), .A2(G146), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n336), .A2(G128), .B1(new_n211), .B2(G146), .ZN(new_n337));
  XNOR2_X1  g151(.A(G143), .B(G146), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n335), .A2(new_n337), .B1(G128), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n276), .A3(G104), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n340), .A2(new_n342), .A3(new_n330), .A4(new_n326), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n332), .A2(KEYINPUT10), .A3(new_n339), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n342), .A3(new_n326), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n333), .A2(new_n334), .ZN(new_n348));
  NOR2_X1   g162(.A1(KEYINPUT0), .A2(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT0), .A2(G128), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n338), .A2(new_n350), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n355), .A3(G101), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n347), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n358));
  XNOR2_X1  g172(.A(G104), .B(G107), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n329), .B1(new_n359), .B2(new_n330), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n237), .A2(G107), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n276), .A2(G104), .ZN(new_n362));
  OAI211_X1 g176(.A(KEYINPUT79), .B(G101), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n343), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n211), .A2(G146), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n187), .A2(G143), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n336), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n337), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n367), .A2(new_n368), .B1(new_n281), .B2(new_n348), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n358), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  AND4_X1   g184(.A1(new_n324), .A2(new_n344), .A3(new_n357), .A4(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT78), .B(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n209), .A2(G227), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT77), .B(G110), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n314), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n344), .A2(new_n357), .A3(new_n370), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n323), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n344), .A2(new_n357), .A3(new_n370), .A4(new_n324), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT80), .A3(new_n376), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n364), .A2(new_n369), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n339), .A2(new_n343), .A3(new_n363), .A4(new_n360), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n324), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT12), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT12), .ZN(new_n388));
  AOI211_X1 g202(.A(new_n388), .B(new_n324), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n381), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n377), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n313), .B1(new_n392), .B2(new_n265), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n312), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n376), .B(new_n381), .C1(new_n387), .C2(new_n389), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g213(.A(KEYINPUT82), .B(new_n376), .C1(new_n380), .C2(new_n381), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n313), .B(new_n265), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n383), .B2(new_n391), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n401), .B(KEYINPUT81), .C1(new_n313), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G119), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G116), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT64), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n405), .B2(G116), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n271), .A2(KEYINPUT64), .A3(G119), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT2), .B(G113), .Z(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n406), .ZN(new_n415));
  INV_X1    g229(.A(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n356), .A3(new_n347), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n360), .A2(new_n343), .A3(new_n363), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT5), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n407), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(G113), .B(new_n422), .C1(new_n415), .C2(new_n421), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n423), .A3(new_n413), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G110), .B(G122), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n426), .B(KEYINPUT83), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(new_n433), .A3(new_n428), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n352), .A2(new_n353), .A3(new_n221), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n339), .B2(new_n221), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n209), .A2(G224), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT84), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n428), .A2(KEYINPUT8), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G113), .B1(new_n406), .B2(KEYINPUT5), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT85), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n415), .A2(new_n421), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n420), .B(new_n413), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n413), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n445), .B1(new_n411), .B2(KEYINPUT5), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n364), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n444), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n437), .A2(KEYINPUT7), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n436), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n435), .B(new_n455), .C1(new_n339), .C2(new_n221), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n458), .B2(new_n431), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n440), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n440), .B2(new_n459), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n404), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n213), .A2(G210), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(G101), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n269), .A2(G137), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n318), .A2(G134), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n322), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT65), .B1(new_n369), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n323), .A2(new_n354), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n339), .A2(new_n481), .A3(new_n322), .A4(new_n477), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(KEYINPUT30), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n339), .A2(new_n322), .A3(new_n477), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n418), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n418), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n479), .A2(new_n489), .A3(new_n480), .A4(new_n482), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n474), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n480), .B1(new_n369), .B2(new_n478), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n418), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n418), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n496), .C1(new_n493), .C2(new_n490), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n492), .B1(new_n497), .B2(new_n473), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n483), .A2(new_n418), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n493), .B1(new_n500), .B2(new_n490), .ZN(new_n501));
  INV_X1    g315(.A(new_n495), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n474), .A2(KEYINPUT29), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n265), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G472), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n487), .B1(KEYINPUT30), .B2(new_n483), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n474), .B(new_n490), .C1(new_n507), .C2(new_n489), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT31), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n488), .A2(new_n510), .A3(new_n474), .A4(new_n490), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n497), .A2(new_n473), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT32), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT67), .B(KEYINPUT32), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT68), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n521), .B(new_n518), .C1(new_n513), .C2(new_n514), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n516), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n224), .A2(new_n227), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n405), .B2(G128), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n405), .A2(G128), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n281), .A2(KEYINPUT23), .A3(G119), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT24), .B(G110), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n281), .A2(G119), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n532), .A2(new_n527), .A3(KEYINPUT70), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT70), .B1(new_n532), .B2(new_n527), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n531), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n527), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n532), .A2(new_n527), .A3(KEYINPUT70), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n529), .A2(G110), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT73), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n524), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n542), .A3(new_n538), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n529), .A2(G110), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n246), .B2(new_n224), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT74), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n224), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n547), .B(new_n548), .C1(new_n552), .C2(new_n245), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n543), .A2(KEYINPUT73), .A3(new_n544), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n536), .B1(new_n530), .B2(new_n535), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n553), .B(new_n554), .C1(new_n557), .C2(new_n524), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n209), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT22), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(G137), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n551), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n553), .B(new_n561), .C1(new_n557), .C2(new_n524), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n265), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT76), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G234), .ZN(new_n570));
  OAI21_X1  g384(.A(G217), .B1(new_n570), .B2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT69), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT25), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n565), .B2(new_n566), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n569), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n573), .A2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n563), .A2(new_n564), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n310), .A2(new_n468), .A3(new_n523), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  AND2_X1   g397(.A1(new_n258), .A2(new_n260), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n254), .B1(new_n251), .B2(KEYINPUT20), .ZN(new_n585));
  AOI211_X1 g399(.A(KEYINPUT88), .B(new_n256), .C1(new_n249), .C2(new_n250), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n584), .A2(new_n587), .B1(G475), .B2(new_n266), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n295), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n294), .A2(KEYINPUT33), .A3(new_n291), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(G478), .A3(new_n265), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n296), .A2(new_n299), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT92), .B1(new_n588), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n261), .B2(new_n267), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n308), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n601), .B(new_n464), .C1(new_n461), .C2(new_n462), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n578), .A2(new_n580), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n513), .A2(new_n265), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n395), .A2(new_n606), .A3(new_n403), .A4(new_n517), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  NAND3_X1  g425(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n612), .A2(new_n267), .A3(new_n301), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n513), .B2(new_n265), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n514), .B2(new_n513), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n551), .A2(new_n558), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n579), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(KEYINPUT25), .A3(new_n575), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n572), .B1(new_n577), .B2(new_n568), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n310), .A2(new_n468), .A3(new_n619), .A4(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT37), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT93), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(G110), .Z(G12));
  NOR2_X1   g447(.A1(new_n305), .A2(G900), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT94), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n303), .B(KEYINPUT95), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n267), .A2(new_n612), .A3(new_n301), .A4(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n523), .A3(new_n468), .A4(new_n629), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  XNOR2_X1  g454(.A(new_n637), .B(KEYINPUT39), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n395), .A2(new_n403), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT40), .ZN(new_n643));
  INV_X1    g457(.A(new_n301), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n261), .B2(new_n267), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n463), .B(KEYINPUT38), .Z(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n464), .A4(new_n628), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n500), .A2(new_n490), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n473), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n508), .A2(KEYINPUT96), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n265), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT96), .B1(new_n508), .B2(new_n649), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n515), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n517), .A2(new_n519), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n521), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n517), .A2(KEYINPUT68), .A3(new_n519), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n643), .A2(new_n647), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n628), .B1(new_n661), .B2(new_n516), .ZN(new_n662));
  INV_X1    g476(.A(new_n637), .ZN(new_n663));
  AOI211_X1 g477(.A(new_n663), .B(new_n595), .C1(new_n261), .C2(new_n267), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n664), .A3(new_n468), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  OAI21_X1  g480(.A(new_n265), .B1(new_n399), .B2(new_n400), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n401), .A4(new_n311), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n401), .A3(new_n311), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n523), .A2(new_n581), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n600), .A2(new_n673), .A3(new_n603), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT98), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT41), .B(G113), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND2_X1  g491(.A1(new_n578), .A2(new_n580), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n661), .B2(new_n516), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n672), .A2(new_n670), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n603), .A3(new_n613), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  AND3_X1   g496(.A1(new_n672), .A2(new_n466), .A3(new_n670), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n662), .A2(new_n310), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  OAI21_X1  g499(.A(new_n473), .B1(new_n501), .B2(new_n502), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n509), .A2(new_n511), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(KEYINPUT99), .A3(new_n514), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT99), .B1(new_n687), .B2(new_n514), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n688), .A2(new_n618), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n581), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n672), .A2(new_n601), .A3(new_n670), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n261), .A2(new_n267), .ZN(new_n694));
  AND4_X1   g508(.A1(KEYINPUT100), .A2(new_n694), .A3(new_n301), .A4(new_n466), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT100), .B1(new_n645), .B2(new_n466), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT101), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  NOR2_X1   g513(.A1(new_n628), .A2(new_n663), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n683), .A2(new_n597), .A3(new_n690), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n384), .A2(new_n385), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n388), .B1(new_n704), .B2(new_n324), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n386), .A2(KEYINPUT12), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n371), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n703), .B1(new_n707), .B2(new_n376), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n390), .A2(KEYINPUT102), .A3(new_n377), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(G469), .A3(new_n383), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(G469), .A2(G902), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n401), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n401), .A2(new_n710), .A3(KEYINPUT103), .A4(new_n711), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n311), .A2(new_n464), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n461), .A2(new_n462), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n716), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n597), .A2(new_n637), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT32), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n517), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n516), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n581), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n724), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n716), .A2(new_n721), .A3(new_n718), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n721), .B1(new_n716), .B2(new_n718), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n679), .B(new_n664), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n723), .A2(new_n730), .B1(new_n733), .B2(new_n729), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n217), .ZN(G33));
  NAND3_X1  g549(.A1(new_n723), .A2(new_n679), .A3(new_n638), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n392), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n383), .A4(new_n709), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(G469), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n711), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT46), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n711), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n401), .A3(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(new_n311), .A3(new_n641), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n464), .A3(new_n463), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n694), .A2(new_n595), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n628), .A2(new_n619), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT105), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n747), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NAND2_X1  g571(.A1(new_n745), .A2(new_n311), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT47), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n463), .A2(new_n464), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n523), .A2(new_n581), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n664), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT106), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  NAND3_X1  g578(.A1(new_n694), .A2(new_n594), .A3(new_n690), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n720), .B2(new_n722), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n404), .A2(new_n760), .A3(new_n301), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n612), .A2(new_n267), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n523), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n700), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n261), .A2(new_n267), .A3(new_n301), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n608), .B1(new_n771), .B2(new_n597), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(new_n582), .A3(new_n630), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n736), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n674), .A2(new_n697), .A3(new_n684), .A4(new_n681), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n774), .A2(new_n775), .A3(new_n734), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n716), .A2(new_n628), .A3(new_n311), .A4(new_n637), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n658), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n695), .B2(new_n696), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT107), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n778), .B(new_n781), .C1(new_n695), .C2(new_n696), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n665), .A2(new_n701), .A3(new_n639), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n787), .B(new_n784), .C1(new_n780), .C2(new_n782), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n776), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT109), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n674), .A2(new_n697), .A3(new_n681), .A4(new_n684), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n730), .A2(new_n723), .ZN(new_n796));
  INV_X1    g610(.A(new_n733), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(KEYINPUT42), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT111), .B1(new_n775), .B2(new_n734), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n774), .A2(KEYINPUT110), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n770), .A2(new_n773), .A3(new_n803), .A4(new_n736), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n786), .A2(new_n788), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n789), .A2(new_n809), .A3(new_n790), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n792), .A2(new_n793), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n776), .B(KEYINPUT53), .C1(new_n786), .C2(new_n788), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n791), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT108), .B1(new_n813), .B2(KEYINPUT54), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT108), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n815), .B(new_n793), .C1(new_n791), .C2(new_n812), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n811), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT112), .B(new_n811), .C1(new_n814), .C2(new_n816), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n750), .A2(new_n636), .ZN(new_n821));
  INV_X1    g635(.A(new_n680), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n760), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n629), .A2(new_n690), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n581), .A3(new_n304), .A4(new_n658), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n588), .A2(new_n595), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n824), .A2(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n821), .A2(new_n581), .A3(new_n690), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n822), .A2(new_n464), .A3(new_n646), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n760), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n668), .A2(new_n401), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(new_n312), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n759), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n829), .A2(new_n467), .A3(new_n822), .ZN(new_n840));
  INV_X1    g654(.A(new_n600), .ZN(new_n841));
  OAI211_X1 g655(.A(G952), .B(new_n209), .C1(new_n826), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  INV_X1    g658(.A(new_n728), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n821), .A2(new_n845), .A3(new_n823), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT48), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n843), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n836), .A2(new_n312), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT113), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n835), .B1(new_n759), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT51), .B1(new_n834), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n819), .A2(new_n820), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(G952), .A2(G953), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n646), .A2(new_n678), .A3(new_n717), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n836), .B(KEYINPUT49), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n658), .A3(new_n748), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n858), .A2(KEYINPUT115), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(G75));
  NAND2_X1  g680(.A1(new_n432), .A2(new_n434), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT116), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n439), .B(KEYINPUT55), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n791), .A2(KEYINPUT109), .B1(new_n806), .B2(new_n807), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n265), .B1(new_n873), .B2(new_n810), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(G210), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n209), .A2(G952), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n870), .B1(new_n875), .B2(new_n871), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G51));
  NAND2_X1  g695(.A1(new_n792), .A2(new_n808), .ZN(new_n882));
  INV_X1    g696(.A(new_n810), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT54), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n811), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n711), .B(KEYINPUT57), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n886), .A2(new_n887), .B1(new_n400), .B2(new_n399), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n874), .A2(G469), .A3(new_n739), .A4(new_n740), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n879), .B1(new_n888), .B2(new_n889), .ZN(G54));
  NAND3_X1  g704(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n891));
  INV_X1    g705(.A(new_n249), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n879), .ZN(G60));
  INV_X1    g709(.A(new_n879), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n590), .A2(new_n591), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n299), .A2(new_n265), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n897), .B1(new_n885), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n902), .ZN(new_n904));
  AOI211_X1 g718(.A(KEYINPUT119), .B(new_n904), .C1(new_n884), .C2(new_n811), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n896), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n898), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n819), .A2(new_n820), .ZN(new_n908));
  INV_X1    g722(.A(new_n901), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT120), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n811), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n793), .B1(new_n873), .B2(new_n810), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n902), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT119), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n885), .A2(new_n897), .A3(new_n902), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n879), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n901), .B1(new_n819), .B2(new_n820), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n918), .C1(new_n907), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n911), .A2(new_n920), .ZN(G63));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n896), .B1(new_n922), .B2(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n882), .B2(new_n883), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n563), .A2(new_n564), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT121), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n923), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n622), .B2(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(G66));
  INV_X1    g746(.A(G224), .ZN(new_n933));
  OAI21_X1  g747(.A(G953), .B1(new_n307), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT123), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n794), .A2(new_n773), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n868), .B1(G898), .B2(new_n209), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n938), .B(new_n941), .ZN(G69));
  NAND3_X1  g756(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n204), .A2(new_n206), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n507), .B(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n642), .A2(new_n760), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n679), .B(new_n947), .C1(new_n597), .C2(new_n771), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n756), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n785), .A2(new_n659), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n763), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n943), .B(new_n946), .C1(new_n953), .C2(G953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n746), .B(new_n845), .C1(new_n696), .C2(new_n695), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n955), .A2(new_n798), .A3(new_n736), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n763), .A2(new_n756), .A3(new_n785), .A4(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n209), .ZN(new_n959));
  INV_X1    g773(.A(G227), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(G900), .A3(G953), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n945), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n954), .B1(new_n959), .B2(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n488), .A2(new_n490), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n473), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n813), .B(new_n965), .C1(new_n967), .C2(new_n491), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n896), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n474), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n953), .A2(new_n936), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n965), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n965), .B1(new_n958), .B2(new_n936), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n966), .A2(new_n474), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n969), .B(new_n972), .C1(new_n973), .C2(new_n974), .ZN(G57));
endmodule


