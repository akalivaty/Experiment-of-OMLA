

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U553 ( .A(KEYINPUT74), .B(n576), .Z(n519) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n805) );
  INV_X1 U555 ( .A(G2105), .ZN(n536) );
  NOR2_X1 U556 ( .A1(G651), .A2(n652), .ZN(n664) );
  XNOR2_X1 U557 ( .A(n535), .B(KEYINPUT64), .ZN(n889) );
  XOR2_X1 U558 ( .A(KEYINPUT17), .B(n541), .Z(n893) );
  AND2_X1 U559 ( .A1(n546), .A2(n545), .ZN(G160) );
  XOR2_X1 U560 ( .A(G543), .B(KEYINPUT0), .Z(n652) );
  NAND2_X1 U561 ( .A1(G51), .A2(n664), .ZN(n524) );
  INV_X1 U562 ( .A(G651), .ZN(n520) );
  NOR2_X1 U563 ( .A1(n520), .A2(G543), .ZN(n521) );
  XOR2_X1 U564 ( .A(KEYINPUT68), .B(n521), .Z(n522) );
  XNOR2_X2 U565 ( .A(KEYINPUT1), .B(n522), .ZN(n663) );
  NAND2_X1 U566 ( .A1(G63), .A2(n663), .ZN(n523) );
  NAND2_X1 U567 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U568 ( .A(KEYINPUT6), .B(n525), .ZN(n533) );
  NOR2_X1 U569 ( .A1(n652), .A2(n520), .ZN(n658) );
  NAND2_X1 U570 ( .A1(G76), .A2(n658), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n659) );
  NAND2_X1 U572 ( .A1(G89), .A2(n659), .ZN(n527) );
  XNOR2_X1 U573 ( .A(KEYINPUT80), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U575 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U576 ( .A(n530), .B(KEYINPUT81), .ZN(n531) );
  XNOR2_X1 U577 ( .A(n531), .B(KEYINPUT5), .ZN(n532) );
  NOR2_X1 U578 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U579 ( .A(KEYINPUT7), .B(n534), .Z(G168) );
  XOR2_X1 U580 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U581 ( .A1(n536), .A2(G2104), .ZN(n535) );
  NAND2_X1 U582 ( .A1(G125), .A2(n889), .ZN(n539) );
  AND2_X1 U583 ( .A1(n536), .A2(G2104), .ZN(n892) );
  NAND2_X1 U584 ( .A1(n892), .A2(G101), .ZN(n537) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n537), .Z(n538) );
  NAND2_X1 U586 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n540), .B(KEYINPUT65), .ZN(n546) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n541) );
  NAND2_X1 U589 ( .A1(G137), .A2(n893), .ZN(n544) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U591 ( .A1(G113), .A2(n888), .ZN(n542) );
  XNOR2_X1 U592 ( .A(KEYINPUT66), .B(n542), .ZN(n543) );
  AND2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U594 ( .A1(G102), .A2(n892), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G138), .A2(n893), .ZN(n547) );
  NAND2_X1 U596 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U597 ( .A1(n888), .A2(G114), .ZN(n550) );
  NAND2_X1 U598 ( .A1(G126), .A2(n889), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U600 ( .A1(n552), .A2(n551), .ZN(G164) );
  XNOR2_X1 U601 ( .A(G2451), .B(G2446), .ZN(n562) );
  XOR2_X1 U602 ( .A(G2430), .B(KEYINPUT112), .Z(n554) );
  XNOR2_X1 U603 ( .A(G2454), .B(G2435), .ZN(n553) );
  XNOR2_X1 U604 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U605 ( .A(G2438), .B(KEYINPUT111), .Z(n556) );
  XNOR2_X1 U606 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U607 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U608 ( .A(n558), .B(n557), .Z(n560) );
  XNOR2_X1 U609 ( .A(G2443), .B(G2427), .ZN(n559) );
  XNOR2_X1 U610 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U611 ( .A(n562), .B(n561), .ZN(n563) );
  AND2_X1 U612 ( .A1(n563), .A2(G14), .ZN(G401) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  XOR2_X1 U615 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n565) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U617 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U618 ( .A(KEYINPUT72), .B(n566), .Z(n916) );
  NAND2_X1 U619 ( .A1(n916), .A2(G567), .ZN(n567) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U621 ( .A1(n659), .A2(G81), .ZN(n568) );
  XNOR2_X1 U622 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G68), .A2(n658), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U625 ( .A(n571), .B(KEYINPUT13), .ZN(n573) );
  NAND2_X1 U626 ( .A1(G43), .A2(n664), .ZN(n572) );
  NAND2_X1 U627 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U628 ( .A1(G56), .A2(n663), .ZN(n575) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n574) );
  XNOR2_X1 U630 ( .A(n575), .B(n574), .ZN(n576) );
  NOR2_X1 U631 ( .A1(n577), .A2(n519), .ZN(n578) );
  XOR2_X2 U632 ( .A(KEYINPUT76), .B(n578), .Z(n929) );
  XNOR2_X1 U633 ( .A(G860), .B(KEYINPUT77), .ZN(n608) );
  OR2_X1 U634 ( .A1(n929), .A2(n608), .ZN(G153) );
  NAND2_X1 U635 ( .A1(G77), .A2(n658), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G90), .A2(n659), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U638 ( .A(KEYINPUT9), .B(n581), .ZN(n585) );
  NAND2_X1 U639 ( .A1(n663), .A2(G64), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G52), .A2(n664), .ZN(n582) );
  AND2_X1 U641 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G301), .A2(G868), .ZN(n586) );
  XNOR2_X1 U644 ( .A(n586), .B(KEYINPUT78), .ZN(n596) );
  INV_X1 U645 ( .A(G868), .ZN(n679) );
  NAND2_X1 U646 ( .A1(G66), .A2(n663), .ZN(n593) );
  NAND2_X1 U647 ( .A1(G54), .A2(n664), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G92), .A2(n659), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G79), .A2(n658), .ZN(n589) );
  XNOR2_X1 U651 ( .A(KEYINPUT79), .B(n589), .ZN(n590) );
  NOR2_X1 U652 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U654 ( .A(KEYINPUT15), .B(n594), .ZN(n924) );
  INV_X1 U655 ( .A(n924), .ZN(n706) );
  NAND2_X1 U656 ( .A1(n679), .A2(n706), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n596), .A2(n595), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G91), .A2(n659), .ZN(n597) );
  XNOR2_X1 U659 ( .A(n597), .B(KEYINPUT69), .ZN(n603) );
  NAND2_X1 U660 ( .A1(G65), .A2(n663), .ZN(n598) );
  XNOR2_X1 U661 ( .A(n598), .B(KEYINPUT70), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G53), .A2(n664), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U664 ( .A(KEYINPUT71), .B(n601), .Z(n602) );
  NOR2_X1 U665 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U666 ( .A1(n658), .A2(G78), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n605), .A2(n604), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n679), .ZN(n607) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U670 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n608), .A2(G559), .ZN(n609) );
  NAND2_X1 U672 ( .A1(n609), .A2(n924), .ZN(n610) );
  XNOR2_X1 U673 ( .A(n610), .B(KEYINPUT82), .ZN(n611) );
  XNOR2_X1 U674 ( .A(KEYINPUT16), .B(n611), .ZN(G148) );
  NOR2_X1 U675 ( .A1(n706), .A2(n679), .ZN(n612) );
  XOR2_X1 U676 ( .A(KEYINPUT84), .B(n612), .Z(n613) );
  NOR2_X1 U677 ( .A1(G559), .A2(n613), .ZN(n616) );
  NOR2_X1 U678 ( .A1(n929), .A2(G868), .ZN(n614) );
  XOR2_X1 U679 ( .A(KEYINPUT83), .B(n614), .Z(n615) );
  NOR2_X1 U680 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U681 ( .A1(n889), .A2(G123), .ZN(n617) );
  XNOR2_X1 U682 ( .A(n617), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U683 ( .A1(G99), .A2(n892), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G135), .A2(n893), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U686 ( .A1(G111), .A2(n888), .ZN(n620) );
  XNOR2_X1 U687 ( .A(KEYINPUT85), .B(n620), .ZN(n621) );
  NOR2_X1 U688 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U689 ( .A1(n624), .A2(n623), .ZN(n976) );
  XNOR2_X1 U690 ( .A(G2096), .B(n976), .ZN(n625) );
  NOR2_X1 U691 ( .A1(G2100), .A2(n625), .ZN(n626) );
  XOR2_X1 U692 ( .A(KEYINPUT86), .B(n626), .Z(G156) );
  XOR2_X1 U693 ( .A(n929), .B(KEYINPUT87), .Z(n628) );
  NAND2_X1 U694 ( .A1(G559), .A2(n924), .ZN(n627) );
  XNOR2_X1 U695 ( .A(n628), .B(n627), .ZN(n676) );
  NOR2_X1 U696 ( .A1(G860), .A2(n676), .ZN(n635) );
  NAND2_X1 U697 ( .A1(G55), .A2(n664), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G67), .A2(n663), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U700 ( .A1(G80), .A2(n658), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G93), .A2(n659), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n678) );
  XNOR2_X1 U704 ( .A(n635), .B(n678), .ZN(G145) );
  NAND2_X1 U705 ( .A1(G48), .A2(n664), .ZN(n637) );
  NAND2_X1 U706 ( .A1(G86), .A2(n659), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U708 ( .A1(G73), .A2(n658), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(KEYINPUT2), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n639), .B(KEYINPUT89), .ZN(n640) );
  NOR2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U712 ( .A1(G61), .A2(n663), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G50), .A2(n664), .ZN(n645) );
  NAND2_X1 U715 ( .A1(G88), .A2(n659), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n658), .A2(G75), .ZN(n646) );
  XOR2_X1 U718 ( .A(KEYINPUT90), .B(n646), .Z(n647) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U720 ( .A1(G62), .A2(n663), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(G303) );
  NAND2_X1 U722 ( .A1(G49), .A2(n664), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n651), .B(KEYINPUT88), .ZN(n657) );
  NAND2_X1 U724 ( .A1(G87), .A2(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n663), .A2(n655), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n657), .A2(n656), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G72), .A2(n658), .ZN(n661) );
  NAND2_X1 U730 ( .A1(G85), .A2(n659), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(KEYINPUT67), .B(n662), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n663), .A2(G60), .ZN(n666) );
  NAND2_X1 U734 ( .A1(G47), .A2(n664), .ZN(n665) );
  AND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U736 ( .A1(n668), .A2(n667), .ZN(G290) );
  XNOR2_X1 U737 ( .A(n678), .B(G305), .ZN(n674) );
  XNOR2_X1 U738 ( .A(KEYINPUT92), .B(KEYINPUT19), .ZN(n670) );
  XNOR2_X1 U739 ( .A(G288), .B(KEYINPUT91), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U741 ( .A(G303), .B(n671), .Z(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(G290), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n675) );
  XOR2_X1 U744 ( .A(G299), .B(n675), .Z(n905) );
  XNOR2_X1 U745 ( .A(n905), .B(n676), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n677), .A2(G868), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(KEYINPUT93), .B(n682), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n683) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n683), .Z(n684) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(KEYINPUT95), .Z(n688) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U759 ( .A(n689), .B(KEYINPUT94), .ZN(n690) );
  NOR2_X1 U760 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U761 ( .A1(G96), .A2(n691), .ZN(n839) );
  NAND2_X1 U762 ( .A1(n839), .A2(G2106), .ZN(n695) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n692) );
  NOR2_X1 U764 ( .A1(G237), .A2(n692), .ZN(n693) );
  NAND2_X1 U765 ( .A1(G108), .A2(n693), .ZN(n840) );
  NAND2_X1 U766 ( .A1(n840), .A2(G567), .ZN(n694) );
  NAND2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n915) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n696) );
  NOR2_X1 U769 ( .A1(n915), .A2(n696), .ZN(n838) );
  NAND2_X1 U770 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U771 ( .A(G301), .ZN(G171) );
  INV_X1 U772 ( .A(G299), .ZN(n921) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n804) );
  INV_X1 U774 ( .A(n805), .ZN(n697) );
  NOR2_X4 U775 ( .A1(n804), .A2(n697), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n724), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U777 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U778 ( .A(G1956), .ZN(n922) );
  NOR2_X1 U779 ( .A1(n922), .A2(n724), .ZN(n699) );
  NOR2_X1 U780 ( .A1(n700), .A2(n699), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n921), .A2(n710), .ZN(n701) );
  XOR2_X1 U782 ( .A(n701), .B(KEYINPUT28), .Z(n721) );
  AND2_X1 U783 ( .A1(n724), .A2(G1996), .ZN(n702) );
  XNOR2_X1 U784 ( .A(KEYINPUT26), .B(n702), .ZN(n703) );
  NOR2_X1 U785 ( .A1(n929), .A2(n703), .ZN(n705) );
  INV_X1 U786 ( .A(n724), .ZN(n740) );
  NAND2_X1 U787 ( .A1(G1341), .A2(n740), .ZN(n704) );
  NAND2_X1 U788 ( .A1(n705), .A2(n704), .ZN(n717) );
  NOR2_X1 U789 ( .A1(n717), .A2(n706), .ZN(n707) );
  XNOR2_X1 U790 ( .A(n707), .B(KEYINPUT103), .ZN(n713) );
  NOR2_X1 U791 ( .A1(G2067), .A2(n740), .ZN(n709) );
  NOR2_X1 U792 ( .A1(n724), .A2(G1348), .ZN(n708) );
  NOR2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U794 ( .A1(n921), .A2(n710), .ZN(n714) );
  AND2_X1 U795 ( .A1(n711), .A2(n714), .ZN(n712) );
  NAND2_X1 U796 ( .A1(n713), .A2(n712), .ZN(n719) );
  INV_X1 U797 ( .A(n714), .ZN(n715) );
  NOR2_X1 U798 ( .A1(n924), .A2(n715), .ZN(n716) );
  NAND2_X1 U799 ( .A1(n717), .A2(n716), .ZN(n718) );
  AND2_X1 U800 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U801 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U802 ( .A(KEYINPUT29), .B(n722), .Z(n728) );
  NOR2_X1 U803 ( .A1(n724), .A2(G1961), .ZN(n723) );
  XOR2_X1 U804 ( .A(KEYINPUT102), .B(n723), .Z(n726) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n1002) );
  NAND2_X1 U806 ( .A1(n724), .A2(n1002), .ZN(n725) );
  NAND2_X1 U807 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U808 ( .A1(n732), .A2(G171), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n728), .A2(n727), .ZN(n738) );
  NAND2_X1 U810 ( .A1(G8), .A2(n740), .ZN(n781) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n781), .ZN(n752) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n740), .ZN(n749) );
  NOR2_X1 U813 ( .A1(n752), .A2(n749), .ZN(n729) );
  NAND2_X1 U814 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U816 ( .A1(G168), .A2(n731), .ZN(n734) );
  NOR2_X1 U817 ( .A1(G171), .A2(n732), .ZN(n733) );
  NOR2_X1 U818 ( .A1(n734), .A2(n733), .ZN(n736) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(KEYINPUT104), .Z(n735) );
  XNOR2_X1 U820 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n738), .A2(n737), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n750), .A2(G286), .ZN(n745) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n781), .ZN(n739) );
  XOR2_X1 U824 ( .A(KEYINPUT105), .B(n739), .Z(n742) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U828 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U829 ( .A(n746), .B(KEYINPUT106), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n747), .A2(G8), .ZN(n748) );
  XNOR2_X1 U831 ( .A(n748), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U832 ( .A1(G8), .A2(n749), .ZN(n754) );
  INV_X1 U833 ( .A(n750), .ZN(n751) );
  NOR2_X1 U834 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U835 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U836 ( .A1(n756), .A2(n755), .ZN(n774) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n937) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n757) );
  XOR2_X1 U839 ( .A(n757), .B(KEYINPUT107), .Z(n758) );
  NOR2_X1 U840 ( .A1(n937), .A2(n758), .ZN(n760) );
  INV_X1 U841 ( .A(KEYINPUT33), .ZN(n759) );
  AND2_X1 U842 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U843 ( .A1(n774), .A2(n761), .ZN(n770) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n918) );
  NAND2_X1 U845 ( .A1(G288), .A2(G1976), .ZN(n762) );
  XNOR2_X1 U846 ( .A(n762), .B(KEYINPUT108), .ZN(n934) );
  INV_X1 U847 ( .A(n934), .ZN(n763) );
  NOR2_X1 U848 ( .A1(n763), .A2(n781), .ZN(n764) );
  NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n764), .ZN(n767) );
  NAND2_X1 U850 ( .A1(n937), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U851 ( .A1(n765), .A2(n781), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U853 ( .A1(n918), .A2(n768), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U855 ( .A(KEYINPUT109), .B(n771), .Z(n777) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n781), .A2(n775), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n777), .A2(n776), .ZN(n825) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XNOR2_X1 U862 ( .A(n778), .B(KEYINPUT24), .ZN(n779) );
  XNOR2_X1 U863 ( .A(n779), .B(KEYINPUT101), .ZN(n780) );
  NOR2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n823) );
  INV_X1 U865 ( .A(G1996), .ZN(n998) );
  NAND2_X1 U866 ( .A1(G141), .A2(n893), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT100), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G105), .A2(n892), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT38), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n888), .A2(G117), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G129), .A2(n889), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n880) );
  AND2_X1 U875 ( .A1(n998), .A2(n880), .ZN(n987) );
  XOR2_X1 U876 ( .A(KEYINPUT99), .B(G1991), .Z(n1008) );
  NAND2_X1 U877 ( .A1(G95), .A2(n892), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G107), .A2(n888), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G119), .A2(n889), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(KEYINPUT98), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G131), .A2(n893), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n881) );
  NOR2_X1 U885 ( .A1(n1008), .A2(n881), .ZN(n975) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n797) );
  XNOR2_X1 U887 ( .A(KEYINPUT110), .B(n797), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n975), .A2(n798), .ZN(n801) );
  AND2_X1 U889 ( .A1(n881), .A2(n1008), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n880), .A2(n998), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n826) );
  INV_X1 U892 ( .A(n826), .ZN(n979) );
  NOR2_X1 U893 ( .A1(n801), .A2(n979), .ZN(n802) );
  NOR2_X1 U894 ( .A1(n987), .A2(n802), .ZN(n803) );
  XNOR2_X1 U895 ( .A(n803), .B(KEYINPUT39), .ZN(n818) );
  NOR2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n827) );
  XNOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NAND2_X1 U898 ( .A1(n892), .A2(G104), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(KEYINPUT96), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G140), .A2(n893), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n809), .ZN(n814) );
  NAND2_X1 U903 ( .A1(n888), .A2(G116), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G128), .A2(n889), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n815), .ZN(n885) );
  NOR2_X1 U909 ( .A1(n819), .A2(n885), .ZN(n973) );
  NAND2_X1 U910 ( .A1(n827), .A2(n973), .ZN(n816) );
  XNOR2_X1 U911 ( .A(KEYINPUT97), .B(n816), .ZN(n829) );
  INV_X1 U912 ( .A(n829), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n819), .A2(n885), .ZN(n971) );
  NAND2_X1 U915 ( .A1(n820), .A2(n971), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n821), .A2(n827), .ZN(n832) );
  INV_X1 U917 ( .A(n832), .ZN(n822) );
  OR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n834) );
  XOR2_X1 U920 ( .A(G1986), .B(G290), .Z(n928) );
  NAND2_X1 U921 ( .A1(n928), .A2(n826), .ZN(n828) );
  AND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n830) );
  OR2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  AND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n835), .ZN(G329) );
  INV_X1 U927 ( .A(G303), .ZN(G166) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n916), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U930 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U934 ( .A(G132), .ZN(G219) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G82), .ZN(G220) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XOR2_X1 U941 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U942 ( .A(KEYINPUT113), .B(G2678), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2096), .B(G2100), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U950 ( .A(G2084), .B(G2078), .Z(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U952 ( .A(G1991), .B(G1986), .Z(n852) );
  XOR2_X1 U953 ( .A(G1961), .B(n922), .Z(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U955 ( .A(G1976), .B(G1981), .Z(n854) );
  XNOR2_X1 U956 ( .A(G1966), .B(G1971), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U958 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2474), .B(KEYINPUT41), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(KEYINPUT115), .B(n859), .ZN(n860) );
  XOR2_X1 U962 ( .A(n860), .B(G1996), .Z(G229) );
  NAND2_X1 U963 ( .A1(n889), .A2(G124), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n861), .B(KEYINPUT44), .ZN(n862) );
  XNOR2_X1 U965 ( .A(KEYINPUT116), .B(n862), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G100), .A2(n892), .ZN(n863) );
  XOR2_X1 U967 ( .A(KEYINPUT117), .B(n863), .Z(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G112), .A2(n888), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G136), .A2(n893), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n879) );
  NAND2_X1 U974 ( .A1(G103), .A2(n892), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G139), .A2(n893), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n888), .A2(G115), .ZN(n873) );
  NAND2_X1 U978 ( .A1(G127), .A2(n889), .ZN(n872) );
  NAND2_X1 U979 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  XNOR2_X1 U981 ( .A(KEYINPUT118), .B(n875), .ZN(n876) );
  NOR2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n982) );
  XNOR2_X1 U983 ( .A(G164), .B(n982), .ZN(n878) );
  XNOR2_X1 U984 ( .A(n879), .B(n878), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n882), .B(n976), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n885), .B(G162), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n901) );
  NAND2_X1 U990 ( .A1(n888), .A2(G118), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G106), .A2(n892), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G142), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT45), .B(n896), .Z(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(G160), .B(n899), .Z(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U1001 ( .A(G286), .B(n929), .Z(n904) );
  XOR2_X1 U1002 ( .A(G301), .B(n924), .Z(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n915), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT119), .B(n908), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT120), .B(n912), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n915), .ZN(G319) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n916), .ZN(G223) );
  XNOR2_X1 U1018 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n917) );
  XOR2_X1 U1019 ( .A(G16), .B(n917), .Z(n944) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G168), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(n920), .B(KEYINPUT57), .ZN(n942) );
  XOR2_X1 U1023 ( .A(n922), .B(n921), .Z(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(KEYINPUT124), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G171), .B(G1961), .Z(n926) );
  XOR2_X1 U1026 ( .A(n924), .B(G1348), .Z(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G1341), .B(n929), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G303), .B(G1971), .Z(n935) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT125), .B(n938), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n969) );
  INV_X1 U1039 ( .A(G16), .ZN(n967) );
  XOR2_X1 U1040 ( .A(G20), .B(G1956), .Z(n948) );
  XNOR2_X1 U1041 ( .A(G1341), .B(G19), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G6), .B(G1981), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT59), .B(G1348), .Z(n949) );
  XNOR2_X1 U1046 ( .A(G4), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n952), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G1961), .B(G5), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT126), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n965), .B(KEYINPUT61), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n970), .B(KEYINPUT127), .ZN(n997) );
  INV_X1 U1065 ( .A(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n981) );
  XOR2_X1 U1067 ( .A(G2084), .B(G160), .Z(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n992) );
  XOR2_X1 U1072 ( .A(G2072), .B(n982), .Z(n984) );
  XOR2_X1 U1073 ( .A(G164), .B(G2078), .Z(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(KEYINPUT50), .B(n985), .ZN(n990) );
  XOR2_X1 U1076 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1078 ( .A(KEYINPUT51), .B(n988), .Z(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n993), .ZN(n994) );
  INV_X1 U1082 ( .A(KEYINPUT55), .ZN(n1017) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n1017), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n995), .A2(G29), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1024) );
  XOR2_X1 U1086 ( .A(n998), .B(G32), .Z(n1000) );
  XNOR2_X1 U1087 ( .A(G26), .B(G2067), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1007) );
  XOR2_X1 U1089 ( .A(G2072), .B(G33), .Z(n1001) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(G28), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G27), .B(n1002), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(KEYINPUT121), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G25), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(KEYINPUT53), .B(n1011), .Z(n1014) );
  XOR2_X1 U1098 ( .A(KEYINPUT54), .B(G34), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(G2084), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G35), .B(G2090), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(n1018), .B(n1017), .Z(n1020) );
  INV_X1 U1104 ( .A(G29), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(G11), .A2(n1021), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(KEYINPUT122), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .Z(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
endmodule

