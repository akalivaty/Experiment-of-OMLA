//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0002(.A(G50), .B1(G58), .B2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G13), .ZN(new_n205));
  OR3_X1    g0005(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n206), .B(new_n210), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(KEYINPUT1), .B2(new_n217), .ZN(G361));
  XNOR2_X1  g0019(.A(G238), .B(G244), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT2), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(G250), .B(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G264), .B(G270), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n224), .B(new_n227), .ZN(G358));
  XOR2_X1   g0028(.A(G68), .B(G77), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G50), .B(G58), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G351));
  INV_X1    g0037(.A(G33), .ZN(new_n238));
  INV_X1    g0038(.A(G41), .ZN(new_n239));
  OAI211_X1 g0039(.A(G1), .B(G13), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G274), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G45), .ZN(new_n244));
  AOI21_X1  g0044(.A(G1), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G226), .ZN(new_n247));
  OR2_X1    g0047(.A1(new_n241), .A2(new_n245), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n252));
  AND3_X1   g0052(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT67), .ZN(new_n253));
  AOI21_X1  g0053(.A(KEYINPUT67), .B1(new_n251), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G222), .B1(new_n255), .B2(G77), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n250), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G1698), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n257), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n249), .B1(new_n267), .B2(new_n241), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G190), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n205), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n238), .A2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n272), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G50), .A2(G58), .ZN(new_n279));
  INV_X1    g0079(.A(G68), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n204), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n271), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n270), .A2(new_n205), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G1), .B2(new_n204), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n282), .B(new_n287), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G200), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n269), .B(new_n294), .C1(new_n295), .C2(new_n268), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n268), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n268), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n290), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT12), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n284), .B2(G68), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n285), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n306), .B(new_n307), .C1(new_n289), .C2(new_n280), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n280), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n274), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n314), .A2(new_n271), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n317));
  AND4_X1   g0117(.A1(new_n310), .A2(new_n311), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT73), .A2(G169), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  OAI211_X1 g0123(.A(G226), .B(new_n323), .C1(new_n253), .C2(new_n254), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT70), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n263), .A2(new_n326), .A3(G226), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n223), .B1(new_n261), .B2(new_n262), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n241), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n246), .B1(new_n333), .B2(new_n248), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n322), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n240), .B1(new_n328), .B2(new_n330), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n337), .A2(KEYINPUT13), .A3(new_n334), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n320), .B(new_n321), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(new_n322), .A3(new_n335), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT13), .B1(new_n337), .B2(new_n334), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(G179), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n341), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n320), .B1(new_n344), .B2(new_n321), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n319), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(new_n341), .A3(G190), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT71), .B1(new_n344), .B2(G200), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  AOI211_X1 g0149(.A(new_n349), .B(new_n295), .C1(new_n340), .C2(new_n341), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n318), .B(new_n347), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT68), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n264), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G238), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n329), .A2(new_n323), .B1(new_n255), .B2(G107), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n240), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n246), .ZN(new_n359));
  INV_X1    g0159(.A(new_n248), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(G244), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n353), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT15), .B(G87), .Z(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n273), .B1(G20), .B2(G77), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n272), .B2(new_n277), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n271), .ZN(new_n367));
  INV_X1    g0167(.A(new_n289), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G77), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n369), .C1(G77), .C2(new_n284), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n357), .B1(new_n265), .B2(new_n333), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n241), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n361), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n363), .B(new_n370), .C1(G179), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n370), .B1(new_n373), .B2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n373), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n304), .A2(new_n352), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(G58), .B(G68), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n204), .A2(KEYINPUT7), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT74), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT74), .A2(G33), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n250), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n252), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n261), .A2(new_n204), .A3(new_n262), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n380), .B1(new_n388), .B2(new_n280), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT75), .B1(new_n389), .B2(new_n390), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n238), .ZN(new_n394));
  NAND2_X1  g0194(.A1(KEYINPUT74), .A2(G33), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(KEYINPUT3), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(G20), .B1(new_n396), .B2(new_n251), .ZN(new_n397));
  OAI21_X1  g0197(.A(G68), .B1(new_n397), .B2(new_n387), .ZN(new_n398));
  AOI211_X1 g0198(.A(KEYINPUT7), .B(G20), .C1(new_n396), .C2(new_n251), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT16), .B(new_n380), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n271), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n391), .A2(new_n392), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n272), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n284), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n368), .B2(new_n403), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT76), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT75), .ZN(new_n408));
  INV_X1    g0208(.A(new_n380), .ZN(new_n409));
  INV_X1    g0209(.A(new_n385), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n253), .A2(new_n254), .A3(G20), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(KEYINPUT7), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(G68), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n413), .B2(KEYINPUT16), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n415));
  INV_X1    g0215(.A(new_n401), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n405), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n246), .B1(new_n223), .B2(new_n248), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n382), .A2(new_n383), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n259), .B1(new_n421), .B2(KEYINPUT3), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G223), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n247), .B2(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n240), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G179), .ZN(new_n429));
  OAI21_X1  g0229(.A(G169), .B1(new_n420), .B2(new_n427), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n407), .A2(new_n419), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT18), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n428), .A2(new_n295), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n420), .A2(new_n427), .A3(new_n376), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n417), .A2(new_n405), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n389), .A2(new_n390), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n401), .B1(new_n408), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n406), .B1(new_n440), .B2(new_n415), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n436), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n407), .A2(new_n445), .A3(new_n419), .A4(new_n431), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n433), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n378), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n388), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n388), .B2(new_n449), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n454));
  INV_X1    g0254(.A(G97), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G97), .A2(G107), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n458), .B2(KEYINPUT6), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n451), .A2(new_n453), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n271), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  INV_X1    g0263(.A(G244), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n263), .A2(new_n323), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n396), .A2(new_n251), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n463), .B1(new_n468), .B2(new_n464), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G250), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n255), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(G1698), .B1(new_n472), .B2(new_n463), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n240), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n283), .B(G45), .C1(new_n239), .C2(KEYINPUT5), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n243), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n475), .A2(new_n476), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G257), .A3(new_n240), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(G200), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n285), .A2(new_n455), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n288), .B(new_n284), .C1(G1), .C2(new_n238), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n455), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n263), .A2(G250), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n323), .B1(new_n488), .B2(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n241), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n481), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(G190), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n462), .A2(new_n482), .A3(new_n486), .A4(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n353), .B1(new_n474), .B2(new_n481), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n300), .A3(new_n491), .ZN(new_n495));
  INV_X1    g0295(.A(new_n460), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n450), .B2(KEYINPUT77), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n288), .B1(new_n497), .B2(new_n453), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n494), .B(new_n495), .C1(new_n498), .C2(new_n485), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n364), .A2(new_n284), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n422), .A2(new_n204), .A3(G68), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT19), .B1(new_n273), .B2(G97), .ZN(new_n502));
  INV_X1    g0302(.A(G87), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n455), .A3(new_n449), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G97), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(new_n204), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n502), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n500), .B1(new_n509), .B2(new_n271), .ZN(new_n510));
  INV_X1    g0310(.A(new_n364), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n484), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n283), .A2(new_n242), .A3(G45), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n471), .B1(new_n244), .B2(G1), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n240), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(G116), .B1(new_n382), .B2(new_n383), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n464), .A2(G1698), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G238), .B2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(new_n468), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n520), .B2(new_n241), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n300), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n521), .A2(G169), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n512), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n484), .A2(new_n503), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n500), .B(new_n525), .C1(new_n509), .C2(new_n271), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(G190), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n295), .C2(new_n521), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n493), .A2(new_n499), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT79), .B1(new_n484), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n285), .B1(new_n283), .B2(G33), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(G116), .A4(new_n288), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n532), .A2(new_n535), .B1(new_n531), .B2(new_n285), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT80), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(G20), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n271), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n271), .B2(new_n538), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n467), .B(new_n204), .C1(G33), .C2(new_n455), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT20), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(KEYINPUT20), .B(new_n542), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n536), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n255), .A2(G303), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n323), .A2(G264), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G257), .A2(G1698), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n422), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n240), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n479), .A2(G270), .A3(new_n240), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n478), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT78), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G303), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n263), .A2(new_n556), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n468), .A2(new_n548), .A3(new_n549), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n241), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT78), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n478), .A2(new_n553), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n546), .A2(new_n555), .A3(G169), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n552), .A2(new_n300), .A3(new_n554), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n563), .A2(new_n564), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n546), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n555), .A2(new_n562), .A3(G200), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n552), .A2(KEYINPUT78), .A3(new_n554), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n567), .B(new_n568), .C1(new_n571), .C2(new_n376), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n571), .A2(KEYINPUT21), .A3(G169), .A4(new_n546), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n471), .A2(new_n323), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G257), .B2(new_n323), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n468), .A2(new_n576), .B1(new_n577), .B2(new_n421), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n241), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT86), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n479), .A2(new_n580), .A3(G264), .A4(new_n240), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n240), .B(G264), .C1(new_n475), .C2(new_n476), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT86), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(new_n584), .A3(new_n478), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n241), .A2(new_n578), .B1(new_n581), .B2(new_n583), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G179), .A3(new_n478), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n449), .A2(G20), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n593), .A2(KEYINPUT23), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n204), .B(G116), .C1(new_n382), .C2(new_n383), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(KEYINPUT23), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n594), .A2(new_n595), .A3(new_n599), .A4(new_n596), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT83), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n598), .A2(new_n600), .B1(new_n601), .B2(KEYINPUT24), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n503), .A2(KEYINPUT22), .A3(G20), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n253), .B2(new_n254), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n263), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n396), .A2(new_n204), .A3(G87), .A4(new_n251), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT22), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n602), .B(new_n610), .C1(new_n601), .C2(KEYINPUT24), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n271), .A3(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT84), .B(KEYINPUT25), .C1(new_n284), .C2(G107), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT25), .ZN(new_n618));
  AOI21_X1  g0418(.A(G107), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n285), .B(new_n619), .C1(new_n617), .C2(new_n618), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n616), .B(new_n620), .C1(new_n484), .C2(new_n449), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT85), .Z(new_n622));
  AOI22_X1  g0422(.A1(new_n591), .A2(new_n592), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n585), .A2(new_n376), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n295), .B1(new_n587), .B2(new_n478), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n615), .A2(new_n626), .A3(new_n622), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n448), .A2(new_n530), .A3(new_n574), .A4(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n524), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n529), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n499), .ZN(new_n633));
  INV_X1    g0433(.A(new_n499), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n529), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n630), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n627), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n566), .A2(new_n573), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n615), .A2(new_n622), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n589), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n530), .B(new_n637), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n448), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n431), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT18), .B1(new_n441), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n445), .B(new_n431), .C1(new_n402), .C2(new_n406), .ZN(new_n646));
  INV_X1    g0446(.A(new_n346), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n374), .A2(KEYINPUT88), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n358), .A2(new_n362), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n300), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT88), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n363), .A4(new_n370), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n647), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n351), .A2(new_n444), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n645), .B(new_n646), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n298), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n303), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n643), .A2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n283), .A2(new_n204), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n567), .A2(new_n665), .ZN(new_n666));
  MUX2_X1   g0466(.A(new_n574), .B(new_n638), .S(new_n666), .Z(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n639), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n628), .B1(new_n669), .B2(new_n665), .ZN(new_n670));
  INV_X1    g0470(.A(new_n623), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n638), .A2(new_n665), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n628), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n640), .A2(new_n665), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(KEYINPUT89), .A3(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n673), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n208), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n504), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n203), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n521), .A2(new_n579), .A3(new_n584), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n565), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n474), .A2(new_n481), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT92), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n587), .A2(new_n696), .A3(new_n521), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n694), .A2(KEYINPUT30), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n490), .A2(new_n491), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n521), .A2(G179), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n571), .A2(new_n699), .A3(new_n585), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n693), .A2(new_n565), .A3(new_n697), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n699), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n664), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT91), .B(KEYINPUT31), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n706), .A2(KEYINPUT93), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT93), .B1(new_n706), .B2(new_n707), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n530), .A2(new_n574), .A3(new_n628), .A4(new_n665), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n708), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n664), .B1(new_n636), .B2(new_n641), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n671), .A2(new_n573), .A3(new_n566), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n493), .A2(new_n499), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n528), .A4(new_n637), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n664), .B1(new_n720), .B2(new_n636), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n715), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  INV_X1    g0524(.A(G13), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G45), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n686), .A2(G1), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n668), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G330), .B2(new_n667), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n205), .B1(G20), .B2(new_n353), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n255), .A2(new_n684), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT94), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n739), .A2(G355), .B1(new_n531), .B2(new_n684), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n422), .A2(new_n684), .ZN(new_n741));
  INV_X1    g0541(.A(new_n203), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n244), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n741), .B(new_n743), .C1(new_n232), .C2(new_n244), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n737), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n204), .A2(new_n300), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(new_n376), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n376), .A2(new_n295), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n204), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n748), .A2(G322), .B1(G303), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n747), .A2(new_n295), .A3(G190), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT33), .B(G317), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n754), .A2(new_n755), .B1(new_n758), .B2(G311), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n750), .A2(new_n756), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G329), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n753), .B(new_n759), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n746), .A2(new_n749), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n750), .A2(new_n376), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G326), .A2(new_n768), .B1(new_n770), .B2(G283), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n376), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n204), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n771), .B(new_n255), .C1(new_n577), .C2(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n748), .A2(G58), .B1(G107), .B2(new_n770), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n754), .A2(G68), .B1(new_n768), .B2(G50), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G77), .A2(new_n758), .B1(new_n752), .B2(G87), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n775), .A2(new_n776), .A3(new_n263), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  OR3_X1    g0579(.A1(new_n760), .A2(KEYINPUT32), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT32), .B1(new_n760), .B2(new_n779), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n780), .B(new_n781), .C1(new_n455), .C2(new_n773), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n766), .A2(new_n774), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n728), .B(new_n745), .C1(new_n735), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n734), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n667), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n731), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n370), .A2(new_n664), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n648), .A2(new_n652), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n377), .A2(new_n374), .A3(new_n789), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n716), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n793), .B(KEYINPUT98), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n716), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n729), .B1(new_n796), .B2(new_n714), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n714), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n735), .A2(new_n732), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n729), .B1(G77), .B2(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n767), .A2(new_n556), .B1(new_n751), .B2(new_n449), .ZN(new_n802));
  INV_X1    g0602(.A(new_n754), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n255), .B1(new_n503), .B2(new_n769), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(G116), .C2(new_n758), .ZN(new_n806));
  INV_X1    g0606(.A(new_n773), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G294), .A2(new_n748), .B1(new_n807), .B2(G97), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT96), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n806), .B(new_n809), .C1(new_n810), .C2(new_n764), .ZN(new_n811));
  INV_X1    g0611(.A(new_n764), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n468), .B1(new_n812), .B2(G132), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT97), .Z(new_n814));
  AOI22_X1  g0614(.A1(new_n754), .A2(G150), .B1(new_n768), .B2(G137), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  INV_X1    g0616(.A(new_n748), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n779), .C2(new_n757), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n751), .A2(new_n286), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n769), .A2(new_n280), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(G58), .C2(new_n807), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n811), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n801), .B1(new_n826), .B2(new_n735), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n793), .B2(new_n733), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n798), .A2(new_n828), .ZN(G384));
  NOR2_X1   g0629(.A1(new_n726), .A2(new_n283), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n380), .B1(new_n398), .B2(new_n399), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(new_n390), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n405), .B1(new_n832), .B2(new_n401), .ZN(new_n833));
  INV_X1    g0633(.A(new_n662), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n447), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n407), .A2(new_n419), .A3(new_n834), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n437), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n432), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n833), .B1(new_n431), .B2(new_n834), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n437), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n837), .A2(KEYINPUT38), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n838), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n442), .B1(new_n441), .B2(new_n436), .ZN(new_n849));
  AND4_X1   g0649(.A1(new_n442), .A2(new_n417), .A3(new_n405), .A4(new_n436), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n645), .A2(new_n646), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n432), .A2(new_n838), .A3(new_n841), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n417), .A2(new_n405), .A3(new_n436), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n644), .B1(new_n417), .B2(new_n405), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n839), .B1(new_n857), .B2(new_n838), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n853), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n847), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n432), .A2(KEYINPUT18), .B1(new_n438), .B2(new_n443), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n835), .B1(new_n864), .B2(new_n446), .ZN(new_n865));
  AOI211_X1 g0665(.A(KEYINPUT76), .B(new_n406), .C1(new_n440), .C2(new_n415), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n418), .B1(new_n417), .B2(new_n405), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n840), .B1(new_n868), .B2(new_n431), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n844), .B1(new_n869), .B2(new_n838), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n860), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n862), .B1(new_n871), .B2(new_n847), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT100), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n865), .A2(new_n870), .A3(new_n860), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n837), .B2(new_n846), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT39), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n847), .A2(new_n861), .A3(new_n862), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n647), .A2(new_n665), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n873), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n374), .A2(new_n664), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n794), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n318), .A2(new_n665), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n346), .A2(new_n351), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n343), .B2(new_n345), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n871), .A2(new_n847), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n893), .A2(new_n894), .B1(new_n852), .B2(new_n662), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n882), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n448), .A2(new_n717), .A3(new_n722), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n657), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n706), .A2(new_n707), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n712), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n448), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n891), .A2(new_n793), .A3(new_n902), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT40), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n891), .A2(new_n793), .A3(new_n902), .A4(KEYINPUT40), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n847), .B2(new_n861), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n903), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n909), .A2(G330), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n830), .B1(new_n899), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n899), .B2(new_n912), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n205), .A2(new_n204), .A3(new_n531), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n459), .B(KEYINPUT99), .Z(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT35), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n918), .B2(new_n917), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT36), .Z(new_n921));
  INV_X1    g0721(.A(G58), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n922), .B2(new_n280), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n203), .B1(G50), .B2(new_n280), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n725), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n914), .A2(new_n921), .A3(new_n925), .ZN(G367));
  XOR2_X1   g0726(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n927));
  XOR2_X1   g0727(.A(new_n685), .B(new_n927), .Z(new_n928));
  OAI21_X1  g0728(.A(new_n676), .B1(new_n672), .B2(new_n675), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(new_n668), .ZN(new_n930));
  INV_X1    g0730(.A(new_n682), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n664), .B1(new_n498), .B2(new_n485), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n719), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n634), .A2(new_n664), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT44), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(KEYINPUT106), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n931), .B(new_n937), .C1(KEYINPUT106), .C2(new_n936), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT106), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(KEYINPUT44), .C1(new_n682), .C2(new_n935), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n682), .A2(new_n935), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT45), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT45), .B1(new_n682), .B2(new_n935), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n938), .B(new_n940), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n673), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n723), .B(new_n930), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(KEYINPUT107), .A3(new_n946), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n723), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n928), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n727), .A2(G1), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT104), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n935), .A2(new_n628), .A3(new_n675), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n499), .B1(new_n933), .B2(new_n671), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n959), .A2(KEYINPUT42), .B1(new_n665), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT42), .B2(new_n959), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n526), .A2(new_n665), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n524), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT101), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(KEYINPUT101), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n529), .A2(new_n963), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n962), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT102), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n958), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n970), .A2(KEYINPUT104), .A3(new_n973), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n946), .A2(new_n935), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT103), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n971), .B2(new_n974), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n970), .A2(KEYINPUT103), .A3(new_n973), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n982), .C1(new_n975), .C2(new_n976), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n978), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n957), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n769), .A2(new_n455), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n817), .A2(new_n556), .B1(new_n757), .B2(new_n804), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(G311), .C2(new_n768), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n752), .A2(KEYINPUT46), .A3(G116), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT46), .B1(new_n752), .B2(G116), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G107), .B2(new_n807), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n760), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n996), .B(new_n422), .C1(G294), .C2(new_n754), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n991), .A2(new_n992), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n807), .A2(G68), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n817), .B2(new_n275), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT108), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n754), .A2(G159), .B1(G77), .B2(new_n770), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G143), .A2(new_n768), .B1(new_n752), .B2(G58), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G50), .A2(new_n758), .B1(new_n761), .B2(G137), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n263), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n998), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT109), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n735), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n968), .A2(new_n785), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n737), .B1(new_n684), .B2(new_n364), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n227), .A2(new_n741), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n728), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n988), .A2(new_n1014), .ZN(G387));
  OR2_X1    g0815(.A1(new_n672), .A2(new_n785), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n224), .A2(G45), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n403), .A2(new_n286), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n687), .B(new_n244), .C1(new_n280), .C2(new_n313), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1017), .B(new_n741), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n687), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n739), .A2(new_n1022), .B1(new_n449), .B2(new_n684), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n737), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n817), .A2(new_n286), .B1(new_n767), .B2(new_n779), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G150), .B2(new_n761), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n989), .B1(G77), .B2(new_n752), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n754), .A2(new_n403), .B1(G68), .B2(new_n758), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n468), .B1(new_n807), .B2(new_n364), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT110), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n803), .A2(new_n810), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n817), .A2(new_n995), .B1(new_n757), .B2(new_n556), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G322), .C2(new_n768), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1034), .A2(KEYINPUT48), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(KEYINPUT48), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n773), .A2(new_n804), .B1(new_n751), .B2(new_n577), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT49), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n770), .A2(G116), .B1(new_n761), .B2(G326), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n468), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1038), .A2(KEYINPUT49), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1031), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n728), .B(new_n1024), .C1(new_n1043), .C2(new_n735), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n930), .A2(new_n955), .B1(new_n1016), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n723), .A2(new_n930), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n685), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n723), .A2(new_n930), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(G393));
  XNOR2_X1  g0849(.A(new_n941), .B(new_n942), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1050), .A2(new_n673), .A3(new_n940), .A4(new_n938), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT111), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n948), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n945), .A2(KEYINPUT111), .A3(new_n946), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n950), .A2(new_n951), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n685), .C1(new_n1056), .C2(new_n947), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n933), .A2(new_n734), .A3(new_n934), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n736), .B1(new_n455), .B2(new_n208), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n236), .B2(new_n741), .ZN(new_n1061));
  INV_X1    g0861(.A(G322), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n769), .A2(new_n449), .B1(new_n760), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n263), .B(new_n1063), .C1(G283), .C2(new_n752), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT113), .Z(new_n1065));
  AOI22_X1  g0865(.A1(new_n748), .A2(G311), .B1(new_n768), .B2(G317), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT52), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n807), .A2(G116), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n754), .A2(G303), .B1(G294), .B2(new_n758), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n754), .A2(G50), .B1(G68), .B2(new_n752), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n816), .B2(new_n760), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n817), .A2(new_n779), .B1(new_n767), .B2(new_n275), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1074));
  AOI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G87), .A2(new_n770), .B1(new_n758), .B2(new_n403), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n807), .A2(G77), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n422), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1065), .A2(new_n1070), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n728), .B(new_n1061), .C1(new_n1080), .C2(new_n735), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1058), .A2(new_n955), .B1(new_n1059), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1057), .A2(new_n1082), .ZN(G390));
  AOI21_X1  g0883(.A(new_n881), .B1(new_n885), .B2(new_n891), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n863), .A2(new_n872), .A3(KEYINPUT100), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n793), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n714), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n891), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n883), .B1(new_n721), .B2(new_n793), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n880), .B1(new_n1092), .B2(new_n892), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n847), .A2(new_n861), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1091), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1088), .A2(KEYINPUT114), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT114), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1084), .B1(new_n873), .B2(new_n879), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n1096), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1088), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n892), .A2(new_n1089), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n902), .A2(G330), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1098), .A2(new_n1101), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT115), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1092), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n795), .A2(new_n1107), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n892), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n892), .B1(new_n714), .B2(new_n1089), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1108), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1114), .A2(new_n1091), .B1(new_n1116), .B2(new_n885), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n448), .A2(new_n1107), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n897), .A2(new_n657), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1111), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n685), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1109), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT114), .B1(new_n1088), .B2(new_n1097), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1100), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1120), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT116), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1120), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n686), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT116), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1125), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n732), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n728), .B1(new_n272), .B2(new_n799), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n812), .A2(G125), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n751), .A2(new_n275), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n748), .A2(G132), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G50), .A2(new_n770), .B1(new_n758), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n754), .A2(G137), .B1(new_n768), .B2(G128), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n263), .C1(new_n779), .C2(new_n773), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n803), .A2(new_n449), .B1(new_n767), .B2(new_n804), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n817), .A2(new_n531), .B1(new_n757), .B2(new_n455), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n812), .A2(G294), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n823), .B(new_n263), .C1(G87), .C2(new_n752), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1078), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1148), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1135), .B1(new_n1156), .B2(new_n735), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1110), .A2(new_n955), .B1(new_n1133), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1127), .A2(new_n1132), .A3(new_n1158), .ZN(G378));
  NAND2_X1  g0959(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G50), .B1(new_n1160), .B2(new_n239), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT119), .Z(new_n1162));
  AOI22_X1  g0962(.A1(G97), .A2(new_n754), .B1(new_n748), .B2(G107), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n922), .B2(new_n769), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n511), .A2(new_n757), .B1(new_n531), .B2(new_n767), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n1165), .C1(G77), .C2(new_n752), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n468), .A3(new_n999), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1164), .B(new_n1167), .C1(G283), .C2(new_n812), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n1168), .B2(KEYINPUT58), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n768), .A2(G125), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n817), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G137), .A2(new_n758), .B1(new_n752), .B2(new_n1141), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n275), .B2(new_n773), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G132), .C2(new_n754), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n238), .B(new_n239), .C1(new_n769), .C2(new_n779), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G124), .B2(new_n761), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT59), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1169), .B1(KEYINPUT58), .B2(new_n1168), .C1(new_n1177), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n735), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT120), .Z(new_n1184));
  AOI211_X1 g0984(.A(new_n728), .B(new_n1184), .C1(new_n286), .C2(new_n799), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n298), .A2(new_n303), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n298), .B2(new_n303), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1188), .A2(new_n290), .A3(new_n834), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n290), .A2(new_n834), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1189), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n1187), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n732), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1185), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  INV_X1    g0998(.A(G330), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n906), .A2(new_n1199), .A3(new_n908), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1198), .B1(new_n1200), .B2(new_n1194), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n907), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1094), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n904), .B1(new_n871), .B2(new_n847), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(G330), .C1(KEYINPUT40), .C2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1205), .A2(new_n1195), .A3(KEYINPUT122), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1205), .A2(KEYINPUT121), .A3(new_n1195), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT121), .B1(new_n1205), .B2(new_n1195), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1201), .A2(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n896), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1200), .A2(new_n1198), .A3(new_n1194), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT122), .B1(new_n1205), .B2(new_n1195), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n896), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n1208), .C2(new_n1207), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1197), .B1(new_n1216), .B2(new_n956), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1117), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1122), .B(new_n1218), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1119), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n686), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1222), .A3(KEYINPUT57), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1217), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n928), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n892), .A2(new_n732), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n729), .B1(G68), .B2(new_n800), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G77), .A2(new_n770), .B1(new_n752), .B2(G97), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n255), .C1(new_n511), .C2(new_n773), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n754), .A2(G116), .B1(G107), .B2(new_n758), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n748), .A2(G283), .B1(new_n768), .B2(G294), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n764), .C2(new_n556), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n754), .A2(new_n1141), .B1(G150), .B2(new_n758), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n748), .A2(G137), .B1(new_n768), .B2(G132), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n764), .C2(new_n1171), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G58), .A2(new_n770), .B1(new_n752), .B2(G159), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n422), .C1(new_n286), .C2(new_n773), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1235), .A2(new_n1238), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1233), .B1(new_n1244), .B2(new_n735), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1218), .A2(new_n955), .B1(new_n1232), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1231), .A2(new_n1246), .ZN(G381));
  OAI21_X1  g1047(.A(new_n1158), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1057), .A2(new_n1082), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n988), .A2(new_n1249), .A3(new_n1014), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G375), .A2(new_n1248), .A3(new_n1250), .A4(new_n1251), .ZN(G407));
  INV_X1    g1052(.A(new_n1248), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n663), .A2(G213), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1227), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(G213), .A3(new_n1256), .ZN(G409));
  AOI21_X1  g1057(.A(new_n986), .B1(new_n954), .B2(new_n956), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1014), .ZN(new_n1259));
  OAI21_X1  g1059(.A(G390), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(G393), .B(new_n787), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1250), .A2(new_n1260), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1250), .B2(new_n1260), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1222), .A2(new_n955), .B1(new_n1196), .B2(new_n1185), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1221), .A2(new_n1222), .A3(new_n928), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1248), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1227), .B2(G378), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1230), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n1119), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1229), .A3(new_n685), .A4(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(G384), .A3(new_n1246), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT123), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1246), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n798), .A3(new_n828), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(KEYINPUT123), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1270), .A2(KEYINPUT124), .A3(new_n1255), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1119), .B1(new_n1110), .B2(new_n1218), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1224), .B1(new_n1216), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n685), .A3(new_n1226), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(G378), .A3(new_n1267), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1269), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1255), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1280), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1282), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1281), .A2(new_n1290), .A3(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1254), .A3(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1255), .A2(G2897), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .A4(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1280), .A2(G2897), .A3(new_n1255), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1297), .B(new_n1298), .C1(new_n1270), .C2(new_n1255), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(new_n1295), .A3(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1266), .B1(new_n1291), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(KEYINPUT124), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1288), .A2(new_n1282), .A3(new_n1289), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT63), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1254), .A4(new_n1289), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1299), .A2(new_n1306), .A3(new_n1295), .A4(new_n1265), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1281), .B2(new_n1290), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1298), .A2(new_n1297), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1265), .B(new_n1295), .C1(new_n1288), .C2(new_n1311), .ZN(new_n1312));
  NOR4_X1   g1112(.A1(new_n1270), .A2(new_n1309), .A3(new_n1255), .A4(new_n1280), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT125), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1301), .B1(new_n1308), .B2(new_n1315), .ZN(G405));
  OAI21_X1  g1116(.A(new_n1286), .B1(new_n1227), .B2(new_n1248), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT126), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT127), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1317), .A2(KEYINPUT126), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1265), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1317), .A2(KEYINPUT126), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1266), .A3(new_n1321), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1323), .A2(new_n1289), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1289), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1319), .A2(new_n1266), .A3(new_n1321), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1266), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1327), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1326), .A2(new_n1330), .ZN(G402));
endmodule


