//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n187), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n193), .B2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(KEYINPUT73), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT73), .B1(new_n197), .B2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(KEYINPUT23), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G110), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n195), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n202), .A2(KEYINPUT74), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT74), .B1(new_n202), .B2(new_n205), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(G146), .B(new_n211), .C1(new_n215), .C2(new_n209), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT75), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  XNOR2_X1  g033(.A(G125), .B(G140), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n211), .B1(new_n215), .B2(new_n209), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n221), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n226), .A2(new_n216), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n196), .A2(new_n200), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n228), .A2(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n192), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n232), .B(new_n191), .C1(new_n208), .C2(new_n223), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  AOI21_X1  g048(.A(G902), .B1(new_n234), .B2(KEYINPUT76), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(KEYINPUT76), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n231), .A2(new_n233), .A3(new_n239), .A4(new_n235), .ZN(new_n240));
  OAI21_X1  g054(.A(G217), .B1(new_n189), .B2(G902), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT72), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(new_n233), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT31), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT2), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G116), .B(G119), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n257), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n221), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT0), .A4(G128), .ZN(new_n265));
  XNOR2_X1  g079(.A(G143), .B(G146), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G137), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(G134), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n269), .C2(G134), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n273), .B(new_n281), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n268), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n263), .B(G146), .C1(new_n193), .C2(KEYINPUT1), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n193), .A2(new_n221), .A3(G143), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n262), .A3(new_n264), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n269), .A3(G134), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n272), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n282), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n283), .A2(new_n295), .A3(KEYINPUT30), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n297));
  INV_X1    g111(.A(new_n268), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n270), .A2(new_n272), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n276), .B1(new_n271), .B2(G137), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT64), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n275), .A2(new_n274), .A3(new_n276), .ZN(new_n302));
  AOI211_X1 g116(.A(G131), .B(new_n299), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n281), .B1(new_n304), .B2(new_n273), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n298), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n282), .A2(new_n289), .A3(new_n294), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n261), .B1(new_n296), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n261), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G101), .ZN(new_n312));
  NOR2_X1   g126(.A1(G237), .A2(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G210), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n312), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n309), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT67), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n283), .A2(new_n295), .A3(new_n261), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT30), .B1(new_n283), .B2(new_n295), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n306), .A2(new_n297), .A3(new_n307), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n323), .B2(new_n261), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT67), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n317), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n250), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(new_n250), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n310), .B1(new_n306), .B2(new_n307), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n320), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n311), .A2(KEYINPUT68), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n317), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT69), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n336), .A2(KEYINPUT69), .A3(new_n337), .ZN(new_n339));
  OAI22_X1  g153(.A1(new_n327), .A2(new_n329), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(G472), .A2(G902), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT70), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n310), .B1(new_n321), .B2(new_n322), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n337), .B1(new_n346), .B2(new_n320), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(new_n347), .C1(new_n336), .C2(new_n337), .ZN(new_n348));
  INV_X1    g162(.A(new_n335), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT68), .B1(new_n311), .B2(new_n334), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n337), .A2(new_n345), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n261), .B1(new_n283), .B2(new_n295), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n334), .B1(new_n353), .B2(new_n311), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n354), .A2(KEYINPUT71), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(KEYINPUT71), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n351), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n357), .A3(new_n245), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n340), .A2(new_n344), .B1(G472), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n325), .B1(new_n324), .B2(new_n317), .ZN(new_n360));
  NOR4_X1   g174(.A1(new_n346), .A2(KEYINPUT67), .A3(new_n320), .A4(new_n337), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT31), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n349), .A2(new_n354), .A3(new_n350), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(new_n317), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n336), .A2(KEYINPUT69), .A3(new_n337), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n362), .A2(new_n328), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n343), .B1(new_n367), .B2(new_n342), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n249), .B1(new_n359), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G140), .ZN(new_n370));
  INV_X1    g184(.A(G953), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G227), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n370), .B(new_n372), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n288), .A2(KEYINPUT78), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n266), .A2(new_n375), .A3(new_n287), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n286), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(G107), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  XNOR2_X1  g200(.A(G104), .B(G107), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n383), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n378), .A2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n381), .A2(G104), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT77), .B(G101), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n377), .A2(new_n385), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n379), .A2(new_n382), .A3(new_n384), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n383), .A2(new_n396), .B1(new_n388), .B2(new_n391), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n286), .B2(new_n288), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n393), .A2(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n280), .A2(new_n282), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n395), .A2(new_n404), .A3(G101), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n298), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n399), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n401), .B1(new_n399), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n373), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n377), .A2(new_n385), .A3(new_n392), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n289), .B1(new_n392), .B2(new_n385), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n400), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT12), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n373), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n393), .B1(new_n289), .B2(new_n397), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT79), .A3(new_n413), .A4(new_n400), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n399), .A2(new_n401), .A3(new_n406), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n416), .A2(new_n417), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n409), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n245), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n416), .A2(new_n420), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n373), .ZN(new_n426));
  INV_X1    g240(.A(new_n408), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n417), .A3(new_n420), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(G469), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G469), .A2(G902), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT9), .B(G234), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n188), .B1(new_n433), .B2(new_n245), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n268), .A2(G125), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n286), .A2(new_n213), .A3(new_n288), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G224), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G953), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n441), .B(new_n443), .Z(new_n444));
  NAND3_X1  g258(.A1(new_n403), .A2(new_n261), .A3(new_n405), .ZN(new_n445));
  INV_X1    g259(.A(G116), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(G119), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n251), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n197), .A2(G116), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(G119), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT5), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n449), .A2(new_n452), .B1(new_n257), .B2(new_n255), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n392), .A2(new_n453), .A3(new_n385), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n445), .A2(new_n454), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n455), .B(KEYINPUT80), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n444), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n455), .B(KEYINPUT8), .Z(new_n464));
  AOI21_X1  g278(.A(new_n453), .B1(new_n392), .B2(new_n385), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n392), .A2(new_n385), .A3(new_n453), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(KEYINPUT81), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n454), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n441), .B1(new_n471), .B2(new_n443), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n443), .A2(new_n471), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n439), .A2(new_n440), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n456), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n245), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n438), .B1(new_n463), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n475), .ZN(new_n478));
  INV_X1    g292(.A(new_n464), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n392), .A2(new_n385), .ZN(new_n480));
  INV_X1    g294(.A(new_n453), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n468), .B2(new_n454), .ZN(new_n483));
  INV_X1    g297(.A(new_n469), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n441), .B(new_n443), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n456), .A2(KEYINPUT6), .B1(new_n458), .B2(new_n459), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n490), .A3(new_n437), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n477), .A2(KEYINPUT82), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G214), .B1(G237), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT82), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n486), .A2(new_n490), .A3(new_n494), .A4(new_n437), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G122), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n497), .B2(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n446), .A2(G122), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT14), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(G116), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT86), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n446), .A3(G122), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n446), .B2(G122), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n508), .A2(new_n501), .B1(G116), .B2(new_n497), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT86), .B1(new_n509), .B2(new_n499), .ZN(new_n510));
  OAI21_X1  g324(.A(G107), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n263), .A2(G128), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n193), .A2(G143), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G134), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n513), .A3(new_n271), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n500), .A2(new_n503), .A3(new_n381), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n520));
  INV_X1    g334(.A(new_n518), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n381), .B1(new_n500), .B2(new_n503), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n263), .A2(G128), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n512), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n263), .A2(KEYINPUT13), .A3(G128), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n271), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n520), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n522), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n518), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n512), .A2(new_n525), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n513), .A3(new_n527), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G134), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT84), .A4(new_n516), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n433), .A2(G217), .A3(new_n371), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n519), .A2(new_n529), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n517), .A2(new_n518), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n502), .A2(new_n503), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n508), .A2(new_n501), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n506), .A3(new_n504), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n539), .B1(new_n544), .B2(G107), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n529), .A2(new_n535), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n536), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT87), .B1(new_n548), .B2(new_n245), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n550), .B(G902), .C1(new_n538), .C2(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n549), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n245), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n553), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n371), .A2(G952), .ZN(new_n560));
  NAND2_X1  g374(.A1(G234), .A2(G237), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(G902), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n313), .A2(G143), .A3(G214), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(G143), .B1(new_n313), .B2(G214), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT18), .B(G131), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n215), .A2(G146), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n222), .ZN(new_n574));
  INV_X1    g388(.A(new_n571), .ZN(new_n575));
  NAND2_X1  g389(.A1(KEYINPUT18), .A2(G131), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n579));
  OAI21_X1  g393(.A(G131), .B1(new_n570), .B2(new_n571), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n226), .B(new_n216), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n575), .A2(new_n281), .A3(new_n569), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n580), .A2(new_n582), .A3(new_n579), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n578), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(G113), .B(G122), .Z(new_n585));
  XOR2_X1   g399(.A(KEYINPUT83), .B(G104), .Z(new_n586));
  XOR2_X1   g400(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n578), .B(new_n587), .C1(new_n581), .C2(new_n583), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G475), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT20), .ZN(new_n594));
  INV_X1    g408(.A(new_n578), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n216), .B(KEYINPUT75), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n220), .B(KEYINPUT19), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n597), .A2(new_n221), .B1(new_n580), .B2(new_n582), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n595), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n590), .B1(new_n599), .B2(new_n587), .ZN(new_n600));
  NOR2_X1   g414(.A1(G475), .A2(G902), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n594), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n594), .A3(new_n601), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n593), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n558), .A2(new_n559), .A3(new_n568), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n556), .A2(new_n550), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n548), .A2(KEYINPUT87), .A3(new_n245), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n553), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n557), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n568), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT88), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n496), .B1(new_n606), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n369), .A2(new_n436), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  INV_X1    g430(.A(KEYINPUT89), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n367), .B2(G902), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n340), .A2(KEYINPUT89), .A3(new_n245), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(G472), .ZN(new_n620));
  INV_X1    g434(.A(new_n342), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n340), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n249), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n436), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n607), .A2(new_n552), .A3(new_n608), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n548), .A2(KEYINPUT33), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n538), .B2(new_n547), .ZN(new_n630));
  OAI211_X1 g444(.A(G478), .B(new_n245), .C1(new_n628), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n605), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n493), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n477), .B2(new_n491), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n633), .A2(new_n567), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  OAI21_X1  g455(.A(new_n604), .B1(new_n602), .B2(KEYINPUT91), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT91), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n600), .A2(new_n643), .A3(new_n594), .A4(new_n601), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n593), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n611), .A2(new_n568), .A3(new_n635), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n626), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(KEYINPUT92), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n208), .A2(new_n223), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n232), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n224), .A2(KEYINPUT92), .A3(new_n230), .ZN(new_n653));
  OAI22_X1  g467(.A1(new_n652), .A2(new_n653), .B1(KEYINPUT36), .B2(new_n192), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n651), .A2(new_n650), .A3(new_n232), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT92), .B1(new_n224), .B2(new_n230), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n654), .A2(new_n247), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n244), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT93), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n244), .A2(new_n659), .A3(KEYINPUT93), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n435), .A2(new_n662), .A3(new_n431), .A4(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n620), .A2(new_n614), .A3(new_n664), .A4(new_n622), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n359), .A2(new_n368), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n371), .A2(G900), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(G902), .A3(new_n561), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT94), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(KEYINPUT94), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n562), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n593), .B(new_n674), .C1(new_n642), .C2(new_n644), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n611), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n668), .A2(new_n664), .A3(new_n635), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n673), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n436), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n682));
  INV_X1    g496(.A(new_n604), .ZN(new_n683));
  OAI22_X1  g497(.A1(new_n683), .A2(new_n602), .B1(new_n592), .B2(new_n591), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n555), .B2(new_n557), .ZN(new_n685));
  INV_X1    g499(.A(new_n660), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n493), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n681), .A2(new_n682), .A3(new_n685), .A4(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n317), .B1(new_n353), .B2(new_n311), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT96), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(G472), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n689), .B2(new_n690), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n319), .A2(new_n326), .A3(new_n691), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(G472), .A2(G902), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n694), .A2(KEYINPUT97), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT97), .B1(new_n694), .B2(new_n695), .ZN(new_n697));
  INV_X1    g511(.A(new_n344), .ZN(new_n698));
  OAI22_X1  g512(.A1(new_n696), .A2(new_n697), .B1(new_n367), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT32), .B1(new_n340), .B2(new_n621), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n492), .A2(new_n495), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n688), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR2_X1   g521(.A1(new_n633), .A2(new_n674), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n668), .A2(new_n664), .A3(new_n635), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT98), .B(G146), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G48));
  INV_X1    g525(.A(new_n424), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n423), .B1(new_n422), .B2(new_n245), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n435), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n369), .A2(new_n637), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT99), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n717), .B(new_n719), .ZN(G15));
  NAND3_X1  g534(.A1(new_n369), .A2(new_n646), .A3(new_n716), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NOR2_X1   g536(.A1(new_n715), .A2(new_n636), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n606), .A2(new_n613), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n662), .A2(new_n663), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n668), .A2(new_n723), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT100), .B(G119), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G21));
  NAND2_X1  g542(.A1(new_n319), .A2(new_n326), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n329), .B1(new_n729), .B2(KEYINPUT31), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n339), .A2(new_n338), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n245), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n337), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n327), .B2(new_n329), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n732), .A2(G472), .B1(new_n735), .B2(new_n621), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT101), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n685), .B2(new_n636), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n611), .A2(KEYINPUT101), .A3(new_n684), .A4(new_n635), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n715), .A2(new_n567), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n736), .A2(new_n740), .A3(new_n624), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND4_X1  g557(.A1(new_n736), .A2(new_n723), .A3(new_n660), .A4(new_n708), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  XOR2_X1   g559(.A(new_n430), .B(KEYINPUT102), .Z(new_n746));
  NAND3_X1  g560(.A1(new_n424), .A2(new_n429), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n435), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n747), .B2(new_n435), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n703), .A2(new_n493), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n668), .A3(new_n624), .A4(new_n708), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n358), .A2(G472), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n367), .B2(new_n698), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n624), .B1(new_n700), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n750), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n634), .B1(new_n492), .B2(new_n495), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n747), .A2(new_n748), .A3(new_n435), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT105), .A3(KEYINPUT42), .A4(new_n708), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n369), .A2(KEYINPUT42), .A3(new_n708), .A4(new_n752), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n756), .A2(new_n758), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n281), .ZN(G33));
  NAND3_X1  g586(.A1(new_n369), .A2(new_n676), .A3(new_n752), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NOR2_X1   g588(.A1(new_n623), .A2(new_n686), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT108), .Z(new_n776));
  OR2_X1    g590(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n627), .A2(new_n631), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT43), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n782), .A3(new_n605), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n776), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n776), .A2(KEYINPUT44), .A3(new_n785), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n426), .A2(new_n428), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT45), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(G469), .C1(KEYINPUT45), .C2(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n746), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n746), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n424), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n435), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n679), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n751), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n788), .A2(new_n789), .A3(new_n803), .ZN(new_n804));
  XOR2_X1   g618(.A(KEYINPUT109), .B(G137), .Z(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G39));
  NAND3_X1  g620(.A1(new_n708), .A2(new_n249), .A3(new_n763), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n668), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n799), .A2(new_n435), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n799), .B2(new_n435), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT111), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NAND4_X1  g628(.A1(new_n717), .A2(new_n721), .A3(new_n726), .A4(new_n742), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n753), .A2(new_n757), .A3(new_n754), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n757), .B1(new_n753), .B2(new_n754), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n768), .B(KEYINPUT105), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n677), .A2(new_n744), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n435), .A2(new_n686), .A3(new_n673), .A4(new_n747), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n740), .B(new_n824), .C1(new_n699), .C2(new_n700), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n823), .A3(new_n709), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n684), .B1(new_n609), .B2(new_n610), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n568), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n568), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n605), .B1(new_n555), .B2(new_n557), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT112), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n568), .A3(new_n632), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n830), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n622), .A3(new_n620), .A4(new_n625), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n615), .A3(new_n665), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n752), .A2(new_n736), .A3(new_n660), .A4(new_n708), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n675), .A2(new_n558), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n839), .B1(new_n840), .B2(new_n751), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n763), .A2(new_n675), .A3(KEYINPUT113), .A4(new_n558), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n668), .A2(new_n664), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n773), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n677), .A2(new_n709), .A3(new_n825), .A4(new_n744), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n826), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n677), .A2(new_n744), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n849), .B2(KEYINPUT52), .ZN(new_n850));
  OR3_X1    g664(.A1(new_n821), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n821), .B2(new_n848), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n771), .B2(new_n815), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n852), .B1(new_n849), .B2(KEYINPUT52), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n826), .A2(new_n845), .A3(new_n847), .A4(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT114), .B(new_n816), .C1(new_n819), .C2(new_n820), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n853), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n784), .A2(new_n562), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n624), .A3(new_n736), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n810), .A2(new_n811), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n714), .A2(new_n434), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n751), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n715), .A2(new_n493), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT115), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n866), .A2(new_n871), .A3(new_n705), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT50), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n715), .A2(new_n751), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n701), .A2(new_n624), .A3(new_n563), .A4(new_n874), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n875), .A2(new_n684), .A3(new_n778), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n736), .A2(new_n660), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n865), .A2(new_n874), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT116), .Z(new_n879));
  OAI211_X1 g693(.A(new_n873), .B(new_n876), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n869), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n869), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n761), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT48), .ZN(new_n885));
  INV_X1    g699(.A(new_n723), .ZN(new_n886));
  OAI221_X1 g700(.A(new_n560), .B1(new_n875), .B2(new_n633), .C1(new_n866), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n864), .A2(new_n882), .A3(new_n883), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(G952), .B2(G953), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n780), .A2(new_n249), .A3(new_n434), .A4(new_n634), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n714), .B(KEYINPUT49), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n701), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n705), .B2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n371), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n245), .B1(new_n861), .B2(new_n853), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(G210), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n488), .A2(new_n489), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n487), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n896), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n898), .B2(new_n901), .ZN(G51));
  XNOR2_X1  g717(.A(new_n862), .B(KEYINPUT54), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n746), .B(KEYINPUT57), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n422), .ZN(new_n907));
  INV_X1    g721(.A(new_n794), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n895), .B1(new_n907), .B2(new_n909), .ZN(G54));
  AND3_X1   g724(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n896), .B1(new_n911), .B2(new_n600), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n600), .B2(new_n911), .ZN(G60));
  NOR2_X1   g727(.A1(new_n628), .A2(new_n630), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n904), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT117), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n904), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n914), .B1(new_n864), .B2(new_n916), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n896), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n922), .A2(KEYINPUT118), .A3(new_n896), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT120), .B1(new_n862), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n933), .B(new_n930), .C1(new_n861), .C2(new_n853), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n231), .A2(new_n233), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n895), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n654), .A2(new_n658), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n932), .B2(new_n934), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT121), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n938), .C1(new_n932), .C2(new_n934), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT123), .B1(new_n935), .B2(new_n936), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n935), .A2(KEYINPUT123), .A3(new_n936), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT124), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n862), .A2(new_n931), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n933), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n862), .A2(KEYINPUT120), .A3(new_n931), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n949), .B1(new_n958), .B2(new_n938), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n936), .A3(new_n957), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND4_X1   g776(.A1(KEYINPUT124), .A2(new_n959), .A3(new_n953), .A4(new_n962), .ZN(new_n963));
  OAI22_X1  g777(.A1(new_n946), .A2(new_n947), .B1(new_n954), .B2(new_n963), .ZN(G66));
  OAI21_X1  g778(.A(G953), .B1(new_n566), .B2(new_n442), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n815), .A2(new_n837), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n899), .B1(G898), .B2(new_n371), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  XOR2_X1   g783(.A(new_n597), .B(KEYINPUT125), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n323), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n822), .A2(new_n709), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n773), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n369), .A2(new_n740), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT127), .B1(new_n802), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n801), .A2(new_n977), .A3(new_n679), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n771), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n813), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(G953), .B1(new_n982), .B2(new_n804), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n971), .B1(new_n983), .B2(new_n669), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n973), .A2(new_n706), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT62), .Z(new_n986));
  AOI21_X1  g800(.A(new_n680), .B1(new_n633), .B2(new_n832), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n369), .A3(new_n763), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n813), .A2(new_n804), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n971), .B1(new_n989), .B2(new_n371), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n371), .B1(G227), .B2(G900), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G72));
  NAND3_X1  g809(.A1(new_n982), .A2(new_n804), .A3(new_n966), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n695), .B(KEYINPUT63), .Z(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n324), .A3(new_n337), .ZN(new_n999));
  INV_X1    g813(.A(new_n966), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n997), .B1(new_n989), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n1001), .B(new_n317), .C1(new_n320), .C2(new_n346), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n319), .A2(new_n326), .A3(new_n347), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1003), .A2(new_n997), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n895), .B1(new_n854), .B2(new_n1004), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n999), .A2(new_n1002), .A3(new_n1005), .ZN(G57));
endmodule


