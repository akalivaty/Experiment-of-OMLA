//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n466), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G2105), .B1(new_n469), .B2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  AND2_X1   g047(.A1(new_n463), .A2(new_n465), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n466), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n478), .A2(G124), .B1(G136), .B2(new_n469), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n476), .B2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND3_X1  g058(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .ZN(new_n484));
  NAND2_X1  g059(.A1(G102), .A2(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n476), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n463), .A2(new_n465), .A3(G126), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n476), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n473), .A2(new_n476), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n505), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n502), .A2(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n500), .A2(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT68), .B(G51), .ZN(new_n518));
  OAI221_X1 g093(.A(new_n516), .B1(new_n510), .B2(new_n517), .C1(new_n502), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n497), .A2(G63), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n499), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G168));
  NAND2_X1  g098(.A1(new_n505), .A2(new_n507), .ZN(new_n524));
  INV_X1    g099(.A(G64), .ZN(new_n525));
  INV_X1    g100(.A(G77), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n504), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n529), .B1(new_n526), .B2(new_n504), .C1(new_n524), .C2(new_n525), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(G651), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n502), .A2(new_n532), .B1(new_n510), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n499), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n502), .A2(new_n539), .B1(new_n510), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT70), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  NOR2_X1   g124(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n497), .B2(new_n501), .ZN(new_n552));
  OAI21_X1  g127(.A(G91), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT71), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n504), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n559), .A2(KEYINPUT71), .A3(new_n560), .A4(G53), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n524), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n553), .A2(new_n562), .A3(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n531), .A2(new_n535), .ZN(G301));
  OR2_X1    g143(.A1(new_n519), .A2(new_n522), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n497), .A2(new_n501), .A3(new_n551), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G87), .B1(G49), .B2(new_n559), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n573), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n524), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n559), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n499), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n502), .A2(new_n585), .B1(new_n510), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n573), .B2(G92), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  AOI211_X1 g168(.A(KEYINPUT10), .B(new_n593), .C1(new_n571), .C2(new_n572), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n524), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n559), .A2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g177(.A1(new_n592), .A2(new_n594), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G299), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(G168), .ZN(G297));
  XNOR2_X1  g183(.A(G297), .B(KEYINPUT74), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n473), .A2(new_n459), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n476), .A2(G111), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT75), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n469), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G123), .B2(new_n478), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2435), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2438), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2451), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XNOR2_X1  g217(.A(G2084), .B(G2090), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT77), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  INV_X1    g224(.A(new_n644), .ZN(new_n650));
  INV_X1    g225(.A(new_n645), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n650), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n647), .B(KEYINPUT17), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n644), .B2(new_n645), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n652), .A2(new_n654), .A3(new_n646), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT78), .B(G1981), .Z(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT79), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  NAND2_X1  g255(.A1(G171), .A2(G16), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G5), .B2(G16), .ZN(new_n682));
  INV_X1    g257(.A(G1961), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G11), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT30), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(G28), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(G28), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n684), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n692));
  NOR2_X1   g267(.A1(G16), .A2(G21), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G168), .B2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1966), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n625), .A2(G29), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n691), .A2(new_n692), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n684), .A2(new_n697), .A3(new_n685), .A4(new_n690), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT86), .B1(new_n699), .B2(new_n695), .ZN(new_n700));
  INV_X1    g275(.A(G2072), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n473), .A2(G139), .A3(new_n476), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n459), .A2(G103), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(KEYINPUT82), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n459), .A2(new_n707), .A3(G103), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n706), .A2(new_n708), .A3(KEYINPUT25), .ZN(new_n709));
  AOI21_X1  g284(.A(KEYINPUT25), .B1(new_n706), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(new_n476), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n704), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G29), .B2(G33), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n698), .A2(new_n700), .B1(new_n701), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n689), .A2(G26), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n478), .A2(G128), .B1(G140), .B2(new_n469), .ZN(new_n720));
  OR2_X1    g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n689), .ZN(new_n725));
  MUX2_X1   g300(.A(new_n719), .B(new_n725), .S(KEYINPUT28), .Z(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(G2067), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n689), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n689), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2090), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n726), .A2(G2067), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n542), .B2(new_n734), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1341), .Z(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(KEYINPUT23), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n718), .A2(new_n733), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n603), .B2(G16), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n730), .A2(G2090), .B1(G1348), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(G164), .A2(G29), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G27), .B2(G29), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n743), .A2(new_n746), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G32), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n478), .B2(G129), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n459), .A2(G105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n759));
  INV_X1    g334(.A(G141), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n492), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n469), .A2(KEYINPUT84), .A3(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT85), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n757), .A2(new_n763), .A3(new_n766), .A4(new_n758), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n754), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT27), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1996), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n745), .A2(G1348), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n717), .B2(new_n701), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G34), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n471), .B2(G29), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n682), .A2(new_n683), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n753), .A2(new_n772), .A3(new_n775), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n734), .A2(G23), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G288), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT81), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n734), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n734), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G6), .B(G305), .S(G16), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n789), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n478), .A2(G119), .B1(G131), .B2(new_n469), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G25), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT80), .B1(new_n806), .B2(G29), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n806), .A2(KEYINPUT80), .A3(G29), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT35), .B(G1991), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G24), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n588), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1986), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n799), .A2(new_n800), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n800), .B1(new_n799), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n782), .A2(new_n776), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n784), .A2(new_n818), .A3(new_n819), .ZN(G311));
  AND3_X1   g395(.A1(new_n753), .A2(new_n775), .A3(new_n783), .ZN(new_n821));
  INV_X1    g396(.A(new_n818), .ZN(new_n822));
  INV_X1    g397(.A(new_n819), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n772), .ZN(G150));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n502), .A2(new_n825), .B1(new_n510), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n497), .A2(G67), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n499), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  OAI21_X1  g410(.A(G92), .B1(new_n550), .B2(new_n552), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT10), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n597), .B(KEYINPUT73), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n595), .B2(new_n524), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n839), .A2(G651), .B1(G54), .B2(new_n559), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n573), .A2(new_n591), .A3(G92), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n610), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT88), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n828), .A2(new_n832), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT88), .B1(new_n827), .B2(new_n831), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n542), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n542), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n845), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n835), .B1(new_n854), .B2(G860), .ZN(G145));
  NAND2_X1  g430(.A1(new_n768), .A2(G164), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n765), .A2(new_n495), .A3(new_n767), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n723), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n724), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n715), .A2(KEYINPUT90), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n617), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n804), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n478), .A2(G130), .B1(G142), .B2(new_n469), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n476), .A2(G118), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G2104), .ZN(new_n867));
  NOR2_X1   g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT89), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n704), .A2(new_n711), .A3(new_n871), .A4(new_n713), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT90), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n864), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n804), .B(new_n617), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n862), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n883), .A2(new_n861), .A3(new_n860), .A4(new_n859), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT91), .ZN(new_n885));
  XNOR2_X1  g460(.A(G162), .B(new_n625), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT91), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G160), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(G160), .A3(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g470(.A(G299), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n842), .A2(KEYINPUT93), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT93), .B1(new_n842), .B2(new_n896), .ZN(new_n898));
  NAND4_X1  g473(.A1(G299), .A2(new_n837), .A3(new_n840), .A4(new_n841), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT94), .B1(new_n901), .B2(KEYINPUT41), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT94), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT93), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n603), .B2(G299), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n842), .A2(KEYINPUT93), .A3(new_n896), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n903), .B(new_n904), .C1(new_n908), .C2(new_n900), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT95), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT92), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n592), .A2(new_n594), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(KEYINPUT92), .A3(G299), .A4(new_n840), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n906), .A2(new_n907), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n911), .B1(new_n916), .B2(new_n904), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n913), .A2(new_n915), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n897), .A2(new_n898), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT95), .A4(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n853), .B(new_n612), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n916), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(KEYINPUT97), .A2(KEYINPUT42), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G288), .B(G290), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT96), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT96), .ZN(new_n932));
  INV_X1    g507(.A(G288), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(G290), .ZN(new_n934));
  NOR2_X1   g509(.A1(G288), .A2(new_n588), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(G303), .B(G305), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(KEYINPUT96), .A3(new_n930), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(KEYINPUT97), .B2(KEYINPUT42), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n924), .B(new_n926), .C1(KEYINPUT97), .C2(KEYINPUT42), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n929), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n929), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n833), .A2(new_n606), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  XOR2_X1   g525(.A(KEYINPUT98), .B(KEYINPUT44), .Z(new_n951));
  XNOR2_X1  g526(.A(G286), .B(G301), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n853), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n847), .A2(new_n542), .A3(new_n848), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n542), .B1(new_n847), .B2(new_n848), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(G301), .B(G168), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n910), .B2(new_n921), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n952), .B2(new_n853), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT99), .B1(new_n956), .B2(new_n957), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT99), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n952), .A2(new_n853), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT100), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n963), .A2(new_n964), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n925), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT101), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n938), .A2(KEYINPUT102), .A3(new_n940), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT102), .B1(new_n938), .B2(new_n940), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n968), .A2(new_n925), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n902), .A2(new_n909), .B1(new_n917), .B2(new_n920), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n960), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n969), .B1(new_n922), .B2(new_n959), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n979), .B2(new_n941), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT41), .B1(new_n908), .B2(new_n900), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n968), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n916), .A2(KEYINPUT41), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n983), .A2(new_n984), .B1(new_n925), .B2(new_n959), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n973), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n974), .B(new_n941), .C1(new_n976), .C2(new_n960), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n892), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n981), .A2(KEYINPUT43), .B1(KEYINPUT103), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n991), .B(new_n988), .C1(new_n978), .C2(new_n980), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n951), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n980), .A2(new_n986), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT104), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n980), .A2(new_n996), .A3(new_n986), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(KEYINPUT43), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT44), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n993), .B1(new_n999), .B2(new_n1000), .ZN(G397));
  AOI21_X1  g576(.A(G1384), .B1(new_n487), .B2(new_n494), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n461), .A2(new_n470), .A3(G40), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G1996), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n769), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1008), .A2(KEYINPUT105), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(KEYINPUT105), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1006), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n723), .B(G2067), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n768), .A3(G1996), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT106), .Z(new_n1015));
  NOR2_X1   g590(.A1(new_n804), .A2(new_n810), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n804), .A2(new_n810), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT125), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OR2_X1    g597(.A1(G290), .A2(G1986), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1006), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT48), .Z(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1013), .A2(new_n1016), .A3(new_n1015), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(G2067), .B2(new_n723), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1011), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1011), .B1(new_n1012), .B2(new_n768), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT124), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1026), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1005), .A2(new_n1002), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  INV_X1    g616(.A(G86), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n581), .B1(new_n1042), .B2(new_n510), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1041), .B1(G1981), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT49), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(KEYINPUT49), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n1040), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(G288), .A2(G1976), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT113), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1040), .B1(new_n1053), .B2(new_n1041), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1040), .B1(new_n1056), .B2(G288), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(KEYINPUT110), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1057), .B(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(G288), .A2(new_n1058), .A3(new_n1056), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1064), .B(G1384), .C1(new_n487), .C2(new_n494), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1003), .A2(new_n1065), .A3(new_n1004), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1066), .A2(G1966), .ZN(new_n1067));
  INV_X1    g642(.A(G1384), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n495), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1004), .B1(new_n1069), .B2(KEYINPUT50), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1002), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n776), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1039), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G168), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G303), .A2(G8), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1076), .B(KEYINPUT55), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1069), .A2(KEYINPUT50), .ZN(new_n1078));
  INV_X1    g653(.A(G2090), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1005), .A4(new_n1072), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT108), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT108), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1070), .A2(new_n1082), .A3(new_n1079), .A4(new_n1072), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1069), .A2(new_n1064), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1005), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n792), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1081), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1077), .B1(new_n1088), .B2(G8), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1063), .A2(new_n1075), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1054), .B1(new_n1055), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1037), .A2(G2067), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1078), .A2(new_n1005), .A3(new_n1072), .ZN(new_n1093));
  INV_X1    g668(.A(G1348), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n842), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1072), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1005), .B1(new_n1002), .B2(new_n1071), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1092), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1099), .A2(new_n1100), .A3(KEYINPUT60), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1096), .B1(new_n1103), .B2(new_n603), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1002), .A2(new_n1106), .A3(new_n1071), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1002), .B2(new_n1071), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1070), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1110), .A2(new_n1111), .B1(new_n1066), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G299), .B(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1105), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT58), .B(G1341), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1086), .A2(G1996), .B1(new_n1038), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(KEYINPUT118), .A3(new_n542), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT59), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1120), .A2(KEYINPUT118), .A3(new_n1123), .A4(new_n542), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1113), .A2(new_n1105), .A3(new_n1115), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1104), .A2(new_n1118), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1066), .A2(new_n1112), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1107), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1956), .B1(new_n1133), .B2(new_n1070), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT117), .B(new_n1114), .C1(new_n1131), .C2(new_n1134), .ZN(new_n1135));
  OR3_X1    g710(.A1(new_n1095), .A2(KEYINPUT116), .A3(new_n842), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT116), .B1(new_n1095), .B2(new_n842), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1129), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1117), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1127), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1088), .A2(G8), .A3(new_n1077), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT109), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1088), .A2(KEYINPUT109), .A3(G8), .A4(new_n1077), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1077), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1079), .B(new_n1070), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n1087), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT115), .B(new_n1146), .C1(new_n1148), .C2(new_n1039), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1039), .B1(new_n1147), .B2(new_n1087), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1077), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1073), .B(G168), .C1(new_n1066), .C2(G1966), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(G8), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(G8), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1155), .A2(new_n1162), .A3(G8), .A4(new_n1156), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1158), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1074), .A2(G286), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1084), .A2(new_n749), .A3(new_n1005), .A4(new_n1085), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT53), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(KEYINPUT121), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(KEYINPUT121), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1167), .A2(KEYINPUT122), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1093), .A2(new_n683), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(G301), .B(KEYINPUT54), .ZN(new_n1177));
  NOR4_X1   g752(.A1(new_n1003), .A2(new_n1065), .A3(new_n1168), .A4(G2078), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1004), .B(KEYINPUT123), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1066), .A2(KEYINPUT53), .A3(new_n749), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1173), .A2(new_n1181), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1176), .A2(new_n1180), .B1(new_n1182), .B2(new_n1177), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1140), .A2(new_n1154), .A3(new_n1166), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1166), .A2(KEYINPUT62), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1182), .A2(G171), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1145), .A2(new_n1153), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1164), .A2(new_n1188), .A3(new_n1165), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1075), .A2(KEYINPUT63), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1191), .A2(new_n1153), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1184), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1063), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1091), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(G290), .A2(G1986), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1006), .B1(new_n1023), .B2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1019), .A2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT107), .Z(new_n1199));
  OAI21_X1  g774(.A(new_n1036), .B1(new_n1195), .B2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(G319), .ZN(new_n1202));
  OR2_X1    g776(.A1(G227), .A2(new_n1202), .ZN(new_n1203));
  OR2_X1    g777(.A1(new_n1203), .A2(KEYINPUT126), .ZN(new_n1204));
  OAI211_X1 g778(.A(new_n679), .B(new_n1204), .C1(new_n990), .C2(new_n992), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1203), .A2(KEYINPUT126), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n894), .A2(new_n641), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n641), .ZN(new_n1209));
  AND3_X1   g783(.A1(new_n887), .A2(G160), .A3(new_n889), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1210), .A2(new_n890), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1209), .B1(new_n1211), .B2(new_n892), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n988), .B1(new_n978), .B2(new_n980), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n1213), .A2(KEYINPUT103), .ZN(new_n1214));
  AND2_X1   g788(.A1(new_n989), .A2(KEYINPUT103), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n1214), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g790(.A1(new_n1212), .A2(new_n1216), .A3(new_n679), .A4(new_n1204), .ZN(G225));
endmodule


