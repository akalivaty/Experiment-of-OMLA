//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1105, new_n1106,
    new_n1107, new_n1108;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  XOR2_X1   g013(.A(KEYINPUT68), .B(G96), .Z(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XOR2_X1   g016(.A(KEYINPUT69), .B(G57), .Z(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT70), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n463), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n464), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n468), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n468), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n478), .B2(G2105), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n464), .A2(new_n468), .A3(new_n466), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G124), .A3(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT73), .ZN(new_n485));
  INV_X1    g060(.A(new_n469), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n482), .B(new_n485), .C1(G136), .C2(new_n486), .ZN(G162));
  NOR2_X1   g062(.A1(new_n467), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT74), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT74), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(new_n468), .A3(new_n464), .A4(new_n466), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n466), .A3(G2105), .A4(new_n468), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n496), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n465), .A2(G2104), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT71), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n468), .A2(new_n472), .A3(new_n473), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n467), .A2(G138), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT4), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n501), .A2(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(G88), .A2(new_n514), .B1(new_n516), .B2(G50), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT76), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI221_X1 g105(.A(new_n528), .B1(new_n515), .B2(new_n529), .C1(new_n530), .C2(new_n513), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(G90), .A2(new_n514), .B1(new_n516), .B2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n518), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n533), .B1(new_n536), .B2(KEYINPUT77), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(KEYINPUT77), .B2(new_n536), .ZN(G171));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n513), .A2(new_n539), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n518), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT78), .Z(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n516), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(new_n512), .ZN(new_n554));
  XOR2_X1   g129(.A(KEYINPUT79), .B(G65), .Z(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(new_n514), .B2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n552), .A2(new_n557), .ZN(G299));
  XNOR2_X1  g133(.A(G171), .B(KEYINPUT80), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n514), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n516), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G288));
  INV_X1    g142(.A(G86), .ZN(new_n568));
  INV_X1    g143(.A(G48), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n513), .A2(new_n568), .B1(new_n515), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n518), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n513), .A2(new_n575), .B1(new_n515), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n518), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(new_n514), .A2(G92), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT10), .Z(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n554), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n516), .B2(G54), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(G868), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n559), .B2(G868), .ZN(G284));
  AOI21_X1  g165(.A(new_n589), .B1(new_n559), .B2(G868), .ZN(G321));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(G299), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(G168), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(new_n592), .B2(G168), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n583), .B(new_n587), .C1(new_n596), .C2(G860), .ZN(G148));
  INV_X1    g172(.A(new_n544), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n592), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n588), .A2(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n592), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g177(.A(KEYINPUT81), .B1(new_n467), .B2(G111), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n603), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n604));
  NOR3_X1   g179(.A1(new_n467), .A2(KEYINPUT81), .A3(G111), .ZN(new_n605));
  INV_X1    g180(.A(G123), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n604), .A2(new_n605), .B1(new_n500), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G135), .B2(new_n486), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2096), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n506), .A2(new_n461), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT13), .Z(new_n612));
  OAI21_X1  g187(.A(new_n609), .B1(new_n612), .B2(G2100), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G2100), .B2(new_n612), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT82), .Z(G156));
  XOR2_X1   g190(.A(G2427), .B(G2430), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT83), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2438), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT14), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT84), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n619), .B2(new_n617), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT85), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(new_n632), .A3(G14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT86), .ZN(G401));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2100), .Z(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n638), .B2(KEYINPUT18), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(G227));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1956), .B(G2474), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n648), .B1(KEYINPUT87), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(KEYINPUT87), .B2(new_n653), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT20), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n650), .A2(new_n652), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n653), .A3(new_n648), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n659), .C1(new_n648), .C2(new_n658), .ZN(new_n660));
  XOR2_X1   g235(.A(G1991), .B(G1996), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1981), .B(G1986), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(G229));
  INV_X1    g242(.A(G16), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(KEYINPUT90), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(KEYINPUT90), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G22), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(G166), .B2(new_n672), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(G1971), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(G1971), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT32), .B(G1981), .ZN(new_n677));
  NOR2_X1   g252(.A1(G6), .A2(G16), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n573), .B2(G16), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT92), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n675), .B(new_n676), .C1(new_n677), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n677), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n668), .A2(G23), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n566), .B2(new_n668), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT93), .Z(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  INV_X1    g268(.A(G119), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n467), .A2(G107), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n696));
  OAI22_X1  g271(.A1(new_n500), .A2(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G131), .B2(new_n486), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n693), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT89), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n671), .A2(G24), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n580), .B2(new_n671), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT91), .B(G1986), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n700), .A2(new_n701), .ZN(new_n707));
  NOR4_X1   g282(.A1(new_n691), .A2(new_n702), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n690), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n690), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G168), .A2(new_n668), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n668), .B2(G21), .ZN(new_n715));
  INV_X1    g290(.A(G1966), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n668), .A2(G4), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n588), .B2(G16), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n720), .B2(G1348), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G1348), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n692), .A2(G27), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT99), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G164), .B2(new_n692), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G2078), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n672), .A2(G20), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT23), .Z(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G299), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1956), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G2078), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n672), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n544), .B2(new_n672), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G28), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n692), .B1(new_n736), .B2(G28), .ZN(new_n738));
  AND2_X1   g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NOR2_X1   g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n608), .B2(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n668), .A2(G5), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G171), .B2(new_n668), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n735), .B(new_n742), .C1(new_n744), .C2(G1961), .ZN(new_n745));
  NOR4_X1   g320(.A1(new_n722), .A2(new_n726), .A3(new_n732), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n692), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n692), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT29), .B(G2090), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n748), .B(new_n749), .Z(new_n750));
  AOI21_X1  g325(.A(KEYINPUT98), .B1(new_n744), .B2(G1961), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n744), .A2(KEYINPUT98), .A3(G1961), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n746), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n692), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n486), .A2(G139), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n506), .A2(G127), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n467), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n756), .B(new_n757), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n754), .B1(new_n764), .B2(new_n692), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  NOR2_X1   g341(.A1(G29), .A2(G32), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n461), .A2(G105), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT95), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n486), .A2(G141), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n483), .A2(G129), .A3(G2105), .ZN(new_n773));
  AND4_X1   g348(.A1(new_n768), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT96), .Z(new_n775));
  AOI21_X1  g350(.A(new_n767), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT27), .B(G1996), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n715), .A2(new_n716), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  AND2_X1   g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n692), .B1(KEYINPUT24), .B2(G34), .ZN(new_n782));
  OAI22_X1  g357(.A1(G160), .A2(new_n692), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n692), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  INV_X1    g362(.A(G128), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n467), .A2(G116), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n500), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G140), .B2(new_n486), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(new_n692), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n780), .A2(new_n785), .A3(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n753), .A2(new_n766), .A3(new_n778), .A4(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n713), .A2(new_n797), .ZN(G311));
  NAND2_X1  g373(.A1(new_n713), .A2(new_n797), .ZN(G150));
  INV_X1    g374(.A(KEYINPUT100), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n544), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT101), .ZN(new_n802));
  AOI22_X1  g377(.A1(G93), .A2(new_n514), .B1(new_n516), .B2(G55), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n518), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n800), .B2(new_n544), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n802), .A2(new_n806), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n588), .A2(new_n596), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n813));
  AOI21_X1  g388(.A(G860), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n805), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(G145));
  INV_X1    g394(.A(new_n764), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(new_n774), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n775), .B2(new_n820), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n483), .A2(new_n497), .B1(new_n490), .B2(new_n495), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n483), .A2(G126), .A3(G2105), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n507), .B1(new_n504), .B2(new_n505), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n823), .B(new_n824), .C1(KEYINPUT4), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n792), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n822), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n698), .B(KEYINPUT103), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n611), .ZN(new_n830));
  INV_X1    g405(.A(G130), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n467), .A2(G118), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n500), .A2(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G142), .B2(new_n486), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n830), .B(new_n835), .Z(new_n836));
  AOI21_X1  g411(.A(KEYINPUT104), .B1(new_n828), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n828), .ZN(new_n838));
  XOR2_X1   g413(.A(G162), .B(G160), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n608), .ZN(new_n840));
  AOI21_X1  g415(.A(G37), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n838), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g418(.A1(new_n805), .A2(new_n592), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n588), .B(G299), .Z(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(KEYINPUT41), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n807), .A2(new_n808), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n600), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n848), .B2(new_n851), .ZN(new_n853));
  XNOR2_X1  g428(.A(G166), .B(G288), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n573), .B(new_n580), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n844), .B1(new_n859), .B2(new_n592), .ZN(G295));
  OAI21_X1  g435(.A(new_n844), .B1(new_n859), .B2(new_n592), .ZN(G331));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n862));
  NOR2_X1   g437(.A1(G171), .A2(G168), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n559), .B2(G168), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n850), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n850), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(new_n864), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n869), .A2(new_n872), .A3(new_n849), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n848), .B1(new_n869), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n856), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n872), .A3(new_n849), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n869), .A2(new_n872), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n856), .B(new_n877), .C1(new_n878), .C2(new_n848), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n862), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n875), .B2(new_n856), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n884));
  INV_X1    g459(.A(new_n856), .ZN(new_n885));
  MUX2_X1   g460(.A(KEYINPUT41), .B(new_n846), .S(new_n845), .Z(new_n886));
  AND3_X1   g461(.A1(new_n869), .A2(new_n872), .A3(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n884), .B(new_n885), .C1(new_n887), .C2(new_n874), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n887), .B2(new_n874), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT108), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n882), .B1(new_n891), .B2(new_n862), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT44), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n883), .A2(new_n890), .A3(new_n862), .A4(new_n888), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n876), .B2(new_n881), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(G397));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n900));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n501), .B2(new_n509), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n905));
  INV_X1    g480(.A(new_n471), .ZN(new_n906));
  INV_X1    g481(.A(new_n477), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n506), .B2(G125), .ZN(new_n908));
  OAI211_X1 g483(.A(G40), .B(new_n906), .C1(new_n908), .C2(new_n467), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT110), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(KEYINPUT110), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G1996), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n900), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n915), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n792), .B(G2067), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n920), .A2(new_n774), .ZN(new_n921));
  OAI22_X1  g496(.A1(new_n918), .A2(new_n919), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT47), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n775), .A2(new_n917), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n924), .B(new_n920), .C1(new_n917), .C2(new_n774), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n916), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT112), .Z(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n701), .A3(new_n698), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n792), .A2(new_n794), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n916), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT48), .Z(new_n933));
  XNOR2_X1  g508(.A(new_n698), .B(new_n701), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n916), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n936), .B2(KEYINPUT126), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n923), .B(new_n930), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n911), .A2(new_n905), .ZN(new_n940));
  INV_X1    g515(.A(new_n902), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G8), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1981), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n573), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT115), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(KEYINPUT49), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT49), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n946), .B2(new_n573), .ZN(new_n952));
  OAI211_X1 g527(.A(G1981), .B(G305), .C1(new_n950), .C2(new_n949), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n945), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1976), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n954), .A2(new_n955), .A3(new_n566), .ZN(new_n956));
  INV_X1    g531(.A(new_n947), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n945), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G303), .A2(G8), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT55), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n962), .B(new_n901), .C1(new_n501), .C2(new_n509), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR4_X1   g541(.A1(new_n965), .A2(new_n910), .A3(new_n966), .A4(new_n471), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n961), .B(new_n963), .C1(new_n964), .C2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G2090), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n940), .A2(new_n971), .A3(new_n904), .ZN(new_n972));
  INV_X1    g547(.A(G1971), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n969), .A2(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n960), .A2(G8), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n566), .A2(G1976), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT114), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n945), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT52), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n955), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n945), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n984), .A3(new_n954), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n958), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n985), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n959), .B(KEYINPUT55), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n944), .B2(new_n974), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n969), .A2(new_n784), .B1(new_n972), .B2(new_n716), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n990), .A2(new_n944), .A3(G286), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n978), .A2(new_n987), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT63), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n977), .A2(G8), .A3(new_n976), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n988), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n991), .A2(KEYINPUT63), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n978), .A3(new_n987), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n986), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n944), .B1(new_n990), .B2(G168), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G168), .B2(new_n990), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT51), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT125), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n978), .A2(new_n987), .A3(new_n989), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n969), .A2(G1961), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n972), .A2(G2078), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(KEYINPUT123), .A2(KEYINPUT53), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(KEYINPUT123), .A3(KEYINPUT53), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n559), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1011), .B(new_n1020), .C1(KEYINPUT62), .C2(new_n1005), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n999), .B1(new_n1010), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n971), .A2(new_n904), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n909), .A2(new_n1025), .A3(G2078), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1012), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(KEYINPUT53), .B2(new_n1013), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1023), .B1(new_n1028), .B2(G171), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1016), .A2(G301), .A3(new_n1017), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1029), .A2(new_n1030), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1027), .B(G301), .C1(KEYINPUT53), .C2(new_n1013), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1019), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT124), .B1(new_n1033), .B2(new_n1023), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT124), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1035), .B(KEYINPUT54), .C1(new_n1019), .C2(new_n1032), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1031), .B(new_n1011), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT57), .B1(new_n557), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(G299), .B(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT116), .B(G1956), .Z(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n968), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT117), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n968), .A2(new_n1046), .A3(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT56), .B(G2072), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1024), .A2(new_n940), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1041), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n963), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n962), .B1(new_n826), .B2(new_n901), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(KEYINPUT117), .B(new_n1042), .C1(new_n1054), .C2(new_n940), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1046), .B1(new_n968), .B2(new_n1043), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1041), .B(new_n1050), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1038), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT58), .B(G1341), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n943), .A2(new_n1060), .B1(new_n972), .B2(G1996), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n544), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT59), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(new_n544), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1041), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1068), .A2(KEYINPUT120), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT120), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1057), .A2(KEYINPUT61), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT121), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1068), .A2(KEYINPUT120), .A3(new_n1069), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(KEYINPUT61), .A3(new_n1078), .A4(new_n1057), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1059), .A4(new_n1066), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n969), .A2(G1348), .B1(G2067), .B2(new_n942), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT119), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  OAI221_X1 g659(.A(new_n1084), .B1(new_n942), .B2(G2067), .C1(new_n969), .C2(G1348), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n588), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n588), .B1(new_n1086), .B2(KEYINPUT60), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1087), .A2(new_n1088), .B1(KEYINPUT60), .B2(new_n1086), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1074), .A2(new_n1081), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1086), .A2(new_n588), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1057), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1037), .B1(new_n1094), .B2(KEYINPUT122), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1090), .A2(new_n1096), .A3(new_n1093), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1022), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G290), .A2(G1986), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n927), .B(new_n935), .C1(new_n915), .C2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n939), .B1(new_n1098), .B2(new_n1102), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g678(.A(G227), .ZN(new_n1105));
  NAND2_X1  g679(.A1(new_n1105), .A2(G319), .ZN(new_n1106));
  XOR2_X1   g680(.A(new_n1106), .B(KEYINPUT127), .Z(new_n1107));
  NOR3_X1   g681(.A1(G401), .A2(G229), .A3(new_n1107), .ZN(new_n1108));
  AND3_X1   g682(.A1(new_n1108), .A2(new_n842), .A3(new_n896), .ZN(G308));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n842), .A3(new_n896), .ZN(G225));
endmodule


