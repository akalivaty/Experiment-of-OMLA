//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT69), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G113gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(KEYINPUT70), .B2(new_n206), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT70), .B2(new_n206), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(new_n204), .A3(new_n202), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT80), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT2), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n216), .A2(new_n219), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n220), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n224), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n215), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n214), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n223), .A2(new_n236), .A3(new_n231), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n237), .A3(new_n214), .ZN(new_n238));
  NAND2_X1  g037(.A1(G225gat), .A2(G233gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n214), .B2(new_n232), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n234), .A2(new_n238), .A3(new_n239), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n214), .A2(new_n232), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n233), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT5), .B1(new_n246), .B2(new_n239), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n242), .ZN(new_n248));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT0), .ZN(new_n250));
  XNOR2_X1  g049(.A(G57gat), .B(G85gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n244), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n244), .B2(new_n248), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT81), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n254), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT6), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n248), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n252), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT81), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n255), .A4(new_n254), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n258), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT22), .ZN(new_n267));
  INV_X1    g066(.A(G211gat), .ZN(new_n268));
  INV_X1    g067(.A(G218gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G211gat), .B(G218gat), .Z(new_n272));
  OR2_X1    g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n272), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT74), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(KEYINPUT74), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n278));
  MUX2_X1   g077(.A(G183gat), .B(new_n278), .S(G190gat), .Z(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n279), .A2(new_n282), .B1(KEYINPUT64), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(KEYINPUT23), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(KEYINPUT23), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(new_n288), .B2(KEYINPUT64), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n280), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n279), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n288), .A2(new_n294), .A3(KEYINPUT25), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n288), .A2(new_n294), .A3(KEYINPUT66), .A4(KEYINPUT25), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n291), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n303), .B2(KEYINPUT26), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n283), .A2(KEYINPUT67), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n286), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(KEYINPUT26), .B2(new_n303), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n307), .A2(new_n309), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n310), .A2(KEYINPUT68), .A3(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n321), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n299), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n277), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n326), .A2(new_n299), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n320), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n321), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n327), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT29), .B1(new_n326), .B2(new_n299), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT75), .B1(new_n339), .B2(new_n327), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n329), .B(new_n333), .C1(new_n341), .C2(new_n277), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT30), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n341), .A2(new_n277), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n333), .B1(new_n345), .B2(new_n329), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n329), .B1(new_n341), .B2(new_n277), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n332), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n265), .A2(new_n344), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT31), .B(G50gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g153(.A(G228gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n237), .A2(new_n320), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n277), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n273), .B2(new_n274), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n232), .B1(new_n360), .B2(KEYINPUT3), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n357), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n358), .B2(new_n277), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n236), .B1(new_n277), .B2(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n232), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT83), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n354), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(G22gat), .B1(new_n371), .B2(KEYINPUT84), .ZN(new_n375));
  INV_X1    g174(.A(new_n362), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n364), .A2(new_n369), .A3(new_n366), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n369), .B1(new_n364), .B2(new_n366), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT85), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT85), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n371), .A2(KEYINPUT84), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n374), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n379), .B(new_n372), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n354), .B(KEYINPUT82), .Z(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n351), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT34), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n210), .A2(new_n213), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n334), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n326), .A2(new_n214), .A3(new_n299), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G227gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n356), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n393), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AOI211_X1 g200(.A(KEYINPUT34), .B(new_n399), .C1(new_n395), .C2(new_n396), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n399), .A3(new_n396), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n404), .B(KEYINPUT32), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n404), .B2(new_n405), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n404), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT71), .B1(new_n404), .B2(KEYINPUT32), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n403), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n416));
  INV_X1    g215(.A(new_n403), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n413), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n411), .A3(new_n410), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT73), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n403), .A4(new_n409), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT36), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(KEYINPUT72), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n403), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n416), .A2(KEYINPUT72), .A3(new_n417), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT36), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n332), .B1(new_n347), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n341), .A2(new_n276), .A3(new_n275), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n322), .A2(new_n328), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n436), .B2(new_n277), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n434), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n262), .A2(new_n255), .A3(new_n254), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n260), .A4(new_n348), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n347), .A2(new_n431), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n333), .A2(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n346), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT87), .B1(new_n444), .B2(new_n433), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n432), .B1(new_n431), .B2(new_n347), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n434), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n239), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n234), .A2(new_n241), .ZN(new_n451));
  INV_X1    g250(.A(new_n238), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n246), .B2(new_n239), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n252), .C1(KEYINPUT39), .C2(new_n453), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT40), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n459), .A2(new_n460), .A3(new_n259), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n344), .A2(new_n350), .A3(new_n346), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n375), .A2(new_n381), .A3(KEYINPUT85), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n373), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n390), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n392), .B(new_n430), .C1(new_n449), .C2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n427), .B(new_n428), .C1(new_n387), .C2(new_n390), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n471), .B2(new_n351), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n440), .A2(new_n260), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n423), .A2(KEYINPUT35), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n462), .B1(new_n467), .B2(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT88), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n470), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(KEYINPUT91), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  AOI21_X1  g285(.A(G1gat), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n482), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n485), .B2(new_n488), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G29gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT14), .ZN(new_n500));
  OR2_X1    g299(.A1(G43gat), .A2(G50gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  NAND2_X1  g301(.A1(G43gat), .A2(G50gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n495), .A2(new_n497), .A3(new_n500), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n498), .B1(new_n492), .B2(new_n493), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n497), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n501), .B(new_n503), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n504), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n509), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n491), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT92), .Z(new_n518));
  NOR2_X1   g317(.A1(new_n489), .A2(new_n490), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n513), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n516), .A2(KEYINPUT18), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n519), .B(new_n520), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n518), .B(KEYINPUT13), .Z(new_n526));
  AOI22_X1  g325(.A1(new_n522), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT12), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n530), .B2(KEYINPUT94), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n528), .A2(new_n539), .A3(new_n529), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n538), .A2(new_n524), .A3(new_n527), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n479), .A2(new_n481), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G57gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G64gat), .ZN(new_n551));
  INV_X1    g350(.A(G64gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n548), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G127gat), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n549), .A2(new_n557), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n519), .B1(KEYINPUT21), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n217), .ZN(new_n568));
  XOR2_X1   g367(.A(G183gat), .B(G211gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT8), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(KEYINPUT95), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n582), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT96), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND4_X1   g391(.A1(KEYINPUT95), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT95), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n590), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n591), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n592), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n514), .B2(new_n515), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n520), .A2(new_n602), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n604), .A2(new_n605), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n579), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(new_n578), .A3(new_n606), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n591), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n589), .A2(KEYINPUT97), .A3(new_n590), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n564), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n558), .A2(new_n592), .A3(new_n599), .A4(new_n598), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G230gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n356), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT10), .B1(new_n617), .B2(new_n618), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n600), .A2(new_n627), .A3(new_n558), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n622), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  INV_X1    g433(.A(new_n629), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n635), .B2(new_n623), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n574), .A2(new_n613), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n543), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n265), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(G1gat), .Z(G1324gat));
  INV_X1    g443(.A(new_n462), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n482), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n648), .B2(new_n650), .ZN(G1325gat));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n425), .B2(new_n429), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n425), .A2(new_n653), .A3(new_n429), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n642), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n423), .A2(G15gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n642), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n642), .A2(new_n468), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT101), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR3_X1   g463(.A1(new_n640), .A2(new_n573), .A3(new_n612), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n543), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n265), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n498), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT45), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n425), .A2(new_n653), .A3(new_n429), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n654), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n392), .B1(new_n449), .B2(new_n469), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n477), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n613), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n612), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n479), .A2(new_n481), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n640), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n680), .A2(new_n542), .A3(new_n574), .A4(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G29gat), .B1(new_n682), .B2(new_n265), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n670), .A2(new_n683), .ZN(G1328gat));
  NOR3_X1   g483(.A1(new_n666), .A2(new_n645), .A3(new_n494), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n494), .B1(new_n682), .B2(new_n645), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1329gat));
  OAI21_X1  g487(.A(G43gat), .B1(new_n682), .B2(new_n657), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n423), .A2(G43gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n666), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1330gat));
  NOR3_X1   g492(.A1(new_n666), .A2(G50gat), .A3(new_n468), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(KEYINPUT102), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G50gat), .B1(new_n682), .B2(new_n468), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1331gat));
  INV_X1    g499(.A(new_n542), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n681), .A2(new_n574), .A3(new_n613), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n674), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n265), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(new_n550), .ZN(G1332gat));
  XNOR2_X1  g504(.A(new_n703), .B(KEYINPUT103), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n462), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT49), .B(G64gat), .Z(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT104), .ZN(G1333gat));
  NAND3_X1  g510(.A1(new_n706), .A2(G71gat), .A3(new_n672), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n703), .A2(new_n423), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(G71gat), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n391), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT106), .B(G78gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1335gat));
  NOR3_X1   g518(.A1(new_n681), .A2(new_n573), .A3(new_n542), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n680), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n265), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n573), .A2(new_n542), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n674), .A2(new_n613), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n674), .A2(KEYINPUT51), .A3(new_n613), .A4(new_n724), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT107), .B1(new_n725), .B2(new_n726), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n668), .A2(new_n585), .A3(new_n640), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n722), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  NAND4_X1  g532(.A1(new_n677), .A2(new_n679), .A3(new_n462), .A4(new_n720), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n734), .A2(G92gat), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n645), .A2(G92gat), .A3(new_n681), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT108), .Z(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n727), .B2(new_n728), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT52), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n729), .B2(new_n730), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT52), .B1(new_n734), .B2(G92gat), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(KEYINPUT110), .B(new_n739), .C1(new_n743), .C2(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n721), .B2(new_n657), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n423), .A2(G99gat), .A3(new_n681), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n731), .B2(new_n751), .ZN(G1338gat));
  NAND3_X1  g551(.A1(new_n680), .A2(new_n391), .A3(new_n720), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n468), .A2(G106gat), .A3(new_n681), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n731), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n727), .B2(new_n728), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n753), .B2(G106gat), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n756), .A2(new_n759), .B1(new_n761), .B2(new_n755), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n619), .A2(new_n627), .ZN(new_n763));
  INV_X1    g562(.A(new_n628), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n764), .A3(new_n621), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT111), .A4(new_n621), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(KEYINPUT54), .A3(new_n629), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n770), .B(new_n622), .C1(new_n626), .C2(new_n628), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(new_n634), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(KEYINPUT55), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n612), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n771), .A2(KEYINPUT55), .A3(new_n634), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n768), .A2(KEYINPUT54), .A3(new_n629), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n626), .A2(new_n628), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT111), .B1(new_n777), .B2(new_n621), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n769), .A2(KEYINPUT112), .A3(new_n775), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n783), .B2(new_n633), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n625), .A2(new_n629), .A3(new_n632), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n785), .B(new_n786), .C1(new_n781), .C2(new_n782), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n774), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n525), .A2(new_n526), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n518), .B1(new_n516), .B2(new_n521), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n535), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n541), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n530), .A2(KEYINPUT94), .ZN(new_n795));
  INV_X1    g594(.A(new_n536), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n540), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n524), .A2(new_n527), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT114), .B(new_n791), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n788), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n782), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT112), .B1(new_n769), .B2(new_n775), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n633), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n785), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n786), .B1(new_n781), .B2(new_n782), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n799), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT114), .B1(new_n541), .B2(new_n791), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n808), .A2(new_n811), .A3(new_n812), .A4(new_n774), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n801), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n640), .A2(new_n541), .A3(new_n791), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n784), .A2(new_n787), .ZN(new_n816));
  INV_X1    g615(.A(new_n773), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n542), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n612), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n573), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n641), .A2(new_n701), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT116), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n801), .A2(new_n813), .B1(new_n819), .B2(new_n612), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n825), .B(new_n822), .C1(new_n826), .C2(new_n573), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n645), .A2(new_n668), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n423), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n468), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n205), .A3(new_n701), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n427), .A2(new_n428), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n828), .A2(new_n668), .A3(new_n833), .A4(new_n475), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n834), .A2(new_n701), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n835), .B2(new_n205), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n831), .B2(new_n681), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n640), .A2(new_n207), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT117), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n834), .B2(new_n839), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n831), .B2(new_n574), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n574), .A2(G127gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n834), .B2(new_n842), .ZN(G1342gat));
  NOR3_X1   g642(.A1(new_n834), .A2(G134gat), .A3(new_n612), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n831), .B2(new_n612), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n847), .B(new_n848), .C1(new_n845), .C2(new_n844), .ZN(G1343gat));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n824), .A2(new_n391), .A3(new_n827), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(KEYINPUT119), .A3(new_n852), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n773), .B(KEYINPUT120), .Z(new_n857));
  NAND2_X1  g656(.A1(new_n542), .A2(new_n806), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n815), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n612), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n814), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n574), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n852), .B(new_n468), .C1(new_n862), .C2(new_n822), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n855), .A2(new_n856), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n672), .A2(new_n829), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n542), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n672), .A2(new_n468), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n645), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n828), .A3(new_n668), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n701), .A2(G141gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(KEYINPUT121), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(new_n874), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n850), .B1(new_n868), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT58), .B1(new_n873), .B2(new_n874), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(new_n867), .B2(G141gat), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n881), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n875), .A2(new_n878), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n867), .B2(G141gat), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n885), .B(new_n886), .C1(new_n888), .C2(new_n850), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n884), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(G148gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n891), .A3(new_n640), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n865), .A2(new_n866), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n891), .C1(new_n893), .C2(new_n640), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n896));
  INV_X1    g695(.A(new_n788), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n800), .B1(new_n897), .B2(KEYINPUT123), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(KEYINPUT123), .B2(new_n897), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n573), .B1(new_n899), .B2(new_n860), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n852), .B(new_n391), .C1(new_n900), .C2(new_n823), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n681), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n866), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n895), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n892), .B1(new_n894), .B2(new_n905), .ZN(G1345gat));
  AOI21_X1  g705(.A(G155gat), .B1(new_n873), .B2(new_n573), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n573), .A2(G155gat), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT124), .Z(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n893), .B2(new_n909), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n873), .B2(new_n613), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n612), .A2(new_n218), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n893), .B2(new_n912), .ZN(G1347gat));
  NAND2_X1  g712(.A1(new_n462), .A2(new_n265), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n423), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n828), .A2(new_n468), .A3(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(new_n301), .A3(new_n701), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n828), .A2(new_n265), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n645), .A3(new_n471), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n542), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(new_n301), .ZN(G1348gat));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n302), .A3(new_n640), .ZN(new_n922));
  OAI21_X1  g721(.A(G176gat), .B1(new_n916), .B2(new_n681), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1349gat));
  NOR2_X1   g723(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n311), .A3(new_n573), .ZN(new_n926));
  OAI21_X1  g725(.A(G183gat), .B1(new_n916), .B2(new_n574), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n928), .B(new_n929), .Z(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n916), .B2(new_n612), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n919), .A2(new_n312), .A3(new_n613), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT126), .ZN(G1351gat));
  INV_X1    g734(.A(new_n902), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n672), .A2(new_n914), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(new_n701), .ZN(new_n940));
  INV_X1    g739(.A(new_n918), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n869), .A2(new_n462), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n542), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n940), .A2(new_n946), .ZN(G1352gat));
  NOR3_X1   g746(.A1(new_n944), .A2(G204gat), .A3(new_n681), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n903), .A2(new_n937), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G204gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n573), .A3(new_n937), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n268), .B1(KEYINPUT127), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT63), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n953), .B(new_n955), .C1(KEYINPUT127), .C2(new_n954), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n945), .A2(new_n268), .A3(new_n573), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n938), .B2(new_n612), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n269), .A3(new_n613), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


