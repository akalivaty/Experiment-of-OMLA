//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n189), .B2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n195), .A2(new_n196), .B1(G143), .B2(new_n189), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n187), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n203), .B1(new_n209), .B2(G137), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n214), .A2(new_n207), .A3(new_n206), .A4(new_n210), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(new_n205), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n190), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n190), .A2(new_n192), .A3(new_n220), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n190), .A2(new_n192), .A3(new_n220), .A4(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n213), .B1(new_n216), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT2), .B(G113), .Z(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n233), .B(new_n234), .Z(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n215), .A2(G131), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n208), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n228), .A3(new_n223), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT30), .A3(new_n213), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n213), .B(new_n235), .C1(new_n216), .C2(new_n229), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G101), .ZN(new_n244));
  NOR2_X1   g058(.A1(G237), .A2(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G210), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n244), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n242), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n235), .B1(new_n239), .B2(new_n213), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT28), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT69), .B1(new_n242), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n249), .B(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n242), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n230), .A2(new_n236), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT71), .A3(new_n242), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n242), .A2(KEYINPUT71), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(KEYINPUT28), .A3(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n242), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(new_n249), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT29), .A4(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n250), .A2(new_n259), .A3(KEYINPUT70), .A4(new_n260), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n263), .A2(new_n264), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G472), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n241), .A2(new_n242), .A3(new_n271), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n241), .A2(KEYINPUT31), .A3(new_n242), .A4(new_n271), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n280));
  INV_X1    g094(.A(new_n257), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NOR4_X1   g097(.A1(new_n282), .A2(new_n283), .A3(G472), .A4(G902), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n279), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n264), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n283), .B1(new_n289), .B2(G472), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n275), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT16), .ZN(new_n292));
  OR2_X1    g106(.A1(KEYINPUT73), .A2(G125), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT73), .A2(G125), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(G140), .A3(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(G125), .A2(G140), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n294), .ZN(new_n298));
  OR2_X1    g112(.A1(KEYINPUT16), .A2(G140), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G146), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n187), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT24), .B(G110), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n304), .B2(G128), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n308), .B1(new_n312), .B2(G110), .ZN(new_n313));
  XNOR2_X1  g127(.A(G125), .B(G140), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n302), .B(new_n313), .C1(G146), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(G110), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(KEYINPUT72), .A3(G110), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n306), .A2(new_n307), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n295), .A2(new_n296), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(new_n300), .ZN(new_n325));
  AOI21_X1  g139(.A(G146), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n297), .A2(new_n189), .A3(new_n300), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n321), .B(new_n322), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n316), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT22), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(G137), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n329), .B1(new_n316), .B2(new_n328), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n330), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n337), .B1(new_n340), .B2(new_n334), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT25), .A3(new_n264), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  INV_X1    g157(.A(new_n330), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n334), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n336), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n343), .B1(new_n346), .B2(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n264), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G902), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n348), .A2(new_n350), .B1(new_n341), .B2(new_n351), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT75), .B1(new_n291), .B2(new_n352), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n304), .A2(G116), .ZN(new_n356));
  INV_X1    g170(.A(G116), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G119), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT5), .ZN(new_n359));
  OR3_X1    g173(.A1(new_n357), .A2(KEYINPUT5), .A3(G119), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G113), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n233), .A2(new_n234), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G104), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n366), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G107), .ZN(new_n374));
  OAI211_X1 g188(.A(G104), .B(new_n365), .C1(new_n367), .C2(KEYINPUT76), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n371), .A2(new_n372), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n366), .A2(new_n374), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G101), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n377), .B1(new_n376), .B2(new_n379), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n364), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n385));
  INV_X1    g199(.A(new_n366), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n374), .B(new_n375), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(G101), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n376), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n236), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(KEYINPUT83), .B(new_n364), .C1(new_n380), .C2(new_n381), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(G110), .B(G122), .Z(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n395), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n384), .A2(new_n397), .A3(new_n392), .A4(new_n393), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n193), .B(new_n298), .C1(new_n197), .C2(new_n198), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT84), .ZN(new_n401));
  INV_X1    g215(.A(new_n198), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n219), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n193), .A4(new_n298), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n298), .B1(new_n223), .B2(new_n228), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT85), .B(G224), .Z(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G953), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n408), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n394), .A2(new_n414), .A3(new_n395), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n399), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n398), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n395), .B(KEYINPUT8), .Z(new_n420));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n363), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n379), .B1(new_n387), .B2(G101), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT78), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n425), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n364), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n420), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n408), .A2(new_n432), .A3(KEYINPUT7), .A4(new_n412), .ZN(new_n433));
  INV_X1    g247(.A(new_n407), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n401), .A3(new_n405), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n411), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n406), .B2(new_n407), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n431), .A2(new_n433), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n419), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n380), .A2(new_n381), .ZN(new_n443));
  OAI22_X1  g257(.A1(new_n443), .A2(new_n424), .B1(new_n429), .B2(new_n364), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n444), .A2(new_n420), .B1(new_n411), .B2(new_n436), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(KEYINPUT89), .A3(new_n439), .A4(new_n433), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n399), .A2(KEYINPUT86), .A3(new_n413), .A4(new_n415), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n418), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n418), .A2(new_n447), .A3(new_n450), .A4(new_n448), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n454), .A2(new_n453), .ZN(new_n456));
  INV_X1    g270(.A(G221), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT9), .B(G234), .Z(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n264), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n238), .B(KEYINPUT79), .ZN(new_n460));
  OAI211_X1 g274(.A(KEYINPUT10), .B(new_n199), .C1(new_n380), .C2(new_n381), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  INV_X1    g276(.A(new_n193), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT77), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n187), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n190), .A2(KEYINPUT77), .A3(KEYINPUT1), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n190), .A2(new_n192), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n462), .B1(new_n469), .B2(new_n425), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n391), .A2(new_n228), .A3(new_n223), .A4(new_n389), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n460), .A2(new_n461), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n199), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n426), .A2(new_n473), .A3(new_n427), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT80), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n469), .A2(new_n425), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n426), .A2(new_n477), .A3(new_n473), .A4(new_n427), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n479), .A2(KEYINPUT12), .A3(new_n238), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT12), .B1(new_n479), .B2(new_n238), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G140), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n331), .A2(G227), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n472), .A2(new_n487), .A3(new_n485), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n472), .B2(new_n485), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n461), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n470), .A2(new_n471), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n238), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n482), .A2(new_n486), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G469), .B1(new_n494), .B2(G902), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n472), .A2(new_n485), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n480), .B2(new_n481), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n485), .B1(new_n493), .B2(new_n472), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G469), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n501), .A2(new_n264), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n459), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G214), .B1(G237), .B2(G902), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n455), .A2(new_n456), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n373), .ZN(new_n511));
  MUX2_X1   g325(.A(new_n315), .B(new_n323), .S(KEYINPUT19), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n189), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n245), .A2(G143), .A3(G214), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G143), .B1(new_n245), .B2(G214), .ZN(new_n516));
  OAI21_X1  g330(.A(G131), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n245), .A2(G214), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n191), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n205), .A3(new_n514), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n301), .A2(G146), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n511), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n314), .B2(new_n189), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n323), .B2(new_n189), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT18), .B(G131), .C1(new_n515), .C2(new_n516), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n295), .A2(new_n523), .A3(G146), .A4(new_n296), .ZN(new_n527));
  NAND2_X1  g341(.A1(KEYINPUT18), .A2(G131), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n519), .A2(new_n514), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT92), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n519), .A2(new_n514), .A3(new_n528), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n519), .B2(new_n514), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n527), .A4(new_n525), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n522), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G475), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n517), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n517), .A2(new_n520), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n540), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n326), .A2(new_n327), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n536), .A2(new_n531), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n511), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n538), .B(new_n539), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n509), .B1(new_n547), .B2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n544), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n537), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n550), .A2(new_n511), .B1(new_n537), .B2(new_n522), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n539), .A4(new_n264), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n511), .A2(KEYINPUT93), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n264), .B1(new_n545), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n537), .A2(new_n549), .A3(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(G475), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n548), .A2(new_n552), .A3(new_n556), .A4(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n331), .A2(G952), .ZN(new_n562));
  NAND2_X1  g376(.A1(G234), .A2(G237), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT21), .B(G898), .Z(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(G902), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT13), .B1(new_n187), .B2(G143), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n209), .ZN(new_n572));
  XNOR2_X1  g386(.A(G128), .B(G143), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT95), .B(G122), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n575), .A2(new_n357), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n357), .A2(G122), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n365), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n575), .A2(new_n357), .ZN(new_n579));
  INV_X1    g393(.A(new_n577), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n579), .A2(G107), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n574), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT14), .ZN(new_n583));
  OAI22_X1  g397(.A1(new_n575), .A2(new_n357), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT96), .B1(new_n577), .B2(KEYINPUT14), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n586), .A2(new_n583), .A3(new_n357), .A4(G122), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(G107), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n576), .A2(new_n365), .A3(new_n577), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n573), .B(new_n209), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n458), .A2(G217), .A3(new_n331), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n582), .A2(new_n596), .A3(new_n592), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n264), .ZN(new_n601));
  INV_X1    g415(.A(G478), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n602), .A2(KEYINPUT15), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n601), .B(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n561), .A2(new_n570), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n508), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n355), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NAND2_X1  g424(.A1(new_n452), .A2(new_n454), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n507), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n495), .A2(new_n505), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n286), .B2(new_n287), .ZN(new_n614));
  AND2_X1   g428(.A1(KEYINPUT98), .A2(G472), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n459), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n613), .A2(new_n352), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n602), .A2(new_n264), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n600), .A2(new_n602), .A3(new_n264), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n582), .A2(new_n596), .A3(new_n592), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n596), .B1(new_n582), .B2(new_n592), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT99), .B1(new_n625), .B2(KEYINPUT33), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n627), .B(new_n628), .C1(new_n623), .C2(new_n624), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n600), .B2(KEYINPUT100), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n598), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n626), .A2(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n621), .B(new_n622), .C1(new_n633), .C2(new_n602), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n559), .B2(new_n560), .ZN(new_n635));
  INV_X1    g449(.A(new_n570), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n557), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n636), .A3(new_n605), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n619), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(new_n616), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT25), .B1(new_n341), .B2(new_n264), .ZN(new_n652));
  AND4_X1   g466(.A1(KEYINPUT25), .A2(new_n345), .A3(new_n264), .A4(new_n336), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n350), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n316), .A2(new_n328), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n351), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NOR4_X1   g473(.A1(new_n508), .A2(new_n607), .A3(new_n651), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT37), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G110), .ZN(G12));
  INV_X1    g476(.A(new_n507), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n452), .B2(new_n454), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n654), .A2(new_n658), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n564), .B1(new_n568), .B2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n642), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n604), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n291), .A2(new_n506), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n455), .A2(new_n674), .A3(new_n456), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n674), .B1(new_n455), .B2(new_n456), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n455), .A2(new_n456), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n455), .A2(new_n674), .A3(new_n456), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(KEYINPUT38), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G472), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT32), .B1(new_n614), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n266), .A2(new_n267), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n276), .B1(new_n685), .B2(new_n257), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n683), .B1(new_n686), .B2(new_n264), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n684), .A2(new_n284), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n665), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n561), .A2(new_n605), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n507), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT103), .B1(new_n682), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n694));
  INV_X1    g508(.A(new_n692), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n677), .A2(new_n681), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n667), .B(KEYINPUT39), .Z(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n506), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT40), .Z(new_n700));
  NAND3_X1  g514(.A1(new_n693), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  INV_X1    g516(.A(new_n622), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n632), .B(KEYINPUT33), .C1(new_n625), .C2(new_n631), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n627), .B1(new_n600), .B2(new_n628), .ZN(new_n705));
  INV_X1    g519(.A(new_n629), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n620), .B(new_n703), .C1(new_n707), .C2(G478), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n561), .A2(new_n708), .A3(new_n667), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n666), .A2(new_n670), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND2_X1  g526(.A1(new_n341), .A2(new_n351), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n654), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n684), .A2(new_n284), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(new_n275), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n479), .A2(new_n238), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT12), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n479), .A2(KEYINPUT12), .A3(new_n238), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n499), .B1(new_n721), .B2(new_n497), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n505), .A3(new_n617), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(new_n505), .A3(KEYINPUT104), .A4(new_n617), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n716), .A2(new_n664), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n637), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT105), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT41), .B(G113), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n727), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n612), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(KEYINPUT106), .A3(new_n716), .A4(new_n647), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  INV_X1    g550(.A(new_n647), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND3_X1  g554(.A1(new_n726), .A2(new_n291), .A3(new_n727), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n611), .A2(new_n606), .A3(new_n507), .A4(new_n665), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n304), .ZN(G21));
  NAND3_X1  g558(.A1(new_n664), .A2(new_n726), .A3(new_n727), .ZN(new_n745));
  NOR2_X1   g559(.A1(G472), .A2(G902), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n268), .A2(new_n747), .A3(new_n270), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n268), .B2(new_n270), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n748), .A2(new_n749), .A3(new_n257), .ZN(new_n750));
  INV_X1    g564(.A(new_n286), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n289), .A2(G472), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n268), .A2(new_n270), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n268), .A2(new_n270), .A3(new_n747), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n281), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n286), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n746), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n753), .A2(new_n352), .A3(new_n754), .A4(new_n761), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n745), .A2(new_n570), .A3(new_n690), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(G122), .Z(G24));
  AOI21_X1  g578(.A(new_n760), .B1(new_n759), .B2(new_n746), .ZN(new_n765));
  INV_X1    g579(.A(new_n746), .ZN(new_n766));
  AOI211_X1 g580(.A(KEYINPUT108), .B(new_n766), .C1(new_n758), .C2(new_n286), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(KEYINPUT109), .A3(new_n665), .A4(new_n754), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n753), .A2(new_n665), .A3(new_n761), .A4(new_n754), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n709), .A2(KEYINPUT110), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n635), .A2(new_n775), .A3(new_n667), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n734), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  AOI21_X1  g593(.A(new_n663), .B1(new_n455), .B2(new_n456), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n716), .A3(new_n777), .A4(new_n506), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NAND4_X1  g601(.A1(new_n780), .A2(new_n716), .A3(new_n506), .A4(new_n669), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G134), .ZN(G36));
  NAND2_X1  g603(.A1(new_n490), .A2(new_n493), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n491), .A2(new_n492), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n719), .A2(new_n720), .B1(new_n791), .B2(new_n460), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n792), .B2(new_n485), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n494), .A2(KEYINPUT45), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(G469), .ZN(new_n797));
  NAND2_X1  g611(.A1(G469), .A2(G902), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n798), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n505), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n617), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n697), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT43), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n561), .B2(new_n634), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n708), .A2(KEYINPUT43), .A3(new_n559), .A4(new_n560), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n616), .B(new_n659), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n806), .B1(new_n810), .B2(KEYINPUT44), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n651), .A3(new_n665), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(KEYINPUT112), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n780), .B1(new_n813), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT111), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n780), .C1(new_n813), .C2(new_n814), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n805), .A2(new_n816), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  NAND2_X1  g636(.A1(new_n804), .A2(KEYINPUT47), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n291), .A2(new_n352), .A3(new_n709), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n803), .A2(new_n825), .A3(new_n617), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n780), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NOR3_X1   g642(.A1(new_n714), .A2(new_n663), .A3(new_n459), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT113), .ZN(new_n830));
  INV_X1    g644(.A(new_n561), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n708), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT114), .Z(new_n833));
  NAND2_X1  g647(.A1(new_n723), .A2(new_n505), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT49), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n836), .A2(KEYINPUT115), .B1(KEYINPUT49), .B2(new_n834), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(KEYINPUT115), .B2(new_n836), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n682), .A3(new_n688), .ZN(new_n839));
  INV_X1    g653(.A(new_n780), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n733), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n564), .B1(new_n808), .B2(new_n809), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n716), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT48), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n714), .A2(new_n564), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n841), .A2(new_n635), .A3(new_n688), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n562), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n733), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n780), .A3(new_n688), .A4(new_n847), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n561), .A3(new_n708), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n842), .A2(new_n352), .A3(new_n754), .A4(new_n768), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n733), .B2(new_n507), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n726), .A2(KEYINPUT119), .A3(new_n663), .A4(new_n727), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n682), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n682), .A2(new_n857), .A3(KEYINPUT50), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n852), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n723), .A2(new_n505), .A3(new_n459), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT117), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n823), .B2(new_n826), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n853), .A2(new_n840), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  INV_X1    g683(.A(new_n826), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n825), .B1(new_n803), .B2(new_n617), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n866), .C1(new_n872), .C2(new_n864), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n841), .A2(new_n773), .A3(new_n842), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n862), .A2(new_n868), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n849), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n878));
  INV_X1    g692(.A(new_n852), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n682), .A2(KEYINPUT50), .A3(new_n857), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT50), .B1(new_n682), .B2(new_n857), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n874), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n876), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n823), .A2(new_n826), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n867), .B1(new_n884), .B2(new_n863), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n878), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n882), .A2(KEYINPUT120), .A3(new_n885), .A4(new_n876), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n877), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n728), .A2(new_n637), .B1(new_n741), .B2(new_n742), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n763), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n660), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n635), .B1(new_n605), .B2(new_n831), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n618), .A2(new_n894), .A3(new_n570), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n678), .A2(new_n663), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n355), .A2(new_n608), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n892), .A2(new_n893), .A3(new_n739), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n668), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n659), .A2(new_n605), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n780), .A2(new_n670), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(new_n788), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n781), .A2(new_n782), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n783), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n773), .A2(new_n777), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n780), .A2(new_n506), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n898), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n666), .B(new_n670), .C1(new_n669), .C2(new_n710), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n612), .A2(new_n690), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n506), .A3(new_n667), .A4(new_n689), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n778), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT52), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT52), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n778), .A2(new_n911), .A3(new_n913), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n910), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n915), .A2(new_n910), .A3(new_n917), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n909), .B(KEYINPUT53), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT53), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n901), .A2(new_n788), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n784), .B2(new_n785), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n739), .A2(new_n897), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n660), .A2(new_n763), .A3(new_n891), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n907), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n915), .A2(new_n917), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n890), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n909), .B(new_n921), .C1(new_n918), .C2(new_n919), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT53), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT54), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n842), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n933), .A2(new_n745), .A3(new_n762), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n889), .A2(new_n929), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n839), .B1(new_n935), .B2(new_n936), .ZN(G75));
  NAND4_X1  g751(.A1(new_n930), .A2(G210), .A3(G902), .A4(new_n931), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n399), .A2(new_n415), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n413), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT55), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n938), .B2(new_n939), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n331), .A2(G952), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G51));
  XOR2_X1   g760(.A(new_n798), .B(KEYINPUT57), .Z(new_n947));
  AND3_X1   g761(.A1(new_n930), .A2(KEYINPUT54), .A3(new_n931), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n932), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n501), .B(KEYINPUT121), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n797), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n930), .A2(G902), .A3(new_n952), .A4(new_n931), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n945), .B1(new_n951), .B2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n930), .A2(KEYINPUT58), .A3(G902), .A4(new_n931), .ZN(new_n955));
  INV_X1    g769(.A(new_n551), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n955), .A2(new_n539), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n945), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n955), .B2(new_n539), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  XNOR2_X1  g774(.A(new_n620), .B(KEYINPUT59), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n929), .B2(new_n932), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n707), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n633), .B(new_n962), .C1(new_n948), .C2(new_n932), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(new_n958), .A3(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n930), .A2(new_n931), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n346), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n657), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n945), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n970), .A2(KEYINPUT122), .A3(new_n346), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n973), .A2(new_n975), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n971), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n958), .B1(new_n970), .B2(new_n974), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n567), .B2(new_n410), .ZN(new_n984));
  INV_X1    g798(.A(new_n898), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n940), .B1(G898), .B2(new_n331), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n986), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n232), .A2(new_n240), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n512), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(G900), .B1(new_n992), .B2(G227), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n331), .B(new_n993), .C1(G227), .C2(new_n992), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n821), .A2(new_n827), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n716), .A2(new_n664), .A3(new_n691), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n803), .A2(new_n997), .A3(new_n617), .A4(new_n698), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n778), .A3(new_n911), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n785), .B2(new_n784), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n995), .A2(new_n996), .A3(new_n788), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n821), .A2(new_n788), .A3(new_n827), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT126), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n1005), .B2(new_n992), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n699), .B(new_n840), .C1(KEYINPUT125), .C2(new_n894), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1007), .B(new_n355), .C1(KEYINPUT125), .C2(new_n894), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n995), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n778), .A2(new_n911), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n1010), .B2(KEYINPUT62), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n701), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1011), .B1(new_n701), .B2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1009), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n991), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n994), .B1(new_n1006), .B2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(new_n920), .A2(new_n928), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n249), .B1(new_n241), .B2(new_n242), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  NOR2_X1   g837(.A1(new_n243), .A2(new_n271), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1001), .A2(new_n1004), .A3(new_n985), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n1027), .A2(new_n1023), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1026), .B(new_n958), .C1(new_n1028), .C2(new_n1025), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1009), .B(new_n985), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT127), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1030), .A2(new_n1031), .A3(new_n1023), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1031), .B1(new_n1030), .B2(new_n1023), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1029), .B1(new_n1020), .B2(new_n1034), .ZN(G57));
endmodule


