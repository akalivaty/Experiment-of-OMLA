//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(G134gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n205), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  AND3_X1   g022(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n218), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n223), .A2(new_n218), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n226), .A2(new_n225), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT65), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n218), .C1(new_n223), .C2(new_n227), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n229), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n225), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(G190gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G183gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT27), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT27), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G183gat), .ZN(new_n252));
  AND4_X1   g051(.A1(new_n245), .A2(new_n250), .A3(new_n252), .A4(new_n247), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n244), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n246), .A2(KEYINPUT28), .A3(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n252), .A3(new_n247), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n250), .A2(new_n252), .A3(new_n245), .A4(new_n247), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT67), .A3(new_n244), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n243), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n217), .B1(new_n238), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G227gat), .ZN(new_n265));
  INV_X1    g064(.A(G233gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n243), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n261), .A2(new_n244), .B1(KEYINPUT67), .B2(new_n255), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n270), .B(KEYINPUT28), .C1(new_n259), .C2(new_n260), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n205), .A2(new_n212), .A3(new_n215), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n215), .B1(new_n205), .B2(new_n212), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n229), .A2(new_n235), .A3(new_n237), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n264), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n280), .A3(new_n267), .A4(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n202), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT33), .B1(new_n279), .B2(new_n281), .ZN(new_n283));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT70), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT71), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n282), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n264), .A2(new_n277), .ZN(new_n292));
  INV_X1    g091(.A(new_n267), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(KEYINPUT34), .B(new_n267), .C1(new_n264), .C2(new_n277), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI221_X4 g096(.A(new_n202), .B1(KEYINPUT33), .B2(new_n288), .C1(new_n279), .C2(new_n281), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n290), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n281), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT33), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n289), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n282), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n282), .B1(new_n283), .B2(new_n289), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT36), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT83), .ZN(new_n308));
  XOR2_X1   g107(.A(G197gat), .B(G204gat), .Z(new_n309));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT72), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(KEYINPUT73), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G211gat), .B(G218gat), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n317), .B(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G141gat), .B(G148gat), .Z(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n325), .A3(KEYINPUT2), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  OR3_X1    g126(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n328), .A2(new_n329), .B1(G155gat), .B2(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n322), .B1(new_n333), .B2(KEYINPUT2), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n327), .A2(new_n330), .B1(new_n321), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n320), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(G22gat), .Z(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT3), .B1(new_n320), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(new_n340), .C1(new_n342), .C2(new_n335), .ZN(new_n343));
  INV_X1    g142(.A(new_n340), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n317), .A2(new_n319), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n309), .B(new_n318), .C1(new_n315), .C2(new_n316), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n335), .B1(new_n347), .B2(new_n336), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n320), .A2(new_n337), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G78gat), .B(G106gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT81), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT31), .B(G50gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n308), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n343), .A2(new_n350), .A3(KEYINPUT83), .A4(new_n355), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n351), .B2(new_n356), .ZN(new_n360));
  AOI211_X1 g159(.A(KEYINPUT82), .B(new_n355), .C1(new_n343), .C2(new_n350), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n357), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n297), .B1(new_n290), .B2(new_n298), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT36), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n304), .A2(new_n296), .A3(new_n305), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n307), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT4), .B1(new_n217), .B2(new_n335), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n335), .B(KEYINPUT4), .C1(new_n273), .C2(new_n274), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n327), .A2(new_n330), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n334), .A2(new_n321), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n335), .A2(new_n336), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n275), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n335), .B1(new_n273), .B2(new_n274), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n370), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n372), .A2(new_n378), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n375), .A2(new_n214), .A3(new_n216), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n384), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n378), .A2(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n370), .ZN(new_n391));
  OAI211_X1 g190(.A(KEYINPUT5), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT77), .ZN(new_n396));
  XNOR2_X1  g195(.A(G57gat), .B(G85gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AND4_X1   g198(.A1(KEYINPUT80), .A2(new_n393), .A3(KEYINPUT6), .A4(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n386), .B2(new_n392), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT80), .B1(new_n401), .B2(KEYINPUT6), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n320), .ZN(new_n408));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n238), .A2(new_n263), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n272), .A2(new_n276), .ZN(new_n412));
  INV_X1    g211(.A(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n412), .B2(new_n341), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n409), .B1(new_n272), .B2(new_n276), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n416), .A2(new_n320), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n407), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n399), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n386), .A2(new_n392), .A3(new_n398), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT37), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n415), .B2(new_n418), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n320), .B1(new_n416), .B2(new_n417), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n272), .B2(new_n276), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n414), .B(new_n408), .C1(new_n413), .C2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(KEYINPUT37), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n426), .A3(new_n406), .A4(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n403), .A2(new_n419), .A3(new_n423), .A4(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT37), .B1(new_n427), .B2(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n406), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(KEYINPUT85), .A3(new_n406), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n426), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(KEYINPUT30), .B(new_n407), .C1(new_n415), .C2(new_n418), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n427), .A2(new_n406), .A3(new_n429), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT74), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n406), .B1(new_n427), .B2(new_n429), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(KEYINPUT30), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n419), .A2(KEYINPUT74), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n372), .A2(new_n378), .A3(new_n382), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n384), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n448), .A2(new_n384), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n387), .A2(new_n379), .A3(new_n383), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT39), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n398), .B(new_n450), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n384), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(KEYINPUT39), .A3(new_n452), .ZN(new_n458));
  INV_X1    g257(.A(new_n455), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n398), .A3(new_n450), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n420), .A3(new_n460), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n432), .A2(new_n438), .B1(new_n447), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n363), .A2(new_n362), .A3(new_n365), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n444), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n439), .A2(new_n440), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n420), .B2(new_n421), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n401), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n469), .A2(new_n470), .A3(new_n423), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n464), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n423), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n463), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT35), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n367), .A2(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n362), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n307), .A2(new_n478), .A3(new_n366), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n422), .A2(new_n421), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n420), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n403), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n447), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n477), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490));
  XOR2_X1   g289(.A(new_n490), .B(KEYINPUT13), .Z(new_n491));
  INV_X1    g290(.A(G8gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT16), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(G1gat), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n495), .B2(KEYINPUT90), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(G1gat), .B2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI221_X1 g297(.A(new_n495), .B1(KEYINPUT90), .B2(new_n492), .C1(G1gat), .C2(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT92), .ZN(new_n501));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  INV_X1    g304(.A(G36gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT89), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT15), .B(new_n502), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n509), .A4(new_n503), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT93), .B1(new_n501), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n500), .A2(KEYINPUT92), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n516), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n500), .A2(KEYINPUT92), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(KEYINPUT93), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n491), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n500), .B(KEYINPUT91), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n520), .B(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n490), .A3(new_n522), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G113gat), .B(G141gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT11), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT87), .Z(new_n537));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n526), .A2(new_n541), .A3(new_n532), .A4(new_n533), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n546));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  OR2_X1    g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n556), .A2(new_n557), .B1(new_n553), .B2(new_n551), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n557), .B2(new_n556), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n552), .A2(KEYINPUT94), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n551), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n559), .A2(KEYINPUT96), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT96), .B1(new_n559), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n555), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n548), .B1(new_n567), .B2(KEYINPUT21), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT21), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n569), .A3(new_n547), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(new_n568), .B2(new_n570), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n546), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(new_n546), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G183gat), .B(G211gat), .Z(new_n579));
  AND3_X1   g378(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n575), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n501), .B1(new_n569), .B2(new_n566), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT98), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR3_X1    g383(.A1(new_n580), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n580), .B2(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT99), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n528), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n600), .B(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n520), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n589), .A2(KEYINPUT41), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n605), .A2(KEYINPUT101), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT101), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n603), .B(new_n612), .C1(new_n607), .C2(new_n608), .ZN(new_n613));
  XOR2_X1   g412(.A(G134gat), .B(G162gat), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n611), .B2(new_n613), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n592), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n591), .A3(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n587), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n566), .A2(new_n602), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n604), .B(new_n555), .C1(new_n564), .C2(new_n565), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n632), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n640), .B2(new_n635), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n489), .A2(new_n545), .A3(new_n623), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT103), .Z(new_n643));
  INV_X1    g442(.A(new_n485), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT104), .B(G1gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1324gat));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n643), .A2(new_n467), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT42), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(new_n467), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(G8gat), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n649), .B2(new_n653), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n299), .A2(new_n306), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n643), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n307), .ZN(new_n658));
  INV_X1    g457(.A(new_n366), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n662), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n643), .A2(new_n478), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NAND3_X1  g465(.A1(new_n587), .A2(new_n622), .A3(new_n641), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT105), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n545), .A3(new_n489), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n505), .A3(new_n644), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n462), .A2(new_n362), .A3(new_n307), .A4(new_n366), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n473), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT86), .B1(new_n447), .B2(new_n473), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n363), .A2(new_n362), .A3(new_n365), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n673), .B1(new_n677), .B2(KEYINPUT35), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n486), .B1(new_n479), .B2(new_n480), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n622), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n622), .C1(new_n678), .C2(new_n679), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n587), .A2(new_n545), .A3(new_n641), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n485), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n688), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n669), .A2(G36gat), .A3(new_n447), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n687), .B2(new_n447), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  NAND3_X1  g492(.A1(new_n686), .A2(G43gat), .A3(new_n661), .ZN(new_n694));
  INV_X1    g493(.A(new_n656), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n669), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(G43gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g497(.A1(new_n686), .A2(new_n478), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G50gat), .ZN(new_n700));
  OR3_X1    g499(.A1(new_n669), .A2(G50gat), .A3(new_n362), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT48), .B1(new_n702), .B2(KEYINPUT106), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n704), .B(new_n705), .C1(new_n700), .C2(new_n701), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n703), .A2(new_n706), .ZN(G1331gat));
  INV_X1    g506(.A(new_n545), .ZN(new_n708));
  INV_X1    g507(.A(new_n641), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n489), .A2(new_n708), .A3(new_n623), .A4(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(new_n485), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n710), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  AND2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n714), .A2(new_n447), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n467), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n715), .B2(new_n719), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n714), .B2(new_n660), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n710), .A2(G71gat), .A3(new_n695), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(KEYINPUT50), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n718), .A2(new_n478), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  INV_X1    g528(.A(new_n587), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n545), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n622), .B(new_n731), .C1(new_n678), .C2(new_n679), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n734), .A2(new_n597), .A3(new_n644), .A4(new_n709), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n730), .A2(new_n545), .A3(new_n641), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n682), .A2(new_n683), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n485), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1336gat));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n682), .A2(new_n467), .A3(new_n683), .A4(new_n736), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G92gat), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n641), .A2(new_n447), .A3(G92gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n734), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(KEYINPUT112), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(KEYINPUT112), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n740), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n743), .B(KEYINPUT108), .Z(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n621), .B1(new_n477), .B2(new_n488), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n731), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n732), .A2(new_n733), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n754), .A2(KEYINPUT110), .B1(G92gat), .B2(new_n741), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n756), .B(new_n749), .C1(new_n752), .C2(new_n753), .ZN(new_n757));
  AOI211_X1 g556(.A(new_n748), .B(new_n740), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(KEYINPUT110), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n757), .A3(new_n742), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT111), .B1(new_n760), .B2(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n747), .B1(new_n758), .B2(new_n761), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n695), .A2(G99gat), .A3(new_n641), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n734), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G99gat), .B1(new_n737), .B2(new_n660), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1338gat));
  NOR3_X1   g565(.A1(new_n641), .A2(new_n362), .A3(G106gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n734), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n682), .A2(new_n478), .A3(new_n683), .A4(new_n736), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n767), .B1(new_n752), .B2(new_n753), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n777), .B2(new_n769), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n623), .A2(new_n708), .A3(new_n641), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  INV_X1    g581(.A(new_n525), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n523), .B2(new_n518), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n529), .A2(new_n522), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n784), .A2(new_n491), .B1(new_n490), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n539), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n544), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n782), .B1(new_n709), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n544), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n790), .A2(new_n641), .A3(KEYINPUT116), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n636), .ZN(new_n793));
  INV_X1    g592(.A(new_n639), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n635), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n631), .A2(new_n795), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n629), .A2(new_n630), .A3(new_n625), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n545), .A2(new_n793), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  INV_X1    g603(.A(new_n801), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT54), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n797), .B2(new_n801), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n803), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n621), .B1(new_n792), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n808), .B(KEYINPUT55), .C1(new_n797), .C2(new_n801), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n618), .A3(new_n620), .A4(new_n793), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n790), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n809), .B2(new_n811), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT115), .B1(new_n820), .B2(new_n788), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n781), .B1(new_n822), .B2(new_n587), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n485), .A2(new_n467), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n823), .A2(new_n676), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n545), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n779), .B1(new_n827), .B2(G113gat), .ZN(new_n828));
  AOI211_X1 g627(.A(KEYINPUT117), .B(new_n208), .C1(new_n826), .C2(new_n545), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(G113gat), .B2(new_n827), .ZN(G1340gat));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n709), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n730), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n809), .A2(new_n811), .ZN(new_n835));
  INV_X1    g634(.A(new_n818), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n788), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n817), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n788), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n816), .A2(new_n803), .B1(new_n789), .B2(new_n791), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n621), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n780), .B1(new_n841), .B2(new_n730), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(new_n463), .A3(new_n622), .A4(new_n824), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT68), .B(G134gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n846), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n843), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n847), .B1(new_n848), .B2(new_n851), .ZN(G1343gat));
  INV_X1    g651(.A(G141gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n661), .A2(new_n825), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n823), .B2(new_n362), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n839), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n803), .A2(new_n810), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n709), .A2(new_n788), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n622), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n730), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT57), .B(new_n478), .C1(new_n863), .C2(new_n781), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n855), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n853), .B1(new_n865), .B2(new_n545), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n823), .A2(new_n479), .A3(new_n825), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n853), .A3(new_n545), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT58), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n842), .B2(new_n478), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n478), .A2(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n858), .A2(new_n862), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n587), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n874), .B2(new_n780), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n854), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G141gat), .B1(new_n876), .B2(new_n708), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n870), .A2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n881), .A3(new_n709), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT119), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n881), .C1(new_n865), .C2(new_n709), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n842), .A2(KEYINPUT57), .A3(new_n478), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n816), .B2(new_n818), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n835), .A2(KEYINPUT120), .A3(new_n836), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n790), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n587), .B1(new_n890), .B2(new_n861), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n362), .B1(new_n891), .B2(new_n780), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(KEYINPUT57), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n709), .A3(new_n854), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n894), .B2(G148gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n883), .B1(new_n884), .B2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n876), .B2(new_n587), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n867), .A2(new_n331), .A3(new_n730), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n876), .B2(new_n621), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n867), .A2(new_n332), .A3(new_n622), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n823), .A2(KEYINPUT121), .A3(new_n644), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n842), .B2(new_n485), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n463), .B(new_n467), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n708), .A2(G169gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n903), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT121), .B1(new_n823), .B2(new_n644), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n842), .A2(new_n905), .A3(new_n485), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n447), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(KEYINPUT122), .A3(new_n463), .A4(new_n908), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n644), .A2(new_n447), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n463), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n823), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n842), .A2(KEYINPUT123), .A3(new_n463), .A4(new_n917), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n545), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT124), .B1(new_n921), .B2(G169gat), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n915), .A2(new_n924), .ZN(G1348gat));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n920), .A3(new_n709), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G176gat), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n641), .A2(G176gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n907), .B2(new_n928), .ZN(G1349gat));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n912), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n730), .A2(new_n246), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n930), .A2(new_n463), .A3(new_n467), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n920), .A3(new_n730), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT60), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n933), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n919), .A2(new_n920), .A3(new_n622), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(G190gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n941), .B2(G190gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n622), .A2(new_n247), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n943), .A2(new_n944), .B1(new_n907), .B2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n660), .A2(new_n917), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT125), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n893), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n708), .ZN(new_n951));
  AOI211_X1 g750(.A(new_n479), .B(new_n447), .C1(new_n911), .C2(new_n912), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n708), .A2(G197gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  OAI21_X1  g754(.A(G204gat), .B1(new_n950), .B2(new_n641), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n641), .A2(G204gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT62), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n479), .ZN(new_n959));
  AND4_X1   g758(.A1(KEYINPUT62), .A2(new_n913), .A3(new_n959), .A4(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n312), .A3(new_n730), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n587), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n893), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  NOR2_X1   g766(.A1(new_n621), .A2(new_n311), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT127), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n948), .B1(new_n970), .B2(new_n886), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n971), .B2(KEYINPUT126), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n950), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n952), .A2(new_n622), .ZN(new_n975));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n972), .A2(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1355gat));
endmodule


