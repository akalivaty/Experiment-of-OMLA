

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XNOR2_X1 U325 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U326 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U327 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U328 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n463) );
  INV_X1 U329 ( .A(KEYINPUT73), .ZN(n441) );
  INV_X1 U330 ( .A(G71GAT), .ZN(n373) );
  XNOR2_X1 U331 ( .A(n464), .B(n463), .ZN(n470) );
  XNOR2_X1 U332 ( .A(n374), .B(n373), .ZN(n381) );
  XNOR2_X1 U333 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n471) );
  XNOR2_X1 U334 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n389) );
  XNOR2_X1 U335 ( .A(n472), .B(n471), .ZN(n482) );
  XNOR2_X1 U336 ( .A(n390), .B(n389), .ZN(n574) );
  XOR2_X1 U337 ( .A(n385), .B(n384), .Z(n490) );
  XNOR2_X1 U338 ( .A(n478), .B(KEYINPUT119), .ZN(n548) );
  XOR2_X1 U339 ( .A(n485), .B(KEYINPUT28), .Z(n539) );
  INV_X1 U340 ( .A(G29GAT), .ZN(n455) );
  XNOR2_X1 U341 ( .A(n479), .B(G127GAT), .ZN(n480) );
  XNOR2_X1 U342 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U343 ( .A(n481), .B(n480), .ZN(G1342GAT) );
  XNOR2_X1 U344 ( .A(n458), .B(n457), .ZN(G1328GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT76), .B(KEYINPUT65), .Z(n294) );
  XOR2_X1 U346 ( .A(G50GAT), .B(G162GAT), .Z(n346) );
  XOR2_X1 U347 ( .A(G134GAT), .B(KEYINPUT78), .Z(n328) );
  XNOR2_X1 U348 ( .A(n346), .B(n328), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT64), .B(KEYINPUT77), .Z(n296) );
  XNOR2_X1 U351 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U353 ( .A(KEYINPUT11), .B(KEYINPUT79), .Z(n298) );
  XNOR2_X1 U354 ( .A(KEYINPUT67), .B(KEYINPUT81), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U356 ( .A(n300), .B(n299), .Z(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT80), .B(G218GAT), .Z(n302) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n359) );
  XOR2_X1 U360 ( .A(G85GAT), .B(G92GAT), .Z(n304) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n437) );
  XNOR2_X1 U363 ( .A(n359), .B(n437), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U365 ( .A(n308), .B(n307), .Z(n310) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U368 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n312) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G29GAT), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U371 ( .A(KEYINPUT71), .B(n313), .ZN(n436) );
  XNOR2_X1 U372 ( .A(n314), .B(n436), .ZN(n560) );
  XNOR2_X1 U373 ( .A(KEYINPUT82), .B(n560), .ZN(n547) );
  XOR2_X1 U374 ( .A(KEYINPUT36), .B(n547), .Z(n588) );
  XOR2_X1 U375 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n316) );
  XNOR2_X1 U376 ( .A(G1GAT), .B(G57GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U378 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n318) );
  XNOR2_X1 U379 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U381 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U382 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n322) );
  NAND2_X1 U383 ( .A1(G225GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U385 ( .A(KEYINPUT93), .B(n323), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n333) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G148GAT), .Z(n327) );
  XNOR2_X1 U388 ( .A(G127GAT), .B(G162GAT), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U390 ( .A(n329), .B(n328), .Z(n331) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(G155GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U393 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U394 ( .A(G120GAT), .B(KEYINPUT87), .Z(n335) );
  XNOR2_X1 U395 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n372) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n336), .B(KEYINPUT2), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n372), .B(n341), .ZN(n337) );
  XOR2_X1 U400 ( .A(n338), .B(n337), .Z(n486) );
  INV_X1 U401 ( .A(n486), .ZN(n572) );
  INV_X1 U402 ( .A(KEYINPUT100), .ZN(n394) );
  XOR2_X1 U403 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n340) );
  XNOR2_X1 U404 ( .A(G211GAT), .B(KEYINPUT91), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U406 ( .A(n341), .B(KEYINPUT23), .Z(n343) );
  NAND2_X1 U407 ( .A1(G228GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n353) );
  XOR2_X1 U410 ( .A(G22GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U411 ( .A(n346), .B(n401), .ZN(n348) );
  XNOR2_X1 U412 ( .A(G78GAT), .B(G204GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n347), .B(G148GAT), .ZN(n450) );
  XNOR2_X1 U414 ( .A(n348), .B(n450), .ZN(n349) );
  XOR2_X1 U415 ( .A(G197GAT), .B(KEYINPUT21), .Z(n366) );
  XOR2_X1 U416 ( .A(n349), .B(n366), .Z(n351) );
  XNOR2_X1 U417 ( .A(G218GAT), .B(G106GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n485) );
  XOR2_X1 U420 ( .A(G92GAT), .B(KEYINPUT97), .Z(n355) );
  NAND2_X1 U421 ( .A1(G226GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n358) );
  XOR2_X1 U423 ( .A(KEYINPUT83), .B(G211GAT), .Z(n357) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(G183GAT), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n407) );
  XOR2_X1 U426 ( .A(n358), .B(n407), .Z(n361) );
  XNOR2_X1 U427 ( .A(G204GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U429 ( .A(G176GAT), .B(G64GAT), .Z(n440) );
  XOR2_X1 U430 ( .A(n362), .B(n440), .Z(n369) );
  XOR2_X1 U431 ( .A(KEYINPUT19), .B(KEYINPUT89), .Z(n364) );
  XNOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U434 ( .A(G169GAT), .B(n365), .Z(n384) );
  INV_X1 U435 ( .A(n384), .ZN(n367) );
  XOR2_X1 U436 ( .A(n367), .B(n366), .Z(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n535) );
  XOR2_X1 U438 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n371) );
  XNOR2_X1 U439 ( .A(G183GAT), .B(G176GAT), .ZN(n370) );
  XOR2_X1 U440 ( .A(n371), .B(n370), .Z(n383) );
  XNOR2_X1 U441 ( .A(n372), .B(KEYINPUT90), .ZN(n374) );
  XOR2_X1 U442 ( .A(G99GAT), .B(G190GAT), .Z(n376) );
  XNOR2_X1 U443 ( .A(G43GAT), .B(G134GAT), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U445 ( .A(G15GAT), .B(G127GAT), .Z(n402) );
  XNOR2_X1 U446 ( .A(n377), .B(n402), .ZN(n379) );
  AND2_X1 U447 ( .A1(G227GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n385) );
  INV_X1 U450 ( .A(n490), .ZN(n537) );
  NAND2_X1 U451 ( .A1(n535), .A2(n537), .ZN(n386) );
  XOR2_X1 U452 ( .A(KEYINPUT99), .B(n386), .Z(n387) );
  NAND2_X1 U453 ( .A1(n485), .A2(n387), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n388), .B(KEYINPUT25), .ZN(n392) );
  NOR2_X1 U455 ( .A1(n485), .A2(n537), .ZN(n390) );
  INV_X1 U456 ( .A(n574), .ZN(n551) );
  XOR2_X1 U457 ( .A(n535), .B(KEYINPUT27), .Z(n473) );
  NOR2_X1 U458 ( .A1(n551), .A2(n473), .ZN(n391) );
  NOR2_X1 U459 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n395) );
  NOR2_X1 U461 ( .A1(n572), .A2(n395), .ZN(n497) );
  XOR2_X1 U462 ( .A(G57GAT), .B(KEYINPUT72), .Z(n397) );
  XNOR2_X1 U463 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n449) );
  XOR2_X1 U465 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n399) );
  XNOR2_X1 U466 ( .A(KEYINPUT14), .B(KEYINPUT86), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U468 ( .A(n449), .B(n400), .Z(n404) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n413) );
  XOR2_X1 U471 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n406) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G78GAT), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n411) );
  XOR2_X1 U474 ( .A(n407), .B(G64GAT), .Z(n409) );
  NAND2_X1 U475 ( .A1(G231GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U477 ( .A(n411), .B(n410), .Z(n412) );
  XOR2_X1 U478 ( .A(n413), .B(n412), .Z(n585) );
  INV_X1 U479 ( .A(n539), .ZN(n476) );
  NAND2_X1 U480 ( .A1(n490), .A2(n476), .ZN(n414) );
  NOR2_X1 U481 ( .A1(n473), .A2(n414), .ZN(n415) );
  NOR2_X1 U482 ( .A1(n486), .A2(n415), .ZN(n496) );
  INV_X1 U483 ( .A(n496), .ZN(n416) );
  NAND2_X1 U484 ( .A1(n585), .A2(n416), .ZN(n417) );
  OR2_X1 U485 ( .A1(n497), .A2(n417), .ZN(n418) );
  NOR2_X1 U486 ( .A1(n588), .A2(n418), .ZN(n419) );
  XNOR2_X1 U487 ( .A(KEYINPUT37), .B(n419), .ZN(n530) );
  XOR2_X1 U488 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n421) );
  XNOR2_X1 U489 ( .A(G8GAT), .B(G1GAT), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n434) );
  XOR2_X1 U491 ( .A(G141GAT), .B(G22GAT), .Z(n423) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(G36GAT), .ZN(n422) );
  XNOR2_X1 U493 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U494 ( .A(G113GAT), .B(G15GAT), .Z(n425) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G197GAT), .ZN(n424) );
  XNOR2_X1 U496 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U497 ( .A(n427), .B(n426), .Z(n432) );
  XOR2_X1 U498 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n429) );
  NAND2_X1 U499 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U500 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U501 ( .A(KEYINPUT69), .B(n430), .ZN(n431) );
  XNOR2_X1 U502 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U503 ( .A(n434), .B(n433), .Z(n435) );
  XOR2_X1 U504 ( .A(n436), .B(n435), .Z(n576) );
  INV_X1 U505 ( .A(n576), .ZN(n563) );
  XNOR2_X1 U506 ( .A(n437), .B(KEYINPUT74), .ZN(n439) );
  AND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U508 ( .A(n439), .B(n438), .ZN(n444) );
  XNOR2_X1 U509 ( .A(G120GAT), .B(n440), .ZN(n442) );
  XOR2_X1 U510 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n446) );
  XNOR2_X1 U511 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U513 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U514 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(n581) );
  NAND2_X1 U516 ( .A1(n563), .A2(n581), .ZN(n500) );
  NOR2_X1 U517 ( .A1(n530), .A2(n500), .ZN(n454) );
  XNOR2_X1 U518 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n453) );
  XNOR2_X1 U519 ( .A(n454), .B(n453), .ZN(n517) );
  AND2_X1 U520 ( .A1(n517), .A2(n572), .ZN(n458) );
  XNOR2_X1 U521 ( .A(KEYINPUT39), .B(KEYINPUT107), .ZN(n456) );
  XNOR2_X1 U522 ( .A(n581), .B(KEYINPUT41), .ZN(n565) );
  NAND2_X1 U523 ( .A1(n563), .A2(n565), .ZN(n460) );
  XOR2_X1 U524 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n459) );
  XNOR2_X1 U525 ( .A(n460), .B(n459), .ZN(n462) );
  XOR2_X1 U526 ( .A(KEYINPUT114), .B(n585), .Z(n569) );
  NOR2_X1 U527 ( .A1(n560), .A2(n569), .ZN(n461) );
  NAND2_X1 U528 ( .A1(n462), .A2(n461), .ZN(n464) );
  XNOR2_X1 U529 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n466) );
  NOR2_X1 U530 ( .A1(n588), .A2(n585), .ZN(n465) );
  XNOR2_X1 U531 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U532 ( .A1(n581), .A2(n467), .ZN(n468) );
  NOR2_X1 U533 ( .A1(n563), .A2(n468), .ZN(n469) );
  NOR2_X1 U534 ( .A1(n470), .A2(n469), .ZN(n472) );
  NOR2_X1 U535 ( .A1(n473), .A2(n486), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n482), .A2(n474), .ZN(n552) );
  NOR2_X1 U537 ( .A1(n552), .A2(n490), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n475), .B(KEYINPUT118), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n548), .A2(n569), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n479) );
  INV_X1 U542 ( .A(G190GAT), .ZN(n494) );
  NAND2_X1 U543 ( .A1(n535), .A2(n482), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n573) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  NOR2_X1 U547 ( .A1(n573), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT55), .ZN(n489) );
  NOR2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n570) );
  NAND2_X1 U550 ( .A1(n570), .A2(n547), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1351GAT) );
  NOR2_X1 U554 ( .A1(n585), .A2(n547), .ZN(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT16), .B(n495), .ZN(n499) );
  NOR2_X1 U556 ( .A1(n497), .A2(n496), .ZN(n498) );
  NAND2_X1 U557 ( .A1(n499), .A2(n498), .ZN(n520) );
  NOR2_X1 U558 ( .A1(n500), .A2(n520), .ZN(n509) );
  NAND2_X1 U559 ( .A1(n509), .A2(n572), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(KEYINPUT34), .ZN(n502) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n502), .ZN(G1324GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n504) );
  NAND2_X1 U563 ( .A1(n509), .A2(n535), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G8GAT), .B(n505), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U567 ( .A1(n509), .A2(n537), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U569 ( .A(G15GAT), .B(n508), .Z(G1326GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n511) );
  NAND2_X1 U571 ( .A1(n509), .A2(n539), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G22GAT), .B(n512), .ZN(G1327GAT) );
  NAND2_X1 U574 ( .A1(n517), .A2(n535), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(KEYINPUT108), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G36GAT), .B(n514), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n537), .A2(n517), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(KEYINPUT40), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n516), .ZN(G1330GAT) );
  XOR2_X1 U580 ( .A(G50GAT), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U581 ( .A1(n517), .A2(n539), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1331GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n522) );
  NAND2_X1 U584 ( .A1(n576), .A2(n565), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n531), .A2(n520), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n527), .A2(n572), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(G57GAT), .B(n523), .Z(G1332GAT) );
  XOR2_X1 U589 ( .A(G64GAT), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U590 ( .A1(n527), .A2(n535), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1333GAT) );
  NAND2_X1 U592 ( .A1(n537), .A2(n527), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U595 ( .A1(n527), .A2(n539), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  XOR2_X1 U597 ( .A(G85GAT), .B(KEYINPUT113), .Z(n534) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT112), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n572), .A2(n540), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(G1336GAT) );
  NAND2_X1 U602 ( .A1(n540), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n537), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n538), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(KEYINPUT44), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n542), .ZN(G1339GAT) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(KEYINPUT120), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n563), .A2(n548), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U613 ( .A1(n548), .A2(n565), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n563), .A2(n561), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U623 ( .A1(n561), .A2(n565), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  INV_X1 U626 ( .A(n585), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n563), .A2(n570), .ZN(n564) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NOR2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

