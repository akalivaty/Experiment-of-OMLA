//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G204gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G197gat), .ZN(new_n203));
  INV_X1    g002(.A(G197gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G204gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT68), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n207), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(new_n203), .A3(new_n205), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT72), .A3(new_n217), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n225));
  AND2_X1   g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n220), .A2(new_n224), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  INV_X1    g029(.A(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n225), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n217), .A3(new_n223), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT69), .B(KEYINPUT29), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n237), .A2(KEYINPUT79), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT79), .B1(new_n237), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n215), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G228gat), .A3(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n244), .A3(new_n214), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT77), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n211), .A2(KEYINPUT77), .A3(new_n214), .A4(new_n244), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n236), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n235), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT78), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n253), .A3(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n243), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n213), .A2(new_n210), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n213), .A2(new_n210), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT76), .B1(new_n258), .B2(new_n238), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n238), .B1(new_n256), .B2(new_n257), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT76), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT3), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n250), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n237), .A2(new_n239), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n215), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n264), .A2(new_n266), .B1(G228gat), .B2(G233gat), .ZN(new_n267));
  OAI21_X1  g066(.A(G22gat), .B1(new_n255), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G228gat), .A2(G233gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n237), .A2(KEYINPUT79), .A3(new_n239), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n273), .B2(new_n215), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n229), .A2(new_n235), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT3), .B1(new_n245), .B2(new_n246), .ZN(new_n276));
  AOI211_X1 g075(.A(KEYINPUT78), .B(new_n275), .C1(new_n276), .C2(new_n248), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n253), .B1(new_n249), .B2(new_n250), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G22gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n275), .B1(new_n259), .B2(new_n262), .ZN(new_n281));
  INV_X1    g080(.A(new_n266), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n269), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT31), .B(G50gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n284), .B2(KEYINPUT80), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n268), .B(new_n284), .C1(KEYINPUT80), .C2(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G127gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G134gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(G127gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n294), .B(new_n298), .C1(new_n299), .C2(KEYINPUT1), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(G127gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n294), .B(new_n301), .C1(KEYINPUT65), .C2(KEYINPUT1), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT1), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n250), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT73), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n300), .A2(new_n308), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n237), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(new_n314), .B2(new_n250), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n275), .A2(KEYINPUT4), .A3(new_n309), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n315), .A2(new_n311), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n321));
  XNOR2_X1  g120(.A(G1gat), .B(G29gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT0), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT74), .ZN(new_n324));
  XOR2_X1   g123(.A(G57gat), .B(G85gat), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  INV_X1    g127(.A(new_n311), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n275), .A2(new_n309), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n250), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n319), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n321), .A2(new_n327), .A3(new_n334), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n336), .A2(new_n311), .B1(new_n332), .B2(KEYINPUT5), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n312), .B2(new_n319), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n326), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n335), .A2(new_n340), .A3(KEYINPUT75), .A4(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(new_n327), .C1(new_n344), .C2(KEYINPUT6), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G169gat), .ZN(new_n347));
  INV_X1    g146(.A(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n349), .A2(KEYINPUT26), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n352), .B2(KEYINPUT26), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n350), .A2(new_n353), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT27), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT27), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT64), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT64), .ZN(new_n361));
  AOI21_X1  g160(.A(G190gat), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT28), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n359), .A2(new_n364), .A3(G190gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n354), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  AND2_X1   g166(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(KEYINPUT23), .ZN(new_n370));
  OR2_X1    g169(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(G190gat), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n351), .A2(KEYINPUT23), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n349), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n370), .A2(new_n373), .A3(new_n375), .A4(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n366), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n215), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n366), .B2(new_n380), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n384), .B(new_n385), .C1(new_n383), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT70), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n381), .A2(new_n244), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n382), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(KEYINPUT70), .A3(new_n384), .A4(new_n385), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n238), .B1(new_n366), .B2(new_n380), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n384), .B1(new_n394), .B2(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n215), .ZN(new_n396));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n389), .A2(new_n392), .B1(new_n395), .B2(new_n215), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT71), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT30), .A4(new_n399), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT30), .B1(new_n402), .B2(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n399), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n401), .A2(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n292), .B1(new_n346), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT36), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(KEYINPUT67), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n366), .A2(new_n380), .A3(new_n314), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n314), .B1(new_n366), .B2(new_n380), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G227gat), .ZN(new_n414));
  INV_X1    g213(.A(G233gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT66), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n418));
  INV_X1    g217(.A(new_n416), .ZN(new_n419));
  NOR4_X1   g218(.A1(new_n411), .A2(new_n412), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT32), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n417), .B2(new_n420), .ZN(new_n423));
  XOR2_X1   g222(.A(G15gat), .B(G43gat), .Z(new_n424));
  XNOR2_X1  g223(.A(G71gat), .B(G99gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n411), .B2(new_n412), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n428), .A2(KEYINPUT34), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(KEYINPUT34), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n426), .ZN(new_n432));
  OAI221_X1 g231(.A(KEYINPUT32), .B1(new_n422), .B2(new_n432), .C1(new_n417), .C2(new_n420), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n427), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n410), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(new_n431), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT67), .B(KEYINPUT36), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n408), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n401), .A2(new_n404), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n405), .A2(new_n406), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n335), .A2(KEYINPUT81), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n343), .A2(new_n449), .A3(new_n327), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OR3_X1    g250(.A1(new_n336), .A2(KEYINPUT39), .A3(new_n311), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n310), .A2(new_n311), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT39), .B(new_n453), .C1(new_n336), .C2(new_n311), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n326), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n447), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n395), .B2(new_n385), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n391), .A2(new_n384), .A3(new_n215), .ZN(new_n463));
  AOI211_X1 g262(.A(KEYINPUT38), .B(new_n399), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n402), .A2(KEYINPUT82), .A3(new_n461), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT82), .B1(new_n402), .B2(new_n461), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n327), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n448), .A2(new_n450), .A3(new_n341), .A4(new_n340), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n468), .A2(new_n406), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n393), .A2(new_n396), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(KEYINPUT37), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n465), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n399), .B1(new_n474), .B2(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n460), .B(new_n292), .C1(new_n471), .C2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n292), .A2(new_n439), .A3(new_n440), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n407), .A2(new_n346), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT35), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT35), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n470), .A2(new_n469), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n407), .A3(new_n292), .A4(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n444), .A2(new_n479), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT11), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(G169gat), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT83), .B(G197gat), .Z(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n489), .B(new_n347), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT12), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n280), .A2(G15gat), .ZN(new_n499));
  INV_X1    g298(.A(G15gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G22gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G1gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(G1gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(new_n499), .A3(new_n501), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n503), .B2(new_n506), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  INV_X1    g310(.A(G43gat), .ZN(new_n512));
  INV_X1    g311(.A(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G43gat), .A2(G50gat), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(G29gat), .ZN(new_n518));
  INV_X1    g317(.A(G36gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n518), .A2(new_n519), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n520), .A2(new_n521), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n514), .A2(new_n526), .A3(new_n515), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(KEYINPUT15), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT15), .B1(new_n525), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n511), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n528), .A4(new_n524), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n510), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT85), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n529), .A2(new_n530), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n510), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n535), .B(new_n510), .C1(new_n531), .C2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n524), .A2(new_n528), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n510), .A2(new_n543), .A3(new_n532), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n529), .A2(new_n530), .B1(new_n508), .B2(new_n509), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n540), .B(KEYINPUT13), .Z(new_n547));
  AOI22_X1  g346(.A1(new_n542), .A2(KEYINPUT18), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(new_n540), .C1(new_n534), .C2(new_n537), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n498), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n538), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n540), .A4(new_n549), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n546), .A2(new_n547), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n552), .A2(new_n555), .A3(new_n498), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n486), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(G57gat), .A2(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G57gat), .A2(G64gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n565), .ZN(new_n571));
  NOR2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n564), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G57gat), .B(G64gat), .Z(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n575), .A2(KEYINPUT87), .A3(new_n576), .A4(new_n567), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n565), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n575), .B2(new_n567), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n565), .B1(new_n572), .B2(new_n578), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n574), .A2(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n563), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n562), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n584), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n561), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n584), .A2(new_n589), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n597));
  INV_X1    g396(.A(new_n561), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n582), .A2(KEYINPUT21), .ZN(new_n600));
  INV_X1    g399(.A(new_n510), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n593), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n593), .B2(new_n599), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT89), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n599), .ZN(new_n610));
  INV_X1    g409(.A(new_n602), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n607), .B1(new_n612), .B2(new_n603), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G134gat), .B(G162gat), .Z(new_n615));
  OR2_X1    g414(.A1(KEYINPUT90), .A2(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(KEYINPUT90), .A2(G85gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n620));
  NAND2_X1  g419(.A1(G85gat), .A2(G92gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(KEYINPUT8), .ZN(new_n623));
  XNOR2_X1  g422(.A(G99gat), .B(G106gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n619), .A2(new_n623), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(KEYINPUT8), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(new_n620), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n627), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n629), .B2(new_n619), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n626), .B1(new_n630), .B2(KEYINPUT91), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n626), .A2(KEYINPUT91), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT92), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n531), .A2(new_n533), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT92), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n636), .A3(new_n632), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT93), .ZN(new_n639));
  NAND3_X1  g438(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n543), .A2(new_n532), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n639), .B(new_n640), .C1(new_n633), .C2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n536), .A2(new_n631), .A3(new_n632), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n639), .B1(new_n644), .B2(new_n640), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n638), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n647), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n638), .B(new_n651), .C1(new_n643), .C2(new_n645), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n648), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n615), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n649), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n658));
  INV_X1    g457(.A(new_n615), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n614), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT94), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT94), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n614), .A2(new_n655), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n631), .A2(new_n587), .A3(new_n632), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n667));
  INV_X1    g466(.A(new_n624), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT95), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n667), .B2(KEYINPUT95), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n582), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT10), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n631), .A2(new_n582), .A3(KEYINPUT10), .A4(new_n632), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n665), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n665), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n666), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(G120gat), .B(G148gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT96), .ZN(new_n681));
  XOR2_X1   g480(.A(G176gat), .B(G204gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n676), .A2(new_n678), .A3(new_n683), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n679), .A2(KEYINPUT97), .A3(new_n684), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n662), .A2(new_n664), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n560), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n346), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT99), .B(G1gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1324gat));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n447), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n700), .B2(new_n507), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n504), .A2(new_n507), .ZN(new_n702));
  NAND2_X1  g501(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  MUX2_X1   g503(.A(KEYINPUT42), .B(new_n701), .S(new_n704), .Z(G1325gat));
  INV_X1    g504(.A(new_n694), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n443), .B(KEYINPUT100), .Z(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n434), .A2(new_n435), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n500), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT101), .Z(G1326gat));
  INV_X1    g512(.A(new_n292), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  AND2_X1   g516(.A1(new_n655), .A2(new_n660), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n486), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n690), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n614), .A2(new_n559), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n518), .A3(new_n695), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n486), .B2(new_n718), .ZN(new_n726));
  INV_X1    g525(.A(new_n718), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n445), .A2(new_n346), .A3(new_n446), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n442), .B(new_n436), .C1(new_n728), .C2(new_n292), .ZN(new_n729));
  INV_X1    g528(.A(new_n478), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n470), .A2(new_n469), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n730), .A2(new_n406), .A3(new_n731), .A4(new_n468), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n451), .A2(new_n458), .A3(new_n457), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n714), .B1(new_n447), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n729), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n439), .A2(new_n440), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n731), .A2(new_n736), .A3(KEYINPUT35), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n714), .A2(new_n447), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n710), .A2(new_n346), .A3(new_n292), .A4(new_n407), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(KEYINPUT35), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT44), .B(new_n727), .C1(new_n735), .C2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n726), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n721), .ZN(new_n743));
  OAI21_X1  g542(.A(G29gat), .B1(new_n743), .B2(new_n346), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n744), .ZN(G1328gat));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n519), .A3(new_n447), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT102), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n743), .B2(new_n407), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  OAI21_X1  g549(.A(G43gat), .B1(new_n743), .B2(new_n708), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n722), .A2(new_n512), .A3(new_n710), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n443), .ZN(new_n755));
  OAI21_X1  g554(.A(G43gat), .B1(new_n743), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n753), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(new_n752), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT103), .ZN(G1330gat));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n513), .A3(new_n292), .ZN(new_n760));
  AOI21_X1  g559(.A(G50gat), .B1(new_n722), .B2(new_n714), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT48), .Z(G1331gat));
  NAND4_X1  g562(.A1(new_n662), .A2(new_n664), .A3(new_n720), .A4(new_n559), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n486), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n695), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768));
  INV_X1    g567(.A(G64gat), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n765), .B(new_n447), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1333gat));
  NAND3_X1  g571(.A1(new_n765), .A2(G71gat), .A3(new_n707), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n486), .A2(new_n736), .A3(new_n764), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G71gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n765), .A2(new_n714), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n444), .A2(new_n479), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n482), .A2(new_n485), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n559), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n614), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n727), .A4(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n727), .B(new_n783), .C1(new_n735), .C2(new_n740), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(KEYINPUT104), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(KEYINPUT104), .B2(new_n787), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n690), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(new_n695), .A3(new_n616), .A4(new_n618), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n616), .A2(new_n618), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n782), .A2(new_n614), .A3(new_n690), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n742), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n794), .B2(new_n346), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(G1336gat));
  OAI21_X1  g595(.A(G92gat), .B1(new_n794), .B2(new_n407), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n407), .A2(G92gat), .A3(new_n690), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n797), .B(new_n798), .C1(new_n789), .C2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n787), .ZN(new_n802));
  INV_X1    g601(.A(new_n784), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n798), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(G1337gat));
  INV_X1    g608(.A(G99gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n810), .A3(new_n710), .ZN(new_n811));
  OAI21_X1  g610(.A(G99gat), .B1(new_n794), .B2(new_n708), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n726), .A2(new_n741), .A3(new_n714), .A4(new_n793), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n292), .A2(G106gat), .A3(new_n690), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n814), .B(new_n816), .C1(new_n789), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT107), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n787), .B2(new_n784), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n816), .B2(KEYINPUT106), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT106), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n823), .A3(G106gat), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n820), .B(new_n814), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n816), .A2(KEYINPUT106), .ZN(new_n826));
  INV_X1    g625(.A(new_n821), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT107), .B1(new_n828), .B2(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n819), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n832), .B(new_n819), .C1(new_n825), .C2(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n835));
  AND4_X1   g634(.A1(new_n662), .A2(new_n664), .A3(new_n690), .A4(new_n559), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  INV_X1    g636(.A(new_n673), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n674), .A3(new_n677), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(new_n676), .A3(KEYINPUT54), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n684), .B1(new_n676), .B2(KEYINPUT54), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n676), .A3(KEYINPUT54), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n676), .A2(KEYINPUT54), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT55), .A4(new_n684), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n687), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n847));
  INV_X1    g646(.A(new_n547), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n544), .A2(new_n545), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n496), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g654(.A(KEYINPUT110), .B(new_n496), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n557), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n559), .A2(new_n846), .B1(new_n857), .B2(new_n690), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n718), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n655), .B2(new_n660), .ZN(new_n860));
  INV_X1    g659(.A(new_n846), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n614), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n835), .B1(new_n836), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n662), .A2(new_n664), .A3(new_n690), .A4(new_n559), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n718), .A2(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(KEYINPUT111), .C1(new_n866), .C2(new_n614), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n447), .A2(new_n346), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n480), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n782), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n870), .A2(new_n874), .A3(new_n871), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n559), .A2(new_n305), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(G1340gat));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n303), .A3(new_n720), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n720), .B1(new_n875), .B2(new_n877), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(KEYINPUT113), .A3(G120gat), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT113), .B1(new_n883), .B2(G120gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1341gat));
  NAND3_X1  g685(.A1(new_n872), .A2(new_n293), .A3(new_n614), .ZN(new_n887));
  INV_X1    g686(.A(new_n614), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n876), .B2(new_n878), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n293), .ZN(G1342gat));
  NAND4_X1  g689(.A1(new_n870), .A2(new_n297), .A3(new_n727), .A4(new_n871), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT114), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(KEYINPUT114), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n893), .A2(new_n894), .B1(KEYINPUT56), .B2(new_n891), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n718), .B1(new_n876), .B2(new_n878), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n297), .B2(new_n896), .ZN(G1343gat));
  XNOR2_X1  g696(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n707), .A2(new_n292), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n868), .A2(new_n869), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n559), .A2(G141gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n292), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n858), .A2(new_n906), .A3(new_n718), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n862), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n858), .B2(new_n718), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n888), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n910), .B2(new_n865), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n864), .A2(new_n714), .A3(new_n867), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n903), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n755), .A2(new_n869), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n559), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n915), .B2(new_n230), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n912), .A2(new_n903), .ZN(new_n918));
  INV_X1    g717(.A(new_n911), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n921));
  INV_X1    g720(.A(new_n914), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT116), .B1(new_n913), .B2(new_n914), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n782), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n917), .B1(new_n925), .B2(G141gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n916), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT118), .B(new_n916), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1344gat));
  XNOR2_X1  g731(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n863), .B1(new_n693), .B2(new_n559), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(KEYINPUT57), .A3(new_n292), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n912), .A2(KEYINPUT57), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n914), .A2(new_n690), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(KEYINPUT120), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G148gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT120), .B1(new_n937), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n231), .A2(KEYINPUT59), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n924), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n690), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR4_X1   g745(.A1(new_n447), .A2(G148gat), .A3(new_n346), .A4(new_n690), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n868), .A2(new_n899), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1345gat));
  OAI21_X1  g748(.A(G155gat), .B1(new_n944), .B2(new_n888), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n900), .A2(new_n221), .A3(new_n614), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1346gat));
  OAI21_X1  g751(.A(G162gat), .B1(new_n944), .B2(new_n718), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n900), .A2(new_n222), .A3(new_n727), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n407), .A2(new_n695), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT122), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n871), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n868), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(new_n347), .A3(new_n559), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n864), .A2(new_n346), .A3(new_n867), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT121), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(new_n447), .A3(new_n871), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n782), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n960), .B1(new_n964), .B2(new_n347), .ZN(G1348gat));
  NAND3_X1  g764(.A1(new_n963), .A2(new_n348), .A3(new_n720), .ZN(new_n966));
  OAI21_X1  g765(.A(G176gat), .B1(new_n959), .B2(new_n690), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1349gat));
  NAND4_X1  g767(.A1(new_n963), .A2(new_n614), .A3(new_n356), .A4(new_n358), .ZN(new_n969));
  OAI21_X1  g768(.A(G183gat), .B1(new_n959), .B2(new_n888), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n963), .A2(new_n367), .A3(new_n727), .ZN(new_n973));
  OAI21_X1  g772(.A(G190gat), .B1(new_n959), .B2(new_n718), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1351gat));
  NAND2_X1  g775(.A1(new_n708), .A2(new_n957), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n937), .A2(new_n978), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n979), .A2(new_n204), .A3(new_n559), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n707), .A2(new_n407), .A3(new_n292), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT123), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n962), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(new_n782), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n980), .B1(new_n986), .B2(new_n204), .ZN(G1352gat));
  NOR3_X1   g786(.A1(new_n982), .A2(G204gat), .A3(new_n690), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  OAI21_X1  g788(.A(G204gat), .B1(new_n979), .B2(new_n690), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1353gat));
  INV_X1    g790(.A(G211gat), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n977), .A2(new_n888), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n937), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT63), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n983), .A2(new_n992), .A3(new_n614), .A4(new_n985), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1354gat));
  NAND2_X1  g796(.A1(new_n727), .A2(G218gat), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT126), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n979), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n727), .A3(new_n985), .ZN(new_n1001));
  INV_X1    g800(.A(G218gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1001), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(G1355gat));
endmodule


