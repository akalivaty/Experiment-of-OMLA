//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT27), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT69), .A3(G116), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n197), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  AOI21_X1  g022(.A(G131), .B1(new_n207), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n208), .A2(new_n209), .A3(new_n214), .A4(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n213), .A2(new_n215), .B1(G131), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT64), .B1(new_n223), .B2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(G146), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT65), .B1(new_n223), .B2(G146), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n221), .A3(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n223), .A2(G146), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .A4(new_n227), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n205), .B1(new_n219), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n231), .A2(new_n233), .A3(new_n234), .A4(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n242));
  OAI21_X1  g056(.A(G128), .B1(new_n225), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n226), .A2(KEYINPUT68), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT68), .B1(new_n226), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n210), .A2(G134), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(new_n216), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n213), .B2(new_n215), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT28), .B1(new_n238), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n241), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n226), .A2(new_n243), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n226), .A2(KEYINPUT68), .A3(new_n243), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n213), .A2(new_n215), .ZN(new_n259));
  INV_X1    g073(.A(new_n249), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n246), .A2(new_n263), .A3(new_n250), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n262), .A2(new_n238), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n205), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(KEYINPUT67), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n250), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n246), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n218), .A2(new_n236), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n266), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT28), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n252), .B1(new_n274), .B2(KEYINPUT72), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(KEYINPUT28), .C1(new_n265), .C2(new_n273), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n193), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n262), .A2(KEYINPUT30), .A3(new_n272), .A4(new_n264), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n268), .B1(new_n259), .B2(new_n260), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n258), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n271), .B1(new_n281), .B2(new_n269), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n279), .B(new_n205), .C1(new_n282), .C2(KEYINPUT30), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n262), .A2(new_n238), .A3(new_n264), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n192), .A2(KEYINPUT71), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n278), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(G472), .A3(G902), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n278), .B2(new_n291), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n298));
  INV_X1    g112(.A(new_n252), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n298), .A2(new_n193), .A3(new_n277), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n283), .A2(new_n284), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n301), .B2(new_n192), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n262), .A2(new_n272), .A3(new_n264), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n284), .B1(new_n304), .B2(new_n266), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n252), .B1(new_n305), .B2(KEYINPUT28), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G472), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n311), .B(new_n295), .C1(new_n278), .C2(new_n291), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n294), .A2(new_n297), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G125), .B(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n221), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT24), .B(G110), .Z(new_n316));
  NAND2_X1  g130(.A1(new_n239), .A2(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n199), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n316), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n199), .A2(G128), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n318), .B(new_n324), .C1(new_n325), .C2(KEYINPUT23), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G110), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n315), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G140), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(KEYINPUT76), .A3(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT16), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n221), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n320), .A2(new_n322), .A3(new_n316), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n326), .A2(G110), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n338), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G146), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n221), .A3(new_n338), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT78), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n346), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n341), .B(new_n342), .C1(new_n349), .C2(new_n339), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n345), .B(new_n315), .C1(new_n327), .C2(new_n323), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT77), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G137), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n348), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n350), .A2(new_n351), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT78), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT74), .B(G217), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G902), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(G234), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G902), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT79), .Z(new_n369));
  NAND2_X1  g183(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n363), .A2(new_n366), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n366), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n331), .B(new_n241), .C1(new_n244), .C2(new_n245), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n236), .A2(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G224), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G953), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT7), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n378), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n385), .ZN(new_n387));
  AOI211_X1 g201(.A(KEYINPUT85), .B(new_n387), .C1(new_n379), .C2(new_n380), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G110), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT8), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G104), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(G107), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n392), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n199), .A3(G116), .ZN(new_n406));
  OAI211_X1 g220(.A(G113), .B(new_n406), .C1(new_n202), .C2(new_n405), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n407), .A3(new_n201), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n404), .B1(new_n201), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n391), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(G101), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n205), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n408), .A3(new_n390), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n379), .A2(new_n380), .A3(new_n387), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n389), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n408), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n390), .B(KEYINPUT83), .Z(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n418), .A2(KEYINPUT6), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n424), .A2(new_n425), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n381), .A2(new_n383), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT84), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n418), .A2(KEYINPUT6), .B1(new_n424), .B2(new_n425), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n425), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT84), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n422), .B(new_n423), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n423), .B(KEYINPUT86), .Z(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n386), .A2(new_n388), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n366), .B1(new_n441), .B2(new_n420), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n445), .B2(new_n436), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n438), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n334), .A2(new_n335), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT87), .B(new_n315), .C1(new_n448), .C2(new_n221), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT18), .A2(G131), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n451));
  AOI21_X1  g265(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G237), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n354), .A3(G214), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n223), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(KEYINPUT18), .A3(G131), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n334), .A2(new_n460), .A3(G146), .A4(new_n335), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n392), .ZN(new_n464));
  OAI21_X1  g278(.A(G131), .B1(new_n451), .B2(new_n452), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n247), .A3(new_n457), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n345), .A2(new_n346), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT17), .B(G131), .C1(new_n451), .C2(new_n452), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n462), .B(new_n464), .C1(new_n469), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n462), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n465), .A2(new_n475), .A3(new_n467), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n465), .B2(new_n467), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n476), .A2(new_n477), .A3(new_n339), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n334), .A2(KEYINPUT19), .A3(new_n335), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT19), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n314), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(KEYINPUT89), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(KEYINPUT89), .B2(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n221), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n474), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n473), .B1(new_n485), .B2(new_n464), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  INV_X1    g304(.A(G475), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n462), .B1(new_n469), .B2(new_n472), .ZN(new_n492));
  INV_X1    g306(.A(new_n464), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n494), .B2(new_n473), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n489), .A2(new_n490), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G478), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n223), .A2(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n239), .A2(G143), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n207), .ZN(new_n502));
  INV_X1    g316(.A(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G116), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n196), .A2(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G107), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n505), .A3(new_n395), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT13), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n501), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT13), .B1(new_n223), .B2(G128), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n510), .B1(new_n239), .B2(G143), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n502), .B(new_n509), .C1(new_n517), .C2(new_n207), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n239), .A2(G143), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n223), .A2(G128), .ZN(new_n520));
  OAI21_X1  g334(.A(G134), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n506), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n521), .A2(new_n502), .B1(new_n522), .B2(new_n395), .ZN(new_n523));
  OR3_X1    g337(.A1(new_n503), .A2(KEYINPUT14), .A3(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n505), .A2(KEYINPUT14), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n504), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT9), .B(G234), .Z(new_n529));
  INV_X1    g343(.A(KEYINPUT80), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT9), .B(G234), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT80), .ZN(new_n533));
  AND4_X1   g347(.A1(new_n354), .A2(new_n531), .A3(new_n364), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n518), .B2(new_n528), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n520), .B1(KEYINPUT13), .B2(new_n519), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n512), .A2(new_n513), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G134), .ZN(new_n543));
  INV_X1    g357(.A(new_n502), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n507), .B2(new_n508), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n543), .A2(new_n545), .B1(new_n523), .B2(new_n527), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n546), .A2(KEYINPUT92), .A3(new_n534), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n366), .B(new_n499), .C1(new_n538), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT92), .B1(new_n546), .B2(new_n534), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n518), .A2(new_n528), .ZN(new_n551));
  INV_X1    g365(.A(new_n534), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n537), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n553), .A3(new_n535), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n499), .B1(new_n554), .B2(new_n366), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G952), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  NAND2_X1  g372(.A1(G234), .A2(G237), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(G902), .A3(G953), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n556), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n496), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G214), .B1(G237), .B2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n447), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n241), .B(new_n403), .C1(new_n244), .C2(new_n245), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n243), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n241), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n404), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n218), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n403), .B1(new_n241), .B2(new_n574), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT82), .B1(new_n580), .B2(KEYINPUT10), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT82), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n403), .A2(new_n583), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n416), .A2(new_n230), .A3(new_n235), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n246), .A2(new_n586), .B1(new_n587), .B2(new_n414), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n588), .A3(new_n218), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n354), .A2(G227), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT81), .ZN(new_n591));
  XNOR2_X1  g405(.A(G110), .B(G140), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n579), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n588), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n219), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n598), .B2(new_n589), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n571), .B(new_n366), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n589), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n593), .B1(new_n579), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n594), .A3(new_n589), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(G469), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(G469), .A2(G902), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n531), .A2(new_n533), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n366), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(G221), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n570), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n313), .A2(new_n377), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT93), .B(G101), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  INV_X1    g429(.A(KEYINPUT28), .ZN(new_n616));
  AOI211_X1 g430(.A(KEYINPUT67), .B(new_n249), .C1(new_n213), .C2(new_n215), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n258), .A2(new_n280), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n205), .B1(new_n618), .B2(new_n271), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n284), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n299), .B1(new_n620), .B2(new_n276), .ZN(new_n621));
  INV_X1    g435(.A(new_n277), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n192), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n283), .A2(new_n289), .A3(new_n286), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n289), .B1(new_n283), .B2(new_n286), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n366), .B1(new_n278), .B2(new_n291), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT94), .B1(new_n631), .B2(G472), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n292), .A2(new_n377), .A3(new_n610), .A4(new_n606), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n494), .A2(new_n473), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n491), .B1(new_n636), .B2(new_n366), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n486), .A2(new_n488), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT20), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  INV_X1    g456(.A(new_n536), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n546), .B2(new_n534), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n554), .A2(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n497), .A2(G902), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n366), .B1(new_n538), .B2(new_n547), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n645), .A2(new_n646), .B1(new_n497), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n635), .B1(new_n641), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n496), .A2(new_n650), .A3(KEYINPUT96), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n422), .B1(new_n433), .B2(new_n437), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n655));
  INV_X1    g469(.A(new_n423), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n438), .A2(KEYINPUT95), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n445), .A2(new_n436), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n423), .B1(new_n659), .B2(new_n422), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n569), .B(new_n657), .C1(new_n658), .C2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n653), .A2(new_n661), .A3(new_n565), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n633), .A2(new_n634), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n637), .B1(new_n489), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n640), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n556), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n654), .A2(new_n656), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(KEYINPUT95), .A3(new_n438), .ZN(new_n672));
  INV_X1    g486(.A(new_n569), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n660), .B2(new_n655), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n566), .A2(new_n670), .A3(new_n672), .A4(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n633), .A2(new_n634), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  AOI21_X1  g492(.A(KEYINPUT25), .B1(new_n363), .B2(new_n366), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n373), .B(G902), .C1(new_n360), .C2(new_n362), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n367), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n359), .A2(KEYINPUT36), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n361), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n369), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n606), .A3(new_n610), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n570), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n687), .B(new_n292), .C1(new_n632), .C2(new_n630), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT98), .B(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n561), .B1(new_n692), .B2(new_n563), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n670), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n691), .B1(new_n695), .B2(new_n661), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n669), .A2(new_n556), .A3(new_n693), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(KEYINPUT99), .A3(new_n672), .A4(new_n674), .ZN(new_n698));
  INV_X1    g512(.A(new_n686), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n313), .A2(new_n696), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  AND2_X1   g515(.A1(new_n606), .A2(new_n610), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n693), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT102), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT40), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n447), .B(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n496), .B1(new_n555), .B2(new_n549), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n710), .A2(new_n673), .A3(new_n685), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n366), .B1(new_n305), .B2(new_n193), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n192), .B1(new_n283), .B2(new_n284), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n294), .A2(new_n717), .A3(new_n297), .A4(new_n312), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n707), .A2(new_n708), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  NAND2_X1  g534(.A1(new_n496), .A2(new_n650), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n693), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n661), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n313), .A2(new_n699), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT103), .B(G146), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G48));
  OAI21_X1  g541(.A(new_n366), .B1(new_n596), .B2(new_n599), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n610), .A3(new_n600), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n662), .A2(new_n313), .A3(new_n377), .A4(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT41), .B(G113), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT105), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT104), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n732), .B(new_n735), .ZN(G15));
  NAND2_X1  g550(.A1(new_n681), .A2(new_n370), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n297), .A2(new_n312), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n293), .A2(new_n292), .B1(new_n309), .B2(G472), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n675), .A4(new_n731), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n313), .A2(new_n377), .A3(new_n675), .A4(new_n731), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G116), .ZN(G18));
  NAND2_X1  g560(.A1(new_n685), .A2(new_n568), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n661), .A2(new_n747), .A3(new_n730), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n313), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NOR2_X1   g564(.A1(new_n661), .A2(new_n565), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n737), .B(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT107), .B(G472), .Z(new_n754));
  OAI21_X1  g568(.A(new_n626), .B1(new_n193), .B2(new_n306), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n631), .A2(new_n754), .B1(new_n755), .B2(new_n187), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n730), .A2(new_n711), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n751), .A2(new_n753), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT109), .B(G122), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G24));
  NOR2_X1   g574(.A1(new_n661), .A2(new_n730), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n685), .A3(new_n722), .A4(new_n756), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n447), .B2(new_n673), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n654), .A2(new_n439), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n569), .A4(new_n438), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n765), .A2(new_n702), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n313), .A3(new_n377), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n294), .A2(new_n310), .A3(new_n296), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n768), .A2(new_n722), .A3(new_n771), .A4(new_n753), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n769), .A2(new_n770), .B1(new_n772), .B2(KEYINPUT42), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n740), .A2(new_n775), .A3(new_n697), .A4(new_n768), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n768), .A2(new_n313), .A3(new_n377), .A4(new_n697), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT111), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  AND2_X1   g594(.A1(new_n765), .A2(new_n767), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n633), .A2(new_n292), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n641), .A2(new_n650), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(KEYINPUT112), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n787));
  MUX2_X1   g601(.A(new_n784), .B(new_n786), .S(new_n787), .Z(new_n788));
  NAND3_X1  g602(.A1(new_n783), .A2(new_n685), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n602), .A2(new_n603), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n571), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n605), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n605), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n600), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n610), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n703), .ZN(new_n803));
  OR4_X1    g617(.A1(new_n782), .A2(new_n791), .A3(new_n792), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  OR4_X1    g619(.A1(new_n313), .A2(new_n782), .A3(new_n377), .A4(new_n723), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n329), .ZN(G42));
  NAND2_X1  g624(.A1(new_n788), .A2(new_n561), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n782), .A2(new_n730), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n771), .A2(new_n753), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT122), .B(KEYINPUT48), .Z(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n755), .A2(new_n187), .ZN(new_n819));
  INV_X1    g633(.A(new_n754), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n627), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n737), .B(KEYINPUT108), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n761), .ZN(new_n825));
  INV_X1    g639(.A(new_n718), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n813), .A2(new_n377), .A3(new_n561), .A4(new_n826), .ZN(new_n827));
  OAI221_X1 g641(.A(new_n558), .B1(new_n824), .B2(new_n825), .C1(new_n827), .C2(new_n653), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n824), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n807), .A2(new_n808), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n729), .A2(new_n600), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n610), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n781), .B(new_n830), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n827), .A2(new_n496), .A3(new_n650), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n756), .A2(new_n685), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n814), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n710), .A2(new_n673), .A3(new_n731), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n824), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n839), .ZN(new_n842));
  INV_X1    g656(.A(new_n840), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n830), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n834), .B(new_n838), .C1(new_n841), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n829), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n838), .B1(new_n844), .B2(new_n841), .ZN(new_n848));
  INV_X1    g662(.A(new_n834), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n845), .A2(new_n852), .A3(new_n846), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n847), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n661), .A2(new_n711), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n611), .A2(new_n685), .A3(new_n693), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n718), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n700), .A2(new_n725), .A3(new_n857), .A4(new_n762), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n858), .B(KEYINPUT52), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n861), .B2(new_n859), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n447), .A2(new_n569), .A3(new_n566), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n549), .B2(new_n555), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n647), .A2(new_n498), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(KEYINPUT115), .A3(new_n548), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n641), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n634), .B(new_n871), .C1(new_n630), .C2(new_n632), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n688), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n688), .B2(new_n872), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n641), .B2(new_n648), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n496), .A2(new_n650), .A3(KEYINPUT114), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n863), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n634), .B(new_n881), .C1(new_n632), .C2(new_n630), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n613), .A2(new_n749), .A3(new_n882), .A4(new_n758), .ZN(new_n883));
  INV_X1    g697(.A(new_n732), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n876), .A2(new_n885), .A3(new_n745), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n669), .A2(new_n693), .A3(new_n868), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n313), .A2(new_n699), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n836), .A2(new_n611), .A3(new_n723), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n781), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n779), .A2(new_n773), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n862), .A2(KEYINPUT53), .A3(new_n886), .A4(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n661), .A2(new_n565), .A3(new_n730), .A4(new_n711), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n823), .A2(new_n895), .B1(new_n313), .B2(new_n748), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n613), .A3(new_n732), .A4(new_n882), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n897), .A2(new_n875), .A3(new_n874), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n892), .A2(new_n898), .A3(new_n899), .A4(new_n745), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n876), .A2(new_n885), .A3(new_n745), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n779), .A2(new_n773), .A3(new_n891), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT117), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n861), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n893), .B(new_n894), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n899), .B1(new_n886), .B2(new_n892), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT117), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n862), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n910), .A2(new_n911), .B1(new_n904), .B2(new_n906), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n854), .B(new_n907), .C1(new_n894), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n557), .A2(new_n354), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n822), .A2(new_n609), .A3(new_n673), .A4(new_n784), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT113), .Z(new_n917));
  XOR2_X1   g731(.A(new_n832), .B(KEYINPUT49), .Z(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n826), .A3(new_n710), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(G75));
  XOR2_X1   g734(.A(new_n429), .B(new_n432), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  INV_X1    g736(.A(new_n861), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n908), .B2(new_n909), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n905), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n366), .B1(new_n925), .B2(new_n893), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G210), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n904), .A2(new_n906), .ZN(new_n930));
  INV_X1    g744(.A(new_n893), .ZN(new_n931));
  OAI211_X1 g745(.A(G902), .B(new_n439), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n928), .A3(new_n922), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n354), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n929), .A2(new_n936), .ZN(G51));
  XOR2_X1   g751(.A(new_n605), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n894), .B1(new_n925), .B2(new_n893), .ZN(new_n939));
  INV_X1    g753(.A(new_n907), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n596), .A2(new_n599), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n926), .B(new_n795), .C1(new_n794), .C2(new_n793), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n934), .B1(new_n943), .B2(new_n944), .ZN(G54));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  AND2_X1   g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  OAI211_X1 g761(.A(G902), .B(new_n947), .C1(new_n930), .C2(new_n931), .ZN(new_n948));
  INV_X1    g762(.A(new_n486), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n934), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n926), .A2(KEYINPUT123), .A3(new_n486), .A4(new_n947), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(G60));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n645), .B(new_n956), .C1(new_n939), .C2(new_n940), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n935), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n907), .B1(new_n912), .B2(new_n894), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n645), .B1(new_n959), .B2(new_n956), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n683), .B(new_n964), .C1(new_n930), .C2(new_n931), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n925), .B2(new_n893), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n363), .B(KEYINPUT124), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n965), .B(new_n935), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n964), .B1(new_n930), .B2(new_n931), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n934), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n965), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(G66));
  XNOR2_X1  g789(.A(new_n886), .B(KEYINPUT125), .ZN(new_n976));
  NAND2_X1  g790(.A1(G224), .A2(G953), .ZN(new_n977));
  OAI22_X1  g791(.A1(new_n976), .A2(G953), .B1(new_n564), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(G898), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n429), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  OAI21_X1  g795(.A(new_n279), .B1(new_n282), .B2(KEYINPUT30), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT126), .Z(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(new_n483), .Z(new_n984));
  INV_X1    g798(.A(new_n719), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n700), .A2(new_n725), .A3(new_n762), .ZN(new_n986));
  OR3_X1    g800(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT62), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n704), .B(new_n782), .C1(new_n880), .C2(new_n870), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n809), .B1(new_n740), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n987), .A2(new_n804), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n984), .B1(new_n991), .B2(new_n354), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n779), .A2(new_n773), .ZN(new_n993));
  NOR4_X1   g807(.A1(new_n803), .A2(new_n661), .A3(new_n711), .A4(new_n815), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n809), .A2(new_n994), .A3(new_n986), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n804), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(G953), .ZN(new_n997));
  INV_X1    g811(.A(new_n984), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n992), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G227), .A2(G900), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(G953), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1000), .B(new_n1002), .ZN(G72));
  NOR2_X1   g817(.A1(new_n991), .A2(new_n976), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT63), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n714), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n301), .A2(new_n193), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT127), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n996), .A2(new_n976), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n1006), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n935), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n912), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1008), .A2(new_n714), .A3(new_n1006), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(G57));
endmodule


