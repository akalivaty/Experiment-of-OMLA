//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n202), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(G77), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G244), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n214), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n213), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT64), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n229), .B(new_n233), .C1(new_n228), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n222), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT66), .Z(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n217), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G222), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n225), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(G1698), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n255), .B1(new_n256), .B2(new_n253), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n259), .B2(new_n260), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n266), .A2(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(new_n216), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n265), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G179), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n209), .B1(new_n213), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(new_n269), .A3(G13), .A4(G20), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(G1), .B2(new_n210), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  OR3_X1    g0087(.A1(new_n286), .A2(new_n287), .A3(new_n202), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n203), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n210), .A2(G33), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n289), .B1(new_n290), .B2(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n281), .A2(new_n283), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(new_n279), .B1(new_n202), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n265), .A2(new_n275), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G169), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n277), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n276), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT71), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n300), .B2(G190), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n298), .B(KEYINPUT9), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n303), .A2(new_n305), .A3(new_n309), .A4(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n217), .A2(G20), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n312), .B1(new_n294), .B2(new_n313), .C1(new_n292), .C2(new_n202), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n279), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT11), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n296), .A2(new_n217), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT12), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n284), .B(G68), .C1(G1), .C2(new_n210), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n253), .A2(G226), .A3(new_n254), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n266), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(G238), .B2(new_n273), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n325), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(G200), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n327), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(G190), .A3(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n320), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n329), .A2(new_n330), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(KEYINPUT72), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT14), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n339), .C1(new_n329), .C2(new_n330), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT73), .B1(new_n337), .B2(G179), .ZN(new_n344));
  AND4_X1   g0144(.A1(KEYINPUT73), .A2(new_n333), .A3(G179), .A4(new_n334), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n341), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n320), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n336), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n221), .A2(new_n217), .ZN(new_n349));
  OAI21_X1  g0149(.A(G20), .B1(new_n349), .B2(new_n201), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n291), .A2(G159), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n253), .B2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT74), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n355), .B2(KEYINPUT74), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT16), .B(new_n353), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n217), .B1(new_n355), .B2(new_n360), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n279), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n293), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n286), .B2(new_n287), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n281), .A2(new_n283), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n293), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n356), .A2(new_n358), .A3(G223), .A4(new_n254), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n356), .A2(new_n358), .A3(G226), .A4(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT75), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n263), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT75), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n263), .A2(G232), .A3(new_n270), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n272), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(G179), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n383), .B1(new_n379), .B2(new_n380), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n338), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n373), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT18), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n367), .A2(new_n372), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G200), .B2(new_n386), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n393), .A3(KEYINPUT17), .ZN(new_n394));
  AOI211_X1 g0194(.A(G190), .B(new_n383), .C1(new_n379), .C2(new_n380), .ZN(new_n395));
  AOI21_X1  g0195(.A(G200), .B1(new_n381), .B2(new_n384), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n367), .B(new_n372), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n373), .A2(new_n387), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n389), .A2(new_n394), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n253), .A2(G232), .A3(new_n254), .ZN(new_n404));
  INV_X1    g0204(.A(G107), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n405), .B2(new_n253), .C1(new_n258), .C2(new_n218), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n266), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n326), .B1(G244), .B2(new_n273), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n338), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n225), .A2(G20), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n411), .B1(new_n293), .B2(new_n292), .C1(new_n294), .C2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n279), .B1(new_n256), .B2(new_n296), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n284), .B(G77), .C1(G1), .C2(new_n210), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(KEYINPUT70), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G179), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n407), .A2(new_n418), .A3(new_n408), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT70), .B1(new_n410), .B2(new_n416), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n416), .B1(G200), .B2(new_n409), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n391), .B2(new_n409), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n311), .A2(new_n348), .A3(new_n403), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n269), .A2(G45), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(G41), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT5), .ZN(new_n434));
  AOI21_X1  g0234(.A(G41), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n438), .A2(KEYINPUT78), .A3(G41), .ZN(new_n439));
  OAI211_X1 g0239(.A(G264), .B(new_n263), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n435), .A2(new_n436), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT78), .B1(new_n438), .B2(G41), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n268), .A4(new_n431), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n356), .A2(new_n358), .A3(G250), .A4(new_n254), .ZN(new_n444));
  INV_X1    g0244(.A(G294), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n278), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n266), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n338), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n440), .A2(new_n418), .A3(new_n448), .A4(new_n443), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n269), .B2(G33), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n278), .A2(KEYINPUT76), .A3(G1), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n284), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n405), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT25), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n370), .B2(G107), .ZN(new_n459));
  AOI22_X1  g0259(.A1(G107), .A2(new_n456), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n279), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n210), .A3(G87), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n359), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n465), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n253), .A3(KEYINPUT22), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n405), .A3(G20), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT82), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n471), .A2(new_n472), .B1(KEYINPUT23), .B2(G107), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n476));
  OR2_X1    g0276(.A1(new_n476), .A2(G20), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT24), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n474), .A2(KEYINPUT82), .B1(new_n470), .B2(new_n405), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n471), .A2(new_n472), .B1(new_n476), .B2(G20), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n466), .A4(new_n468), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n462), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n450), .B(new_n451), .C1(new_n461), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n461), .A2(new_n485), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n449), .A2(G200), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(new_n391), .C2(new_n449), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n479), .A2(new_n484), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n279), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n460), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(new_n451), .A4(new_n450), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n487), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n497), .A2(new_n498), .A3(G107), .ZN(new_n499));
  XNOR2_X1  g0299(.A(G97), .B(G107), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(new_n210), .B1(new_n313), .B2(new_n292), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n405), .B1(new_n355), .B2(new_n360), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n279), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n370), .A2(G97), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n456), .B2(G97), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n356), .A2(new_n358), .A3(G250), .A4(G1698), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n356), .A2(new_n358), .A3(G244), .A4(new_n254), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n266), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(G257), .B(new_n263), .C1(new_n437), .C2(new_n439), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n443), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n507), .B1(G200), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(new_n515), .A3(new_n443), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n338), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n514), .A2(new_n515), .A3(new_n418), .A4(new_n443), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n507), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n356), .A2(new_n358), .A3(G238), .A4(new_n254), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n356), .A2(new_n358), .A3(G244), .A4(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n266), .ZN(new_n528));
  INV_X1    g0328(.A(G250), .ZN(new_n529));
  INV_X1    g0329(.A(G45), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(G1), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n269), .A2(new_n267), .A3(G45), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n263), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(G190), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n210), .ZN(new_n536));
  INV_X1    g0336(.A(G87), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n498), .A3(new_n405), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n294), .B2(new_n498), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n217), .A2(G20), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n356), .A3(new_n358), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n279), .A2(new_n544), .B1(new_n296), .B2(new_n412), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n284), .A2(G87), .A3(new_n455), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n534), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n533), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n527), .B2(new_n266), .ZN(new_n549));
  INV_X1    g0349(.A(G200), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n528), .A2(new_n418), .A3(new_n533), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n544), .A2(new_n279), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n296), .A2(new_n412), .ZN(new_n554));
  INV_X1    g0354(.A(new_n412), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n370), .A2(new_n455), .A3(new_n462), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n549), .A2(G169), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n547), .A2(new_n551), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n520), .A2(new_n523), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n496), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G270), .B(new_n263), .C1(new_n437), .C2(new_n439), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n443), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(KEYINPUT79), .A3(new_n443), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n356), .A2(new_n358), .A3(G264), .A4(G1698), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n356), .A2(new_n358), .A3(G257), .A4(new_n254), .ZN(new_n571));
  INV_X1    g0371(.A(G303), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n253), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n266), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT80), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n564), .A2(KEYINPUT79), .A3(new_n443), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT79), .B1(new_n564), .B2(new_n443), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT80), .B(new_n574), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n456), .A2(G116), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n508), .B(new_n210), .C1(G33), .C2(new_n498), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n582), .B(new_n279), .C1(new_n210), .C2(G116), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G116), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n296), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(G190), .A3(new_n578), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n580), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(G169), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n575), .B2(new_n579), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n578), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n595), .A2(new_n598), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n418), .B1(new_n573), .B2(new_n266), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n588), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n600), .A2(new_n601), .B1(new_n569), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n563), .A2(new_n594), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n428), .A2(new_n605), .ZN(G372));
  NAND2_X1  g0406(.A1(new_n308), .A2(new_n310), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n394), .A2(new_n399), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n346), .A2(new_n347), .ZN(new_n610));
  INV_X1    g0410(.A(new_n336), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n423), .A3(new_n421), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n401), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n400), .B1(new_n373), .B2(new_n387), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n607), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n302), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n428), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n521), .A2(new_n522), .A3(new_n507), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n519), .B2(new_n517), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n391), .B(new_n548), .C1(new_n527), .C2(new_n266), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n546), .A2(new_n553), .A3(new_n554), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT84), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n527), .A2(new_n628), .A3(new_n266), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n548), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n626), .B1(new_n630), .B2(new_n550), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n545), .A2(new_n556), .B1(new_n549), .B2(new_n418), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n630), .B2(G169), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n623), .A2(new_n490), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n601), .B1(new_n575), .B2(new_n579), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n603), .A2(new_n569), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n595), .B1(new_n592), .B2(new_n578), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(KEYINPUT21), .ZN(new_n640));
  INV_X1    g0440(.A(new_n486), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n635), .A2(new_n643), .A3(new_n622), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT26), .B1(new_n523), .B2(new_n560), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n633), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n620), .B1(new_n621), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT85), .ZN(G369));
  INV_X1    g0450(.A(G330), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n637), .A2(new_n638), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT21), .B1(new_n600), .B2(new_n596), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n269), .A2(new_n210), .A3(G13), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n654), .B(new_n594), .C1(new_n589), .C2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n640), .A2(new_n588), .A3(new_n660), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n651), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n641), .A2(KEYINPUT86), .A3(new_n660), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT86), .B1(new_n641), .B2(new_n660), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n488), .A2(new_n661), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n665), .A2(new_n666), .B1(new_n496), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n640), .A3(new_n661), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n641), .A2(new_n661), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n230), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n538), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n207), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n648), .A2(new_n682), .A3(new_n661), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n634), .B2(new_n523), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n622), .A2(new_n561), .A3(new_n643), .ZN(new_n685));
  AND4_X1   g0485(.A1(KEYINPUT87), .A2(new_n684), .A3(new_n633), .A4(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n633), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n523), .A2(new_n560), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n643), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT87), .B1(new_n689), .B2(new_n684), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n487), .A2(new_n495), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n636), .B1(new_n640), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n660), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n683), .B1(new_n682), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n630), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n418), .A3(new_n449), .A4(new_n516), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n575), .B2(new_n579), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n440), .A2(new_n602), .A3(new_n448), .A4(new_n549), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n516), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n569), .A2(new_n701), .A3(KEYINPUT30), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT30), .B1(new_n569), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT31), .B1(new_n705), .B2(new_n660), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n697), .B1(new_n592), .B2(new_n578), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n440), .A2(new_n448), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n602), .A2(new_n549), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n518), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n576), .A2(new_n577), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n569), .A2(new_n701), .A3(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT31), .B(new_n660), .C1(new_n707), .C2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n706), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n654), .A2(new_n594), .A3(new_n563), .A4(new_n661), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n651), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n695), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n681), .B1(new_n721), .B2(G1), .ZN(G364));
  NAND2_X1  g0522(.A1(new_n662), .A2(new_n663), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n210), .A2(G13), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n269), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n676), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n724), .A2(new_n664), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT88), .ZN(new_n731));
  INV_X1    g0531(.A(new_n729), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n253), .A2(G355), .A3(new_n230), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n251), .A2(new_n530), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n675), .A2(new_n253), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G45), .B2(new_n207), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n733), .B1(G116), .B2(new_n230), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT89), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n209), .B1(G20), .B2(new_n338), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n732), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n210), .A2(new_n391), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n418), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n210), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G58), .A2(new_n747), .B1(new_n750), .B2(new_n225), .ZN(new_n751));
  NAND3_X1  g0551(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n391), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n751), .B1(new_n202), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT90), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n550), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n405), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n744), .A2(new_n757), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n359), .B(new_n759), .C1(G87), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n210), .B1(new_n763), .B2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n498), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n752), .A2(G190), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(G68), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n748), .A2(new_n763), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n762), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n766), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n359), .B1(new_n764), .B2(new_n445), .C1(new_n572), .C2(new_n760), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n775), .B(new_n776), .C1(G326), .C2(new_n753), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n746), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n758), .B1(new_n749), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n768), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n779), .B(new_n782), .C1(G329), .C2(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n756), .A2(new_n772), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n741), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n743), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT91), .Z(new_n788));
  XOR2_X1   g0588(.A(new_n740), .B(KEYINPUT92), .Z(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n723), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n731), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  INV_X1    g0593(.A(KEYINPUT95), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n426), .B(new_n794), .C1(new_n420), .C2(new_n422), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n660), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n648), .A2(KEYINPUT96), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT96), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n599), .A2(new_n604), .A3(new_n486), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n646), .B1(new_n799), .B2(new_n636), .ZN(new_n800));
  INV_X1    g0600(.A(new_n796), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n416), .A2(new_n660), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(KEYINPUT95), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n424), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n800), .B2(new_n660), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n720), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n677), .B2(new_n727), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n803), .A2(new_n720), .A3(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G143), .A2(new_n747), .B1(new_n750), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n773), .B2(new_n290), .C1(new_n815), .C2(new_n754), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n253), .B1(new_n760), .B2(new_n202), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n758), .A2(new_n217), .B1(new_n768), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n764), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n822), .C1(G58), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n818), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n359), .B1(new_n760), .B2(new_n405), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT94), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n783), .A2(G311), .ZN(new_n828));
  INV_X1    g0628(.A(new_n758), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G294), .A2(new_n747), .B1(new_n829), .B2(G87), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n765), .B1(new_n753), .B2(G303), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n828), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n773), .A2(new_n780), .B1(new_n749), .B2(new_n586), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT93), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n825), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n741), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n741), .A2(new_n738), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n732), .B1(new_n313), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n795), .A2(new_n804), .B1(new_n424), .B2(new_n806), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n838), .C1(new_n839), .C2(new_n739), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n813), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  NAND3_X1  g0642(.A1(new_n421), .A2(new_n423), .A3(new_n661), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT97), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n797), .B2(new_n802), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  INV_X1    g0647(.A(new_n658), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n373), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n388), .A2(new_n849), .A3(new_n850), .A4(new_n397), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n363), .A2(new_n279), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT7), .B1(new_n359), .B2(new_n210), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT74), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n217), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT74), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n352), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT16), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n372), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n390), .A2(new_n393), .B1(new_n860), .B2(new_n387), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n848), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n852), .B1(KEYINPUT37), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n608), .B2(new_n616), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n847), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n850), .B1(new_n861), .B2(new_n862), .ZN(new_n867));
  OAI221_X1 g0667(.A(KEYINPUT38), .B1(new_n867), .B2(new_n852), .C1(new_n403), .C2(new_n862), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n347), .B(new_n660), .C1(new_n346), .C2(new_n336), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n320), .A2(new_n661), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n336), .B(new_n873), .C1(new_n346), .C2(new_n347), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n846), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n851), .A2(KEYINPUT98), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n388), .A2(new_n849), .A3(new_n397), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n851), .A2(KEYINPUT98), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n402), .A2(new_n373), .A3(new_n848), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n864), .A2(new_n865), .A3(new_n847), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n346), .A2(new_n347), .A3(new_n661), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n866), .A2(new_n868), .A3(KEYINPUT39), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n616), .A2(new_n848), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n876), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n620), .B1(new_n695), .B2(new_n621), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT99), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT40), .B1(new_n884), .B2(new_n885), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n705), .A2(new_n660), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT31), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n716), .C1(new_n605), .C2(new_n660), .ZN(new_n902));
  INV_X1    g0702(.A(new_n874), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n808), .B1(new_n903), .B2(new_n871), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n897), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n881), .A2(new_n880), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n851), .A2(KEYINPUT98), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n883), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n847), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(new_n868), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n839), .B1(new_n872), .B2(new_n874), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n719), .B2(new_n718), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT99), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n869), .A2(new_n902), .A3(new_n904), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n906), .A2(new_n915), .B1(new_n907), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n428), .B1(new_n719), .B2(new_n718), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n651), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n896), .A2(new_n920), .B1(G1), .B2(new_n725), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n896), .B2(new_n920), .ZN(new_n922));
  INV_X1    g0722(.A(new_n501), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n924), .A2(G116), .A3(new_n211), .A4(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT36), .Z(new_n927));
  OAI211_X1 g0727(.A(new_n208), .B(new_n225), .C1(new_n221), .C2(new_n217), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n269), .B(G13), .C1(new_n928), .C2(new_n247), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(new_n930), .ZN(G367));
  OAI21_X1  g0731(.A(new_n742), .B1(new_n230), .B2(new_n412), .ZN(new_n932));
  INV_X1    g0732(.A(new_n735), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n241), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n729), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT102), .B1(new_n761), .B2(G116), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT46), .ZN(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n746), .A2(new_n572), .B1(new_n768), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G283), .B2(new_n750), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n359), .B1(new_n758), .B2(new_n498), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(G311), .B2(new_n753), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n823), .A2(G107), .B1(G294), .B2(new_n766), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n937), .A2(new_n940), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT103), .B(G137), .Z(new_n945));
  OAI22_X1  g0745(.A1(new_n945), .A2(new_n768), .B1(new_n760), .B2(new_n221), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT104), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n359), .B1(new_n829), .B2(new_n225), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G150), .A2(new_n747), .B1(new_n750), .B2(G50), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n823), .A2(G68), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n753), .A2(G143), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(new_n769), .C2(new_n773), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n944), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n935), .B1(new_n957), .B2(new_n741), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n625), .A2(new_n660), .ZN(new_n959));
  MUX2_X1   g0759(.A(new_n633), .B(new_n634), .S(new_n959), .Z(new_n960));
  INV_X1    g0760(.A(new_n789), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT101), .ZN(new_n964));
  INV_X1    g0764(.A(new_n721), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n507), .A2(new_n660), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n623), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n622), .A2(new_n660), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n673), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n672), .A2(KEYINPUT44), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n672), .B2(new_n972), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n669), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n669), .B1(new_n974), .B2(new_n978), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n654), .A2(new_n660), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n668), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n670), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n664), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n965), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n676), .B(KEYINPUT41), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n964), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n974), .A2(new_n978), .ZN(new_n990));
  INV_X1    g0790(.A(new_n669), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n992), .A2(new_n721), .A3(new_n986), .A4(new_n979), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n721), .ZN(new_n994));
  INV_X1    g0794(.A(new_n988), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(KEYINPUT101), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n728), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n670), .A2(new_n972), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT42), .Z(new_n999));
  INV_X1    g0799(.A(new_n692), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n523), .B1(new_n968), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n661), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n960), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  MUX2_X1   g0805(.A(KEYINPUT43), .B(new_n1003), .S(new_n960), .Z(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n669), .B2(new_n972), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n669), .A2(new_n972), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1005), .B(new_n1009), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n963), .B1(new_n997), .B2(new_n1011), .ZN(G387));
  OR2_X1    g0812(.A1(new_n668), .A2(new_n789), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n678), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1014), .A2(new_n230), .A3(new_n253), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(G107), .B2(new_n230), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n238), .A2(new_n530), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n1014), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n293), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n933), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1016), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n742), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n729), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n764), .A2(new_n412), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n359), .B(new_n1025), .C1(G97), .C2(new_n829), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G68), .A2(new_n750), .B1(new_n783), .B2(G150), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n225), .A2(new_n761), .B1(new_n747), .B2(G50), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n368), .A2(new_n766), .B1(G159), .B2(new_n753), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n253), .B1(new_n783), .B2(G326), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n760), .A2(new_n445), .B1(new_n764), .B2(new_n780), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G317), .A2(new_n747), .B1(new_n750), .B2(G303), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n773), .B2(new_n781), .C1(new_n778), .C2(new_n754), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT49), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1031), .B1(new_n586), .B2(new_n758), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1030), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1024), .B1(new_n1041), .B2(new_n741), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT105), .Z(new_n1043));
  AOI22_X1  g0843(.A1(new_n986), .A2(new_n728), .B1(new_n1013), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n986), .A2(new_n721), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n676), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n986), .A2(new_n721), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n980), .B2(new_n981), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n993), .A3(new_n676), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n972), .A2(new_n740), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n245), .A2(new_n933), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n742), .B1(new_n498), .B2(new_n230), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n729), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n747), .A2(G311), .B1(G317), .B2(new_n753), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT52), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n760), .A2(new_n780), .B1(new_n768), .B2(new_n778), .ZN(new_n1057));
  OR4_X1    g0857(.A1(new_n253), .A2(new_n1056), .A3(new_n759), .A4(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n749), .A2(new_n445), .B1(new_n764), .B2(new_n586), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G303), .B2(new_n766), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT108), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G68), .A2(new_n761), .B1(new_n783), .B2(G143), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n253), .C1(new_n537), .C2(new_n758), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT106), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n754), .A2(new_n290), .B1(new_n746), .B2(new_n769), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n750), .A2(new_n368), .B1(G50), .B2(new_n766), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT107), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT107), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n313), .C2(new_n764), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1058), .A2(new_n1061), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1054), .B1(new_n1072), .B2(new_n741), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n982), .A2(new_n728), .B1(new_n1051), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1050), .A2(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(new_n875), .ZN(new_n1076));
  AND4_X1   g0876(.A1(G330), .A2(new_n902), .A3(new_n839), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n887), .B1(new_n884), .B2(new_n885), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n691), .A2(new_n693), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n661), .A3(new_n839), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n844), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1081), .B2(new_n1076), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n887), .B1(new_n846), .B2(new_n875), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n886), .A2(new_n889), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1077), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n720), .A2(new_n839), .A3(new_n1076), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1082), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n728), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n837), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n729), .B1(new_n368), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT111), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n359), .B1(new_n760), .B2(new_n537), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT113), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G116), .A2(new_n747), .B1(new_n829), .B2(G68), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G97), .A2(new_n750), .B1(new_n783), .B2(G294), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n773), .A2(new_n405), .B1(new_n764), .B2(new_n313), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G283), .B2(new_n753), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n253), .B1(new_n758), .B2(new_n202), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT112), .Z(new_n1103));
  NOR2_X1   g0903(.A1(new_n760), .A2(new_n290), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  INV_X1    g0906(.A(G125), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n749), .A2(new_n1106), .B1(new_n768), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G132), .B2(new_n747), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1103), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n823), .A2(G159), .B1(G128), .B2(new_n753), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n773), .B2(new_n945), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1101), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1094), .B1(new_n1113), .B2(new_n741), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1084), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n739), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1091), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT96), .B1(new_n648), .B2(new_n796), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n800), .A2(new_n798), .A3(new_n801), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n844), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n888), .B1(new_n1120), .B2(new_n1076), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1088), .B1(new_n1121), .B2(new_n1115), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1077), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n621), .A2(new_n720), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT109), .B1(new_n895), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n682), .B1(new_n1079), .B2(new_n661), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n800), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n621), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n620), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1128), .A2(KEYINPUT109), .A3(new_n1129), .A4(new_n1124), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1125), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1087), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1076), .B1(new_n720), .B2(new_n839), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1120), .B1(new_n1077), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n902), .A2(G330), .A3(new_n839), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n875), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1137), .A2(new_n844), .A3(new_n1086), .A4(new_n1080), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1123), .A2(new_n1132), .A3(new_n1133), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT110), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1128), .A2(new_n1129), .A3(new_n1124), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT109), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1139), .A2(new_n1145), .A3(new_n1130), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(new_n1123), .A3(KEYINPUT110), .A4(new_n1133), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1146), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1123), .A2(new_n1133), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n677), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1117), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(G378));
  AOI21_X1  g0953(.A(KEYINPUT110), .B1(new_n1090), .B2(new_n1146), .ZN(new_n1154));
  AND4_X1   g0954(.A1(KEYINPUT110), .A2(new_n1146), .A3(new_n1123), .A4(new_n1133), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1132), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n651), .B1(new_n916), .B2(new_n907), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n898), .A2(new_n905), .A3(new_n897), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT99), .B1(new_n912), .B2(new_n914), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n893), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1120), .A2(new_n869), .A3(new_n1076), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n906), .A2(new_n915), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n1158), .C1(new_n876), .C2(new_n893), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n607), .A2(new_n619), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n299), .A2(new_n658), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n311), .B1(new_n299), .B2(new_n658), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT116), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1167), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1175), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1164), .A2(new_n1177), .A3(new_n1166), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1157), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n677), .B1(new_n1156), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1145), .A2(new_n1130), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT117), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1164), .A2(new_n1177), .A3(new_n1166), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1177), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1176), .A2(KEYINPUT117), .A3(new_n1178), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1157), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1180), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n728), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n739), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1174), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n732), .B1(new_n202), .B2(new_n837), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n773), .A2(new_n821), .B1(new_n764), .B2(new_n290), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n747), .A2(G128), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n815), .B2(new_n749), .C1(new_n760), .C2(new_n1106), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G125), .C2(new_n753), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n829), .C2(G159), .ZN(new_n1202));
  INV_X1    g1002(.A(G124), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n768), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT115), .Z(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G107), .A2(new_n747), .B1(new_n783), .B2(G283), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n412), .B2(new_n749), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n758), .A2(new_n221), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT114), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n761), .A2(new_n225), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G97), .A2(new_n766), .B1(new_n753), .B2(G116), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n253), .A2(G41), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n953), .A4(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1208), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT58), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1213), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1215), .A2(KEYINPUT58), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n1206), .A2(new_n1216), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1193), .B(new_n1194), .C1(new_n786), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1191), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1190), .A2(new_n1223), .ZN(G375));
  INV_X1    g1024(.A(KEYINPUT118), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1139), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1181), .A2(new_n1227), .A3(KEYINPUT118), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n1149), .A3(new_n995), .A4(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n729), .B1(G68), .B2(new_n1092), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n253), .B(new_n1025), .C1(G303), .C2(new_n783), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G77), .A2(new_n829), .B1(new_n750), .B2(G107), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n761), .B1(new_n747), .B2(G283), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G116), .A2(new_n766), .B1(new_n753), .B2(G294), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n253), .B1(new_n749), .B2(new_n290), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1236), .B(new_n1210), .C1(G50), .C2(new_n823), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n753), .A2(G132), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n945), .B2(new_n746), .C1(new_n773), .C2(new_n1106), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT119), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G159), .A2(new_n761), .B1(new_n783), .B2(G128), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT120), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1237), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1239), .A2(KEYINPUT119), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1235), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1230), .B1(new_n1245), .B2(new_n741), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n738), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1076), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1227), .B2(new_n727), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1229), .A2(new_n1250), .ZN(G381));
  INV_X1    g1051(.A(G375), .ZN(new_n1252));
  INV_X1    g1052(.A(G387), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n792), .B(new_n1044), .C1(new_n1047), .C2(new_n1046), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(G381), .A2(G384), .A3(G390), .A4(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1152), .A4(new_n1255), .ZN(G407));
  NAND2_X1  g1056(.A1(new_n659), .A2(G213), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1252), .A2(new_n1152), .A3(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(G407), .A2(G213), .A3(new_n1259), .ZN(G409));
  NAND2_X1  g1060(.A1(G396), .A2(G393), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1254), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(G390), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT101), .B1(new_n994), .B2(new_n995), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n964), .B(new_n988), .C1(new_n993), .C2(new_n721), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n727), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1011), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1265), .B1(new_n1270), .B2(new_n963), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n963), .ZN(new_n1272));
  AOI211_X1 g1072(.A(KEYINPUT124), .B(new_n1272), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1264), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(KEYINPUT124), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1270), .A2(new_n1265), .A3(new_n963), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1263), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1226), .B(new_n1228), .C1(new_n1280), .C2(new_n1146), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n677), .B1(new_n1282), .B2(KEYINPUT60), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1250), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n841), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(G384), .A3(new_n1250), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1152), .B(new_n1222), .C1(new_n1180), .C2(new_n1189), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1188), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1156), .A3(new_n995), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n728), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1221), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G378), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1290), .B(new_n1257), .C1(new_n1291), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1279), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT121), .B1(new_n1291), .B2(new_n1297), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G384), .B1(new_n1284), .B2(new_n1250), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n841), .B(new_n1249), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT57), .B1(new_n1292), .B2(new_n1156), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1179), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n676), .B1(new_n1182), .B2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G378), .B(new_n1223), .C1(new_n1304), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT121), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1182), .A2(new_n1188), .A3(new_n988), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1152), .B1(new_n1309), .B2(new_n1295), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1300), .A2(new_n1257), .A3(new_n1303), .A4(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1299), .B1(new_n1312), .B2(new_n1289), .ZN(new_n1313));
  INV_X1    g1113(.A(G2897), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1257), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT122), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1286), .A2(new_n1316), .A3(new_n1287), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT122), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1315), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1315), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1303), .B2(new_n1316), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1311), .A2(new_n1257), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1308), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1324));
  OAI211_X1 g1124(.A(KEYINPUT123), .B(new_n1322), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1300), .A2(new_n1257), .A3(new_n1311), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT123), .B1(new_n1327), .B2(new_n1322), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1313), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  OR2_X1    g1129(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1258), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1275), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1288), .A2(new_n1333), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1331), .A2(KEYINPUT125), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT125), .B1(new_n1331), .B2(new_n1334), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1312), .A2(new_n1333), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1332), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1329), .B1(new_n1339), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT126), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1329), .B(KEYINPUT126), .C1(new_n1339), .C2(new_n1341), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1152), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1307), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1288), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1341), .ZN(G402));
endmodule


