//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n472), .B2(G137), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n473), .B1(new_n478), .B2(KEYINPUT66), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n480), .B(new_n464), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT67), .Z(G160));
  NAND2_X1  g058(.A1(new_n472), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n474), .B2(new_n475), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT68), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n493), .A2(KEYINPUT68), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n498), .A2(new_n500), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT69), .A3(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT69), .A2(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR3_X1    g089(.A1(new_n514), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n516), .A2(KEYINPUT71), .A3(G50), .A4(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(G543), .A3(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XOR2_X1   g099(.A(new_n524), .B(KEYINPUT72), .Z(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n523), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n530), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n513), .A2(G88), .A3(new_n515), .A4(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(G166));
  AND2_X1   g112(.A1(new_n516), .A2(new_n533), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  INV_X1    g114(.A(new_n519), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n544));
  AND2_X1   g119(.A1(G63), .A2(G651), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n533), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n539), .A2(new_n541), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  NAND2_X1  g123(.A1(new_n538), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n540), .A2(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(new_n533), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(new_n523), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n549), .A2(new_n550), .A3(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND2_X1  g132(.A1(new_n540), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(new_n523), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n516), .A2(new_n533), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n558), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g145(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n571));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(new_n538), .A2(G91), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n519), .A2(KEYINPUT9), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n519), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n530), .ZN(new_n580));
  NOR2_X1   g155(.A1(KEYINPUT5), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT75), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n529), .A2(new_n583), .A3(new_n530), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G65), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT76), .B1(new_n588), .B2(G651), .ZN(new_n589));
  INV_X1    g164(.A(G65), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n582), .B2(new_n584), .ZN(new_n591));
  INV_X1    g166(.A(new_n587), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT76), .B(G651), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n575), .B(new_n579), .C1(new_n589), .C2(new_n594), .ZN(G299));
  NAND3_X1  g170(.A1(new_n522), .A2(new_n535), .A3(KEYINPUT77), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n522), .B2(new_n535), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(G303));
  NAND4_X1  g174(.A1(new_n513), .A2(G87), .A3(new_n515), .A4(new_n533), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n601));
  INV_X1    g176(.A(G49), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n600), .B(new_n601), .C1(new_n519), .C2(new_n602), .ZN(G288));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n529), .B2(new_n530), .ZN(new_n605));
  AND2_X1   g180(.A1(G73), .A2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n523), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n513), .A2(G86), .A3(new_n515), .A4(new_n533), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n513), .A2(G48), .A3(G543), .A4(new_n515), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(G305));
  AOI22_X1  g185(.A1(new_n538), .A2(G85), .B1(G47), .B2(new_n540), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n552), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n523), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n616), .B2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT79), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n538), .A2(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n585), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(new_n514), .ZN(new_n626));
  INV_X1    g201(.A(G54), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n519), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n519), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n621), .B1(new_n632), .B2(G868), .ZN(G284));
  OAI21_X1  g208(.A(new_n621), .B1(new_n632), .B2(G868), .ZN(G321));
  NAND2_X1  g209(.A1(G286), .A2(G868), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G297));
  OAI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n632), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n485), .A2(G123), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT81), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  INV_X1    g222(.A(G111), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(G2105), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(G135), .B2(new_n472), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT12), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  INV_X1    g230(.A(G2100), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(G2096), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n652), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2430), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(KEYINPUT14), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XOR2_X1   g244(.A(G1341), .B(G1348), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2443), .B(G2446), .Z(new_n673));
  OAI21_X1  g248(.A(G14), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT83), .ZN(G401));
  XNOR2_X1  g251(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n677), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n656), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT84), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n677), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2096), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n685), .B(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1971), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT20), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n692), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n692), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G4), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n632), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G1348), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G32), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n472), .A2(G141), .ZN(new_n715));
  INV_X1    g290(.A(G105), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n465), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n485), .A2(G129), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(new_n713), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT27), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1996), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT25), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n472), .A2(G139), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(new_n464), .C2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G33), .B(new_n731), .S(G29), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n713), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n472), .A2(G140), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n485), .A2(G128), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n736), .B1(new_n713), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2067), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT29), .B(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n733), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n713), .A2(G27), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G164), .B2(new_n713), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2078), .ZN(new_n751));
  NOR2_X1   g326(.A1(G171), .A2(new_n708), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G5), .B2(new_n708), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND4_X1   g330(.A1(new_n712), .A2(new_n726), .A3(new_n748), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n708), .A2(G21), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G168), .B2(new_n708), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n753), .A2(new_n754), .B1(G1966), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G1966), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n646), .A2(G29), .A3(new_n650), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT93), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT93), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT30), .B(G28), .ZN(new_n764));
  OR2_X1    g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  NAND2_X1  g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n764), .A2(new_n713), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n708), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n636), .B2(new_n708), .ZN(new_n773));
  INV_X1    g348(.A(G1956), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n708), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n568), .B2(new_n708), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  NAND2_X1  g353(.A1(G160), .A2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(G34), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G34), .B2(new_n780), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT92), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n756), .A2(new_n770), .A3(new_n775), .A4(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G6), .B(G305), .S(G16), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G23), .B(G288), .S(G16), .Z(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n708), .A2(G22), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n536), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n791), .B(new_n794), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT89), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT89), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n802), .A2(KEYINPUT34), .A3(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G24), .B(G290), .S(G16), .Z(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(G1986), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(G1986), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n713), .A2(G25), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G107), .B2(new_n464), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT87), .ZN(new_n812));
  AOI22_X1  g387(.A1(G119), .A2(new_n485), .B1(new_n472), .B2(G131), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n713), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  NOR3_X1   g392(.A1(new_n806), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n804), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT34), .B1(new_n802), .B2(new_n803), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT36), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n820), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n822), .A2(new_n823), .A3(new_n804), .A4(new_n818), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n788), .B1(new_n821), .B2(new_n824), .ZN(G311));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n826));
  XNOR2_X1  g401(.A(G311), .B(new_n826), .ZN(G150));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n552), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n538), .A2(G93), .B1(new_n523), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT96), .B(G55), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n519), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n567), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n565), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT38), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n631), .A2(new_n639), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  AOI21_X1  g415(.A(G860), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(KEYINPUT100), .B(G37), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n472), .A2(G142), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n485), .A2(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n464), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT97), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n654), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n814), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT98), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n508), .B(new_n741), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n731), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n722), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G160), .B(new_n489), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n651), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n855), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n847), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n859), .B2(new_n856), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n856), .A2(KEYINPUT99), .A3(new_n859), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g448(.A(KEYINPUT40), .B(new_n868), .C1(new_n873), .C2(new_n862), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n862), .B1(new_n871), .B2(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(new_n868), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n874), .A2(new_n878), .ZN(G395));
  XNOR2_X1  g454(.A(G290), .B(G288), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n536), .B(G305), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(KEYINPUT42), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT103), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n631), .B(new_n636), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n641), .B(new_n836), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n889), .B(new_n896), .ZN(new_n897));
  MUX2_X1   g472(.A(new_n833), .B(new_n897), .S(G868), .Z(G295));
  MUX2_X1   g473(.A(new_n833), .B(new_n897), .S(G868), .Z(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  XNOR2_X1  g475(.A(G301), .B(G286), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n836), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n891), .A2(new_n902), .A3(new_n892), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n836), .B(new_n901), .Z(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n890), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n905), .A3(new_n884), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n884), .B1(new_n903), .B2(new_n905), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n847), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n903), .A2(new_n905), .ZN(new_n913));
  INV_X1    g488(.A(new_n884), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT104), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n909), .B2(G37), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n912), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n900), .B(new_n911), .C1(new_n920), .C2(new_n907), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n908), .B1(new_n917), .B2(new_n919), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n909), .A2(new_n847), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n907), .B1(new_n923), .B2(new_n906), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT44), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n921), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT4), .B1(new_n493), .B2(KEYINPUT68), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n496), .B1(new_n495), .B2(new_n492), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n477), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n495), .B2(G125), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n480), .B1(new_n936), .B2(new_n464), .ZN(new_n937));
  INV_X1    g512(.A(G125), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n470), .B2(new_n471), .ZN(new_n939));
  OAI211_X1 g514(.A(KEYINPUT66), .B(G2105), .C1(new_n939), .C2(new_n935), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n937), .A2(G40), .A3(new_n940), .A4(new_n473), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n741), .B(G2067), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT106), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n944), .B2(new_n722), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n934), .A2(G1996), .A3(new_n941), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT105), .Z(new_n947));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  AND3_X1   g527(.A1(new_n942), .A2(G1996), .A3(new_n722), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n942), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT107), .Z(new_n955));
  AOI211_X1 g530(.A(new_n953), .B(new_n955), .C1(new_n723), .C2(new_n947), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n814), .B(new_n816), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n942), .ZN(new_n958));
  NOR2_X1   g533(.A1(G290), .A2(G1986), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n942), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT48), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n956), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n814), .A2(new_n816), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT127), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n952), .B(new_n962), .C1(new_n942), .C2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n479), .A2(new_n971), .A3(new_n481), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n934), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT108), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n934), .A2(new_n975), .A3(new_n970), .A4(new_n972), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n797), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n506), .B1(new_n499), .B2(new_n929), .ZN(new_n978));
  AOI211_X1 g553(.A(KEYINPUT50), .B(G1384), .C1(new_n978), .C2(new_n498), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n508), .B2(new_n927), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n979), .A2(new_n981), .A3(new_n941), .ZN(new_n982));
  INV_X1    g557(.A(G2090), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT77), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n536), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n988));
  NOR2_X1   g563(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n987), .A2(G8), .A3(new_n596), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n597), .A2(new_n993), .A3(new_n598), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n994), .B2(new_n988), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n985), .A2(G8), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  NAND2_X1  g572(.A1(G305), .A2(KEYINPUT49), .ZN(new_n998));
  INV_X1    g573(.A(G1981), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n607), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n608), .A2(new_n607), .A3(new_n609), .A4(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n998), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n998), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n978), .B2(new_n498), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n972), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1009), .B2(G8), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(G8), .C1(new_n932), .C2(new_n941), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n997), .B(new_n1006), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n932), .B2(new_n941), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1011), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n997), .B1(new_n1017), .B2(new_n1006), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G288), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(new_n1023), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1019), .A2(KEYINPUT113), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1006), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1013), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1025), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1023), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1021), .B(new_n1034), .C1(new_n1016), .C2(new_n1011), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1029), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n996), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g613(.A(G1976), .B(G288), .C1(new_n1031), .C2(new_n1013), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1017), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G2078), .B1(new_n974), .B2(new_n976), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(KEYINPUT53), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n972), .B1(new_n1008), .B2(new_n980), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n979), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n941), .B1(new_n932), .B2(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1008), .A2(new_n980), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(KEYINPUT116), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n754), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2078), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT53), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n973), .A2(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1051), .A2(KEYINPUT120), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT120), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1044), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT121), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1060), .A3(G171), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT114), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1032), .A2(new_n1036), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n985), .A2(new_n995), .A3(G8), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n985), .A2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(new_n995), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n993), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n973), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1048), .A2(new_n785), .A3(new_n1049), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G168), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(G286), .A3(new_n1077), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(G168), .A3(new_n1077), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT51), .B1(new_n1082), .B2(G8), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1071), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1076), .A2(G286), .A3(new_n1077), .ZN(new_n1085));
  AOI21_X1  g660(.A(G286), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1073), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1082), .A2(G8), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1087), .B(KEYINPUT62), .C1(KEYINPUT51), .C2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1070), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1042), .B1(new_n1062), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1079), .A2(new_n993), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1070), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n995), .B1(new_n985), .B2(G8), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n996), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1095), .A2(new_n1093), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1098), .B(new_n1099), .C1(new_n1037), .C2(new_n1028), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1057), .A2(new_n1060), .A3(G171), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1060), .B1(new_n1057), .B2(G171), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n473), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1105), .A2(KEYINPUT122), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(KEYINPUT122), .ZN(new_n1107));
  NOR4_X1   g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n971), .A4(new_n1053), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(G2105), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1108), .A2(new_n934), .A3(new_n970), .A4(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1051), .B(new_n1112), .C1(new_n1043), .C2(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT124), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT54), .B1(new_n1104), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n934), .A2(new_n970), .A3(new_n972), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1956), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT115), .B(new_n575), .C1(new_n589), .C2(new_n594), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n1123));
  NAND3_X1  g698(.A1(G299), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT76), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n591), .A2(new_n592), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n514), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1127), .A2(new_n593), .B1(G91), .B2(new_n538), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n579), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1121), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1047), .A2(new_n711), .A3(new_n1050), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n972), .A2(new_n1008), .A3(new_n966), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n631), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1124), .B(new_n1129), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1131), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT117), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(new_n1131), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1009), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n973), .B2(G1996), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n568), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT59), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n568), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n631), .A4(new_n1133), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1118), .B1(new_n982), .B2(G1956), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1130), .B(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1135), .B2(KEYINPUT119), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1149), .B(new_n1150), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1131), .A2(new_n1156), .A3(new_n1135), .A4(KEYINPUT61), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT60), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n1133), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n632), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1138), .B(new_n1140), .C1(new_n1155), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1070), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1044), .B(G301), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1113), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT125), .B1(new_n1113), .B2(G171), .ZN(new_n1167));
  OAI211_X1 g742(.A(KEYINPUT54), .B(new_n1164), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1162), .A2(new_n1163), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1092), .B(new_n1101), .C1(new_n1116), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n956), .A2(new_n958), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G290), .B(G1986), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n942), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1171), .A2(KEYINPUT126), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT126), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n969), .B1(new_n1175), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g752(.A1(G229), .A2(new_n462), .A3(new_n675), .A4(G227), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n876), .B2(new_n877), .ZN(new_n1180));
  OR2_X1    g754(.A1(new_n920), .A2(new_n907), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1181), .B2(new_n911), .ZN(G308));
  OAI21_X1  g756(.A(new_n868), .B1(new_n873), .B2(new_n862), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n920), .A2(new_n907), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n1183), .B(new_n1179), .C1(new_n1184), .C2(new_n910), .ZN(G225));
endmodule


