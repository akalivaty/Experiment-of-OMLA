

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799;

  AND2_X1 U377 ( .A1(n761), .A2(n718), .ZN(n390) );
  INV_X1 U378 ( .A(n770), .ZN(n355) );
  XNOR2_X1 U379 ( .A(n655), .B(KEYINPUT78), .ZN(n668) );
  AND2_X1 U380 ( .A1(n722), .A2(n588), .ZN(n589) );
  OR2_X1 U381 ( .A1(n741), .A2(n621), .ZN(n641) );
  AND2_X1 U382 ( .A1(n401), .A2(n400), .ZN(n370) );
  XNOR2_X1 U383 ( .A(n433), .B(n771), .ZN(n659) );
  XNOR2_X1 U384 ( .A(n415), .B(n414), .ZN(n425) );
  NOR2_X1 U385 ( .A1(G953), .A2(G237), .ZN(n535) );
  XNOR2_X1 U386 ( .A(n472), .B(KEYINPUT74), .ZN(n505) );
  INV_X1 U387 ( .A(G110), .ZN(n472) );
  INV_X1 U388 ( .A(n354), .ZN(n664) );
  NAND2_X1 U389 ( .A1(n356), .A2(n355), .ZN(n354) );
  XNOR2_X1 U390 ( .A(n661), .B(n357), .ZN(n356) );
  INV_X1 U391 ( .A(n660), .ZN(n357) );
  XNOR2_X2 U392 ( .A(n358), .B(n553), .ZN(n560) );
  NAND2_X2 U393 ( .A1(n581), .A2(n411), .ZN(n358) );
  INV_X1 U394 ( .A(G953), .ZN(n786) );
  AND2_X2 U395 ( .A1(n784), .A2(n421), .ZN(n420) );
  AND2_X2 U396 ( .A1(n423), .A2(n420), .ZN(n387) );
  AND2_X2 U397 ( .A1(n431), .A2(n428), .ZN(n427) );
  OR2_X2 U398 ( .A1(n378), .A2(n602), .ZN(n635) );
  NOR2_X2 U399 ( .A1(n408), .A2(n403), .ZN(n402) );
  AND2_X2 U400 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X2 U401 ( .A1(n578), .A2(n577), .ZN(n579) );
  BUF_X1 U402 ( .A(n744), .Z(n359) );
  INV_X1 U403 ( .A(G140), .ZN(n414) );
  NOR2_X1 U404 ( .A1(n635), .A2(n645), .ZN(n636) );
  XNOR2_X1 U405 ( .A(KEYINPUT105), .B(n584), .ZN(n744) );
  XNOR2_X1 U406 ( .A(n549), .B(G478), .ZN(n585) );
  XNOR2_X1 U407 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(G902), .ZN(n648) );
  NAND2_X2 U409 ( .A1(n370), .A2(n446), .ZN(n413) );
  NAND2_X2 U410 ( .A1(n447), .A2(n517), .ZN(n446) );
  XNOR2_X2 U411 ( .A(n547), .B(n470), .ZN(n783) );
  XNOR2_X2 U412 ( .A(n532), .B(n450), .ZN(n782) );
  XOR2_X1 U413 ( .A(G137), .B(KEYINPUT71), .Z(n478) );
  NAND2_X1 U414 ( .A1(n594), .A2(n515), .ZN(n409) );
  NAND2_X1 U415 ( .A1(n407), .A2(n648), .ZN(n406) );
  INV_X1 U416 ( .A(n515), .ZN(n407) );
  INV_X1 U417 ( .A(G902), .ZN(n514) );
  INV_X1 U418 ( .A(KEYINPUT69), .ZN(n382) );
  XNOR2_X1 U419 ( .A(G131), .B(KEYINPUT4), .ZN(n470) );
  XNOR2_X1 U420 ( .A(G119), .B(G128), .ZN(n454) );
  XOR2_X1 U421 ( .A(KEYINPUT23), .B(KEYINPUT73), .Z(n455) );
  XOR2_X1 U422 ( .A(KEYINPUT79), .B(KEYINPUT96), .Z(n452) );
  XNOR2_X1 U423 ( .A(n783), .B(G146), .ZN(n496) );
  NAND2_X1 U424 ( .A1(n585), .A2(n412), .ZN(n673) );
  INV_X1 U425 ( .A(KEYINPUT39), .ZN(n432) );
  XNOR2_X1 U426 ( .A(G113), .B(G131), .ZN(n530) );
  XNOR2_X1 U427 ( .A(G143), .B(G128), .ZN(n371) );
  XOR2_X1 U428 ( .A(KEYINPUT91), .B(KEYINPUT18), .Z(n511) );
  INV_X1 U429 ( .A(KEYINPUT35), .ZN(n417) );
  INV_X1 U430 ( .A(n670), .ZN(n445) );
  AND2_X1 U431 ( .A1(n670), .A2(KEYINPUT19), .ZN(n443) );
  XNOR2_X1 U432 ( .A(n435), .B(n502), .ZN(n771) );
  XNOR2_X1 U433 ( .A(G107), .B(KEYINPUT95), .ZN(n473) );
  INV_X1 U434 ( .A(KEYINPUT83), .ZN(n422) );
  NAND2_X1 U435 ( .A1(n648), .A2(n422), .ZN(n421) );
  INV_X1 U436 ( .A(G237), .ZN(n513) );
  XOR2_X1 U437 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n486) );
  INV_X1 U438 ( .A(KEYINPUT77), .ZN(n487) );
  XNOR2_X1 U439 ( .A(G116), .B(G137), .ZN(n488) );
  XNOR2_X1 U440 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n499) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n518) );
  NAND2_X1 U442 ( .A1(n404), .A2(n443), .ZN(n400) );
  XNOR2_X1 U443 ( .A(n497), .B(G472), .ZN(n689) );
  NOR2_X1 U444 ( .A1(n673), .A2(n683), .ZN(n411) );
  XNOR2_X1 U445 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U446 ( .A(G122), .B(KEYINPUT103), .ZN(n538) );
  XNOR2_X1 U447 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n540) );
  XOR2_X1 U448 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n541) );
  INV_X1 U449 ( .A(G101), .ZN(n471) );
  OR2_X1 U450 ( .A1(n430), .A2(KEYINPUT39), .ZN(n428) );
  NOR2_X1 U451 ( .A1(n602), .A2(n613), .ZN(n430) );
  OR2_X1 U452 ( .A1(n613), .A2(n432), .ZN(n429) );
  INV_X1 U453 ( .A(n585), .ZN(n552) );
  XNOR2_X1 U454 ( .A(n533), .B(n389), .ZN(n758) );
  XNOR2_X1 U455 ( .A(n534), .B(n360), .ZN(n389) );
  INV_X1 U456 ( .A(KEYINPUT36), .ZN(n372) );
  NOR2_X1 U457 ( .A1(n641), .A2(n645), .ZN(n623) );
  NAND2_X1 U458 ( .A1(n369), .A2(n443), .ZN(n442) );
  INV_X1 U459 ( .A(n606), .ZN(n436) );
  INV_X1 U460 ( .A(KEYINPUT66), .ZN(n438) );
  NAND2_X1 U461 ( .A1(n586), .A2(n585), .ZN(n741) );
  AND2_X1 U462 ( .A1(n709), .A2(n786), .ZN(n710) );
  XNOR2_X1 U463 ( .A(n708), .B(KEYINPUT121), .ZN(n709) );
  AND2_X1 U464 ( .A1(G214), .A2(n535), .ZN(n360) );
  AND2_X1 U465 ( .A1(n639), .A2(n734), .ZN(n361) );
  OR2_X1 U466 ( .A1(n602), .A2(n429), .ZN(n362) );
  AND2_X1 U467 ( .A1(n442), .A2(n444), .ZN(n363) );
  OR2_X1 U468 ( .A1(n525), .A2(n441), .ZN(n364) );
  XNOR2_X1 U469 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n365) );
  XOR2_X1 U470 ( .A(n593), .B(KEYINPUT45), .Z(n366) );
  AND2_X1 U471 ( .A1(n594), .A2(KEYINPUT83), .ZN(n367) );
  BUF_X1 U472 ( .A(n611), .Z(n368) );
  INV_X1 U473 ( .A(n447), .ZN(n369) );
  NAND2_X1 U474 ( .A1(n408), .A2(n405), .ZN(n622) );
  XNOR2_X1 U475 ( .A(n623), .B(n372), .ZN(n624) );
  BUF_X1 U476 ( .A(n555), .Z(n686) );
  XNOR2_X1 U477 ( .A(n611), .B(n484), .ZN(n555) );
  XNOR2_X1 U478 ( .A(n384), .B(n482), .ZN(n611) );
  BUF_X1 U479 ( .A(n711), .Z(n373) );
  BUF_X1 U480 ( .A(n685), .Z(n374) );
  BUF_X1 U481 ( .A(n766), .Z(n375) );
  BUF_X1 U482 ( .A(n798), .Z(n376) );
  AND2_X2 U483 ( .A1(n560), .A2(n619), .ZN(n571) );
  NAND2_X1 U484 ( .A1(n394), .A2(n573), .ZN(n722) );
  XNOR2_X1 U485 ( .A(n395), .B(KEYINPUT87), .ZN(n394) );
  BUF_X1 U486 ( .A(n380), .Z(n377) );
  XNOR2_X1 U487 ( .A(n579), .B(KEYINPUT98), .ZN(n378) );
  XNOR2_X1 U488 ( .A(n579), .B(KEYINPUT98), .ZN(n603) );
  BUF_X1 U489 ( .A(n565), .Z(n379) );
  XNOR2_X2 U490 ( .A(n397), .B(n366), .ZN(n380) );
  BUF_X1 U491 ( .A(n750), .Z(n381) );
  XNOR2_X1 U492 ( .A(n551), .B(n417), .ZN(n565) );
  XNOR2_X1 U493 ( .A(n397), .B(n366), .ZN(n396) );
  XNOR2_X2 U494 ( .A(n383), .B(n382), .ZN(n685) );
  NAND2_X1 U495 ( .A1(n557), .A2(n469), .ZN(n383) );
  NOR2_X1 U496 ( .A1(n750), .A2(G902), .ZN(n384) );
  NAND2_X1 U497 ( .A1(n427), .A2(n426), .ZN(n385) );
  NAND2_X1 U498 ( .A1(n427), .A2(n426), .ZN(n640) );
  OR2_X1 U499 ( .A1(n603), .A2(n362), .ZN(n426) );
  XNOR2_X1 U500 ( .A(n496), .B(n471), .ZN(n481) );
  BUF_X1 U501 ( .A(n680), .Z(n386) );
  XNOR2_X1 U502 ( .A(n500), .B(n499), .ZN(n680) );
  BUF_X1 U503 ( .A(n756), .Z(n765) );
  BUF_X1 U504 ( .A(n557), .Z(n606) );
  NAND2_X2 U505 ( .A1(n591), .A2(n592), .ZN(n397) );
  AND2_X1 U506 ( .A1(n630), .A2(n361), .ZN(n391) );
  NAND2_X1 U507 ( .A1(n387), .A2(n418), .ZN(n424) );
  XNOR2_X1 U508 ( .A(n439), .B(n438), .ZN(n437) );
  NAND2_X1 U509 ( .A1(n437), .A2(n436), .ZN(n711) );
  XNOR2_X1 U510 ( .A(n539), .B(n538), .ZN(n543) );
  XNOR2_X1 U511 ( .A(n388), .B(KEYINPUT48), .ZN(n399) );
  NOR2_X2 U512 ( .A1(n798), .A2(n794), .ZN(n617) );
  NAND2_X1 U513 ( .A1(n419), .A2(n422), .ZN(n418) );
  NAND2_X1 U514 ( .A1(n631), .A2(n391), .ZN(n388) );
  NAND2_X1 U515 ( .A1(n398), .A2(n380), .ZN(n655) );
  XNOR2_X2 U516 ( .A(n425), .B(n393), .ZN(n532) );
  XNOR2_X2 U517 ( .A(n506), .B(G134), .ZN(n547) );
  XNOR2_X1 U518 ( .A(n390), .B(KEYINPUT60), .ZN(G60) );
  OR2_X2 U519 ( .A1(n601), .A2(n600), .ZN(n602) );
  BUF_X2 U520 ( .A(n689), .Z(n392) );
  XNOR2_X1 U521 ( .A(n371), .B(n393), .ZN(n507) );
  XNOR2_X2 U522 ( .A(n449), .B(G146), .ZN(n393) );
  NAND2_X1 U523 ( .A1(n572), .A2(n686), .ZN(n395) );
  NOR2_X1 U524 ( .A1(n654), .A2(n399), .ZN(n398) );
  NOR2_X1 U525 ( .A1(n402), .A2(n364), .ZN(n401) );
  INV_X1 U526 ( .A(n443), .ZN(n403) );
  INV_X1 U527 ( .A(n405), .ZN(n404) );
  OR2_X1 U528 ( .A1(n659), .A2(n406), .ZN(n405) );
  NAND2_X1 U529 ( .A1(n659), .A2(n515), .ZN(n410) );
  INV_X1 U530 ( .A(n586), .ZN(n412) );
  XNOR2_X2 U531 ( .A(n413), .B(n365), .ZN(n580) );
  XNOR2_X2 U532 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n415) );
  INV_X1 U533 ( .A(n379), .ZN(n795) );
  XNOR2_X1 U534 ( .A(n416), .B(n568), .ZN(n570) );
  NAND2_X1 U535 ( .A1(n565), .A2(n567), .ZN(n416) );
  NAND2_X1 U536 ( .A1(n396), .A2(n367), .ZN(n423) );
  INV_X1 U537 ( .A(n380), .ZN(n419) );
  NAND2_X1 U538 ( .A1(n424), .A2(n650), .ZN(n656) );
  NOR2_X2 U539 ( .A1(n680), .A2(n580), .ZN(n526) );
  NOR2_X1 U540 ( .A1(n766), .A2(G902), .ZN(n465) );
  XNOR2_X1 U541 ( .A(n465), .B(n464), .ZN(n557) );
  NAND2_X1 U542 ( .A1(n603), .A2(n432), .ZN(n431) );
  XNOR2_X1 U543 ( .A(n434), .B(n512), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n508), .B(n507), .ZN(n434) );
  XNOR2_X1 U545 ( .A(n503), .B(n539), .ZN(n435) );
  NAND2_X1 U546 ( .A1(n440), .A2(n609), .ZN(n439) );
  XNOR2_X1 U547 ( .A(n556), .B(KEYINPUT107), .ZN(n440) );
  NAND2_X1 U548 ( .A1(n446), .A2(n363), .ZN(n738) );
  INV_X1 U549 ( .A(n444), .ZN(n441) );
  NAND2_X1 U550 ( .A1(n445), .A2(n517), .ZN(n444) );
  INV_X1 U551 ( .A(n622), .ZN(n447) );
  AND2_X2 U552 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U553 ( .A(n782), .B(n453), .ZN(n461) );
  AND2_X1 U554 ( .A1(n662), .A2(G953), .ZN(n770) );
  XNOR2_X1 U555 ( .A(n478), .B(G104), .ZN(n448) );
  INV_X2 U556 ( .A(G125), .ZN(n449) );
  INV_X1 U557 ( .A(n683), .ZN(n469) );
  XNOR2_X1 U558 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U559 ( .A1(n379), .A2(n569), .ZN(n566) );
  XNOR2_X1 U560 ( .A(n490), .B(n489), .ZN(n494) );
  INV_X1 U561 ( .A(n478), .ZN(n450) );
  XNOR2_X1 U562 ( .A(n479), .B(n448), .ZN(n480) );
  XNOR2_X1 U563 ( .A(G110), .B(KEYINPUT97), .ZN(n451) );
  XNOR2_X1 U564 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U566 ( .A(n456), .B(KEYINPUT24), .Z(n459) );
  NAND2_X1 U567 ( .A1(G234), .A2(n786), .ZN(n457) );
  XOR2_X1 U568 ( .A(KEYINPUT8), .B(n457), .Z(n544) );
  AND2_X1 U569 ( .A1(n544), .A2(G221), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n461), .B(n460), .ZN(n766) );
  NAND2_X1 U571 ( .A1(G234), .A2(n648), .ZN(n462) );
  XNOR2_X1 U572 ( .A(KEYINPUT20), .B(n462), .ZN(n466) );
  NAND2_X1 U573 ( .A1(G217), .A2(n466), .ZN(n463) );
  XNOR2_X1 U574 ( .A(KEYINPUT25), .B(n463), .ZN(n464) );
  AND2_X1 U575 ( .A1(n466), .A2(G221), .ZN(n468) );
  INV_X1 U576 ( .A(KEYINPUT21), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n468), .B(n467), .ZN(n683) );
  XNOR2_X2 U578 ( .A(G143), .B(G128), .ZN(n506) );
  XOR2_X1 U579 ( .A(G140), .B(KEYINPUT80), .Z(n474) );
  XNOR2_X1 U580 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U581 ( .A(n505), .B(n475), .Z(n477) );
  NAND2_X1 U582 ( .A1(G227), .A2(n786), .ZN(n476) );
  XNOR2_X1 U583 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n481), .B(n480), .ZN(n750) );
  XNOR2_X1 U585 ( .A(KEYINPUT72), .B(G469), .ZN(n482) );
  INV_X1 U586 ( .A(KEYINPUT67), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n483), .B(KEYINPUT1), .ZN(n484) );
  NOR2_X2 U588 ( .A1(n685), .A2(n555), .ZN(n574) );
  NAND2_X1 U589 ( .A1(n535), .A2(G210), .ZN(n485) );
  XNOR2_X1 U590 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X1 U591 ( .A(G113), .B(G101), .ZN(n492) );
  XNOR2_X1 U592 ( .A(KEYINPUT3), .B(G119), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n492), .B(n491), .ZN(n502) );
  INV_X1 U594 ( .A(n502), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U596 ( .A(n496), .B(n495), .ZN(n715) );
  NAND2_X1 U597 ( .A1(n715), .A2(n514), .ZN(n497) );
  INV_X1 U598 ( .A(KEYINPUT6), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n392), .B(n498), .ZN(n559) );
  NAND2_X1 U600 ( .A1(n574), .A2(n559), .ZN(n500) );
  INV_X1 U601 ( .A(G116), .ZN(n501) );
  XNOR2_X1 U602 ( .A(n501), .B(G107), .ZN(n539) );
  XNOR2_X2 U603 ( .A(G122), .B(G104), .ZN(n529) );
  XNOR2_X1 U604 ( .A(n529), .B(KEYINPUT16), .ZN(n503) );
  XNOR2_X1 U605 ( .A(KEYINPUT81), .B(KEYINPUT4), .ZN(n504) );
  XNOR2_X1 U606 ( .A(n505), .B(n504), .ZN(n508) );
  NAND2_X1 U607 ( .A1(G224), .A2(n786), .ZN(n509) );
  XNOR2_X1 U608 ( .A(n509), .B(KEYINPUT17), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U610 ( .A(n648), .ZN(n594) );
  NAND2_X1 U611 ( .A1(n514), .A2(n513), .ZN(n516) );
  AND2_X1 U612 ( .A1(n516), .A2(G210), .ZN(n515) );
  NAND2_X1 U613 ( .A1(n516), .A2(G214), .ZN(n670) );
  INV_X1 U614 ( .A(KEYINPUT19), .ZN(n517) );
  XNOR2_X1 U615 ( .A(n518), .B(KEYINPUT14), .ZN(n521) );
  NAND2_X1 U616 ( .A1(G952), .A2(n521), .ZN(n702) );
  NOR2_X1 U617 ( .A1(G953), .A2(n702), .ZN(n520) );
  INV_X1 U618 ( .A(KEYINPUT92), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n520), .B(n519), .ZN(n599) );
  NAND2_X1 U620 ( .A1(G902), .A2(n521), .ZN(n596) );
  XNOR2_X1 U621 ( .A(G898), .B(KEYINPUT93), .ZN(n777) );
  NAND2_X1 U622 ( .A1(G953), .A2(n777), .ZN(n772) );
  NOR2_X1 U623 ( .A1(n596), .A2(n772), .ZN(n523) );
  INV_X1 U624 ( .A(KEYINPUT94), .ZN(n522) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n524) );
  AND2_X1 U626 ( .A1(n599), .A2(n524), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n526), .B(KEYINPUT34), .ZN(n550) );
  XOR2_X1 U628 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n528) );
  XNOR2_X1 U629 ( .A(G143), .B(KEYINPUT11), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n528), .B(n527), .ZN(n534) );
  XNOR2_X1 U631 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U632 ( .A(n532), .B(n531), .ZN(n533) );
  NOR2_X1 U633 ( .A1(G902), .A2(n758), .ZN(n537) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(G475), .ZN(n536) );
  XNOR2_X1 U635 ( .A(n537), .B(n536), .ZN(n586) );
  XNOR2_X1 U636 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U637 ( .A(n543), .B(n542), .Z(n546) );
  NAND2_X1 U638 ( .A1(G217), .A2(n544), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n546), .B(n545), .ZN(n548) );
  XNOR2_X1 U640 ( .A(n548), .B(n547), .ZN(n762) );
  NOR2_X1 U641 ( .A1(n762), .A2(G902), .ZN(n549) );
  AND2_X1 U642 ( .A1(n586), .A2(n552), .ZN(n637) );
  NAND2_X1 U643 ( .A1(n550), .A2(n637), .ZN(n551) );
  XNOR2_X1 U644 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n560), .A2(n686), .ZN(n556) );
  INV_X1 U646 ( .A(n392), .ZN(n609) );
  INV_X1 U647 ( .A(KEYINPUT106), .ZN(n558) );
  XNOR2_X1 U648 ( .A(n606), .B(n558), .ZN(n682) );
  INV_X1 U649 ( .A(n682), .ZN(n573) );
  NOR2_X1 U650 ( .A1(n686), .A2(n573), .ZN(n561) );
  INV_X1 U651 ( .A(n559), .ZN(n619) );
  NAND2_X1 U652 ( .A1(n561), .A2(n571), .ZN(n563) );
  INV_X1 U653 ( .A(KEYINPUT32), .ZN(n562) );
  XNOR2_X1 U654 ( .A(n563), .B(n562), .ZN(n797) );
  INV_X1 U655 ( .A(n797), .ZN(n564) );
  AND2_X2 U656 ( .A1(n711), .A2(n564), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n566), .A2(KEYINPUT44), .ZN(n592) );
  INV_X1 U658 ( .A(KEYINPUT44), .ZN(n567) );
  INV_X1 U659 ( .A(KEYINPUT68), .ZN(n568) );
  NAND2_X1 U660 ( .A1(n570), .A2(n569), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n571), .B(KEYINPUT86), .ZN(n572) );
  NAND2_X1 U662 ( .A1(n574), .A2(n392), .ZN(n694) );
  OR2_X1 U663 ( .A1(n694), .A2(n580), .ZN(n576) );
  INV_X1 U664 ( .A(KEYINPUT31), .ZN(n575) );
  XNOR2_X1 U665 ( .A(n576), .B(n575), .ZN(n743) );
  INV_X1 U666 ( .A(n685), .ZN(n578) );
  INV_X1 U667 ( .A(n368), .ZN(n577) );
  NOR2_X1 U668 ( .A1(n378), .A2(n392), .ZN(n582) );
  INV_X1 U669 ( .A(n580), .ZN(n581) );
  NAND2_X1 U670 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U671 ( .A(n583), .B(KEYINPUT100), .ZN(n724) );
  NAND2_X1 U672 ( .A1(n743), .A2(n724), .ZN(n587) );
  NOR2_X1 U673 ( .A1(n586), .A2(n585), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n359), .A2(n741), .ZN(n674) );
  NAND2_X1 U675 ( .A1(n587), .A2(n674), .ZN(n588) );
  INV_X1 U676 ( .A(KEYINPUT64), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n689), .A2(n670), .ZN(n595) );
  XNOR2_X1 U678 ( .A(KEYINPUT30), .B(n595), .ZN(n601) );
  NOR2_X1 U679 ( .A1(G900), .A2(n596), .ZN(n597) );
  NAND2_X1 U680 ( .A1(G953), .A2(n597), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n607) );
  INV_X1 U682 ( .A(n607), .ZN(n600) );
  XNOR2_X1 U683 ( .A(n622), .B(KEYINPUT38), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n640), .A2(n741), .ZN(n605) );
  XOR2_X1 U685 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n604) );
  XNOR2_X1 U686 ( .A(n605), .B(n604), .ZN(n798) );
  NOR2_X1 U687 ( .A1(n683), .A2(n606), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n609), .A2(n618), .ZN(n610) );
  XNOR2_X1 U690 ( .A(KEYINPUT28), .B(n610), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n612), .A2(n577), .ZN(n728) );
  INV_X1 U692 ( .A(n613), .ZN(n671) );
  NAND2_X1 U693 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U694 ( .A1(n673), .A2(n675), .ZN(n615) );
  XNOR2_X1 U695 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n614) );
  XNOR2_X1 U696 ( .A(n615), .B(n614), .ZN(n697) );
  NOR2_X1 U697 ( .A1(n728), .A2(n697), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT42), .ZN(n794) );
  XNOR2_X1 U699 ( .A(n617), .B(KEYINPUT46), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n620), .A2(n670), .ZN(n621) );
  INV_X1 U702 ( .A(n369), .ZN(n645) );
  NOR2_X1 U703 ( .A1(n686), .A2(n624), .ZN(n747) );
  XNOR2_X1 U704 ( .A(KEYINPUT76), .B(n674), .ZN(n626) );
  INV_X1 U705 ( .A(KEYINPUT47), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U707 ( .A1(n728), .A2(n627), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n628), .A2(n738), .ZN(n629) );
  NOR2_X1 U709 ( .A1(n747), .A2(n629), .ZN(n630) );
  INV_X1 U710 ( .A(n728), .ZN(n737) );
  AND2_X1 U711 ( .A1(KEYINPUT76), .A2(n674), .ZN(n632) );
  AND2_X1 U712 ( .A1(n737), .A2(n632), .ZN(n633) );
  INV_X1 U713 ( .A(n738), .ZN(n729) );
  NAND2_X1 U714 ( .A1(n633), .A2(n729), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n634), .A2(KEYINPUT47), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n636), .B(KEYINPUT110), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n734) );
  OR2_X1 U718 ( .A1(n385), .A2(n359), .ZN(n749) );
  XOR2_X1 U719 ( .A(n641), .B(KEYINPUT108), .Z(n642) );
  NAND2_X1 U720 ( .A1(n642), .A2(n686), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n643), .B(KEYINPUT109), .ZN(n644) );
  XOR2_X1 U722 ( .A(n644), .B(KEYINPUT43), .Z(n646) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n712) );
  NAND2_X1 U724 ( .A1(n749), .A2(n712), .ZN(n647) );
  NOR2_X2 U725 ( .A1(n399), .A2(n647), .ZN(n784) );
  XNOR2_X1 U726 ( .A(n648), .B(KEYINPUT85), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n649), .A2(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U728 ( .A1(KEYINPUT2), .A2(n749), .ZN(n651) );
  XNOR2_X1 U729 ( .A(KEYINPUT82), .B(n651), .ZN(n653) );
  INV_X1 U730 ( .A(n712), .ZN(n652) );
  OR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n656), .A2(n668), .ZN(n657) );
  XNOR2_X2 U733 ( .A(n657), .B(KEYINPUT65), .ZN(n756) );
  NAND2_X1 U734 ( .A1(n756), .A2(G210), .ZN(n661) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  INV_X1 U737 ( .A(G952), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n664), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U739 ( .A1(n377), .A2(n784), .ZN(n666) );
  INV_X1 U740 ( .A(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n669), .B(KEYINPUT84), .ZN(n707) );
  NOR2_X1 U744 ( .A1(n697), .A2(n386), .ZN(n705) );
  NOR2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n679) );
  INV_X1 U747 ( .A(n674), .ZN(n676) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U749 ( .A(KEYINPUT119), .B(n677), .Z(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n681), .A2(n386), .ZN(n699) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(n684), .Z(n692) );
  XOR2_X1 U754 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n688) );
  NAND2_X1 U755 ( .A1(n686), .A2(n374), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n688), .B(n687), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n690), .A2(n392), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(n695), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U763 ( .A(KEYINPUT52), .B(KEYINPUT120), .ZN(n700) );
  XNOR2_X1 U764 ( .A(n701), .B(n700), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n710), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U769 ( .A(n373), .B(G110), .ZN(G12) );
  XNOR2_X1 U770 ( .A(n712), .B(G140), .ZN(G42) );
  NAND2_X1 U771 ( .A1(n756), .A2(G472), .ZN(n717) );
  XNOR2_X1 U772 ( .A(KEYINPUT90), .B(KEYINPUT113), .ZN(n713) );
  XOR2_X1 U773 ( .A(n713), .B(KEYINPUT62), .Z(n714) );
  XNOR2_X1 U774 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n717), .B(n716), .ZN(n719) );
  INV_X1 U776 ( .A(n770), .ZN(n718) );
  NAND2_X1 U777 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U778 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n721), .B(n720), .ZN(G57) );
  XNOR2_X1 U780 ( .A(n722), .B(G101), .ZN(G3) );
  NOR2_X1 U781 ( .A1(n724), .A2(n741), .ZN(n723) );
  XOR2_X1 U782 ( .A(G104), .B(n723), .Z(G6) );
  NOR2_X1 U783 ( .A1(n724), .A2(n359), .ZN(n726) );
  XNOR2_X1 U784 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n725) );
  XNOR2_X1 U785 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U786 ( .A(G107), .B(n727), .ZN(G9) );
  XOR2_X1 U787 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n732) );
  NOR2_X1 U788 ( .A1(n728), .A2(n359), .ZN(n730) );
  NAND2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U790 ( .A(n732), .B(n731), .ZN(n733) );
  XOR2_X1 U791 ( .A(G128), .B(n733), .Z(G30) );
  XNOR2_X1 U792 ( .A(G143), .B(KEYINPUT116), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n735), .B(n734), .ZN(G45) );
  INV_X1 U794 ( .A(n741), .ZN(n736) );
  NAND2_X1 U795 ( .A1(n737), .A2(n736), .ZN(n739) );
  NOR2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U797 ( .A(G146), .B(n740), .Z(G48) );
  NOR2_X1 U798 ( .A1(n741), .A2(n743), .ZN(n742) );
  XOR2_X1 U799 ( .A(G113), .B(n742), .Z(G15) );
  NOR2_X1 U800 ( .A1(n359), .A2(n743), .ZN(n746) );
  XNOR2_X1 U801 ( .A(G116), .B(KEYINPUT117), .ZN(n745) );
  XNOR2_X1 U802 ( .A(n746), .B(n745), .ZN(G18) );
  XNOR2_X1 U803 ( .A(G125), .B(n747), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n748), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U805 ( .A(G134), .B(n749), .ZN(G36) );
  NAND2_X1 U806 ( .A1(n765), .A2(G469), .ZN(n754) );
  XOR2_X1 U807 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n752) );
  XNOR2_X1 U808 ( .A(n381), .B(KEYINPUT122), .ZN(n751) );
  XNOR2_X1 U809 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U810 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U811 ( .A1(n770), .A2(n755), .ZN(G54) );
  NAND2_X1 U812 ( .A1(n756), .A2(G475), .ZN(n760) );
  XOR2_X1 U813 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n757) );
  XNOR2_X1 U814 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U815 ( .A1(n765), .A2(G478), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U817 ( .A1(n770), .A2(n764), .ZN(G63) );
  NAND2_X1 U818 ( .A1(n765), .A2(G217), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n375), .B(KEYINPUT124), .ZN(n767) );
  XNOR2_X1 U820 ( .A(n768), .B(n767), .ZN(n769) );
  NOR2_X1 U821 ( .A1(n770), .A2(n769), .ZN(G66) );
  XNOR2_X1 U822 ( .A(n771), .B(G110), .ZN(n773) );
  NAND2_X1 U823 ( .A1(n773), .A2(n772), .ZN(n781) );
  BUF_X1 U824 ( .A(n419), .Z(n774) );
  NOR2_X1 U825 ( .A1(n774), .A2(G953), .ZN(n779) );
  NAND2_X1 U826 ( .A1(G953), .A2(G224), .ZN(n775) );
  XOR2_X1 U827 ( .A(KEYINPUT61), .B(n775), .Z(n776) );
  NOR2_X1 U828 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U829 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U830 ( .A(n781), .B(n780), .ZN(G69) );
  XNOR2_X1 U831 ( .A(n782), .B(n783), .ZN(n788) );
  INV_X1 U832 ( .A(n788), .ZN(n785) );
  XNOR2_X1 U833 ( .A(n785), .B(n784), .ZN(n787) );
  NAND2_X1 U834 ( .A1(n787), .A2(n786), .ZN(n792) );
  XNOR2_X1 U835 ( .A(G227), .B(n788), .ZN(n789) );
  NAND2_X1 U836 ( .A1(n789), .A2(G900), .ZN(n790) );
  NAND2_X1 U837 ( .A1(n790), .A2(G953), .ZN(n791) );
  NAND2_X1 U838 ( .A1(n792), .A2(n791), .ZN(G72) );
  XOR2_X1 U839 ( .A(G137), .B(KEYINPUT126), .Z(n793) );
  XNOR2_X1 U840 ( .A(n794), .B(n793), .ZN(G39) );
  XNOR2_X1 U841 ( .A(G122), .B(n795), .ZN(n796) );
  XNOR2_X1 U842 ( .A(n796), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U843 ( .A(G119), .B(n797), .Z(G21) );
  XNOR2_X1 U844 ( .A(G131), .B(KEYINPUT127), .ZN(n799) );
  XNOR2_X1 U845 ( .A(n799), .B(n376), .ZN(G33) );
endmodule

