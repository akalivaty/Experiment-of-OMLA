

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595;

  NOR2_X1 U325 ( .A1(n394), .A2(n393), .ZN(n493) );
  XOR2_X1 U326 ( .A(KEYINPUT41), .B(n586), .Z(n561) );
  NOR2_X1 U327 ( .A1(n532), .A2(n554), .ZN(n539) );
  XNOR2_X1 U328 ( .A(n419), .B(KEYINPUT104), .ZN(n420) );
  XNOR2_X1 U329 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U330 ( .A(KEYINPUT54), .B(n480), .Z(n293) );
  AND2_X1 U331 ( .A1(n561), .A2(n582), .ZN(n463) );
  INV_X1 U332 ( .A(KEYINPUT47), .ZN(n467) );
  XOR2_X1 U333 ( .A(G99GAT), .B(G85GAT), .Z(n446) );
  XNOR2_X1 U334 ( .A(n467), .B(KEYINPUT113), .ZN(n468) );
  XNOR2_X1 U335 ( .A(n367), .B(KEYINPUT95), .ZN(n368) );
  XNOR2_X1 U336 ( .A(n469), .B(n468), .ZN(n476) );
  XNOR2_X1 U337 ( .A(n369), .B(n368), .ZN(n371) );
  XNOR2_X1 U338 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n477) );
  XNOR2_X1 U339 ( .A(n376), .B(n375), .ZN(n377) );
  NOR2_X1 U340 ( .A1(n527), .A2(n293), .ZN(n579) );
  XNOR2_X1 U341 ( .A(n374), .B(n305), .ZN(n306) );
  XNOR2_X1 U342 ( .A(n421), .B(n420), .ZN(n524) );
  XNOR2_X1 U343 ( .A(n307), .B(n306), .ZN(n311) );
  NOR2_X1 U344 ( .A1(n484), .A2(n483), .ZN(n577) );
  XOR2_X1 U345 ( .A(n481), .B(KEYINPUT28), .Z(n532) );
  XNOR2_X1 U346 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U347 ( .A(n460), .B(G43GAT), .ZN(n461) );
  XNOR2_X1 U348 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  INV_X1 U350 ( .A(KEYINPUT36), .ZN(n312) );
  XOR2_X1 U351 ( .A(G50GAT), .B(G162GAT), .Z(n332) );
  XOR2_X1 U352 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n295) );
  XNOR2_X1 U353 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n294) );
  XNOR2_X1 U354 ( .A(n295), .B(n294), .ZN(n297) );
  INV_X1 U355 ( .A(n297), .ZN(n296) );
  NAND2_X1 U356 ( .A1(n332), .A2(n296), .ZN(n300) );
  INV_X1 U357 ( .A(n332), .ZN(n298) );
  NAND2_X1 U358 ( .A1(n298), .A2(n297), .ZN(n299) );
  NAND2_X1 U359 ( .A1(n300), .A2(n299), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n446), .B(G106GAT), .ZN(n302) );
  AND2_X1 U361 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U362 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n307) );
  XOR2_X1 U364 ( .A(G36GAT), .B(G190GAT), .Z(n374) );
  XNOR2_X1 U365 ( .A(G134GAT), .B(G218GAT), .ZN(n305) );
  XOR2_X1 U366 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n309) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(KEYINPUT69), .B(n310), .Z(n441) );
  XOR2_X1 U370 ( .A(n311), .B(n441), .Z(n568) );
  XNOR2_X1 U371 ( .A(n312), .B(n568), .ZN(n470) );
  XOR2_X1 U372 ( .A(G148GAT), .B(G155GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(G127GAT), .B(G162GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U375 ( .A(n315), .B(G85GAT), .Z(n317) );
  XOR2_X1 U376 ( .A(G113GAT), .B(G1GAT), .Z(n433) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(n433), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U379 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n319) );
  XNOR2_X1 U380 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U382 ( .A(n321), .B(n320), .Z(n326) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(G120GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n322), .B(KEYINPUT0), .ZN(n354) );
  XOR2_X1 U385 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n324) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n354), .B(n336), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n331) );
  XOR2_X1 U390 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n328) );
  NAND2_X1 U391 ( .A1(G225GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U393 ( .A(KEYINPUT1), .B(n329), .Z(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n527) );
  INV_X1 U395 ( .A(KEYINPUT97), .ZN(n388) );
  XOR2_X1 U396 ( .A(G22GAT), .B(G155GAT), .Z(n404) );
  XNOR2_X1 U397 ( .A(n332), .B(n404), .ZN(n335) );
  XOR2_X1 U398 ( .A(G78GAT), .B(G148GAT), .Z(n334) );
  XNOR2_X1 U399 ( .A(G106GAT), .B(G204GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n442) );
  XNOR2_X1 U401 ( .A(n335), .B(n442), .ZN(n340) );
  XOR2_X1 U402 ( .A(n336), .B(KEYINPUT24), .Z(n338) );
  NAND2_X1 U403 ( .A1(G228GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U405 ( .A(n340), .B(n339), .Z(n349) );
  XNOR2_X1 U406 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n341), .B(KEYINPUT89), .ZN(n342) );
  XOR2_X1 U408 ( .A(n342), .B(KEYINPUT21), .Z(n344) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G218GAT), .ZN(n343) );
  XNOR2_X1 U410 ( .A(n344), .B(n343), .ZN(n380) );
  XOR2_X1 U411 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n346) );
  XNOR2_X1 U412 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n380), .B(n347), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n481) );
  INV_X1 U416 ( .A(n481), .ZN(n382) );
  XOR2_X1 U417 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n351) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n369) );
  XOR2_X1 U420 ( .A(G15GAT), .B(G127GAT), .Z(n405) );
  XOR2_X1 U421 ( .A(n369), .B(n405), .Z(n353) );
  XNOR2_X1 U422 ( .A(G43GAT), .B(G99GAT), .ZN(n352) );
  XNOR2_X1 U423 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U424 ( .A(n354), .B(G113GAT), .Z(n356) );
  NAND2_X1 U425 ( .A1(G227GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U426 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U427 ( .A(n358), .B(n357), .Z(n366) );
  XOR2_X1 U428 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n360) );
  XNOR2_X1 U429 ( .A(G190GAT), .B(KEYINPUT86), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U431 ( .A(KEYINPUT84), .B(G71GAT), .Z(n362) );
  XNOR2_X1 U432 ( .A(G183GAT), .B(G176GAT), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n484) );
  AND2_X1 U436 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  INV_X1 U437 ( .A(KEYINPUT94), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n378) );
  XNOR2_X1 U439 ( .A(G176GAT), .B(G92GAT), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n372), .B(G64GAT), .ZN(n445) );
  XNOR2_X1 U441 ( .A(G8GAT), .B(G183GAT), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n373), .B(KEYINPUT78), .ZN(n412) );
  XNOR2_X1 U443 ( .A(n445), .B(n412), .ZN(n376) );
  XNOR2_X1 U444 ( .A(G204GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n479) );
  NOR2_X1 U446 ( .A1(n484), .A2(n479), .ZN(n381) );
  NOR2_X1 U447 ( .A1(n382), .A2(n381), .ZN(n383) );
  XOR2_X1 U448 ( .A(KEYINPUT25), .B(n383), .Z(n386) );
  INV_X1 U449 ( .A(n484), .ZN(n538) );
  NOR2_X1 U450 ( .A1(n481), .A2(n538), .ZN(n384) );
  XNOR2_X1 U451 ( .A(KEYINPUT26), .B(n384), .ZN(n580) );
  INV_X1 U452 ( .A(n479), .ZN(n529) );
  XNOR2_X1 U453 ( .A(KEYINPUT27), .B(n529), .ZN(n390) );
  AND2_X1 U454 ( .A1(n580), .A2(n390), .ZN(n385) );
  NOR2_X1 U455 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n389) );
  NOR2_X1 U457 ( .A1(n527), .A2(n389), .ZN(n394) );
  NAND2_X1 U458 ( .A1(n527), .A2(n390), .ZN(n554) );
  INV_X1 U459 ( .A(KEYINPUT96), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n539), .B(n391), .ZN(n392) );
  NOR2_X1 U461 ( .A1(n538), .A2(n392), .ZN(n393) );
  XOR2_X1 U462 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n396) );
  XNOR2_X1 U463 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U465 ( .A(KEYINPUT80), .B(G64GAT), .Z(n398) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n416) );
  XOR2_X1 U469 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n402) );
  XNOR2_X1 U470 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U472 ( .A(G57GAT), .B(n403), .Z(n454) );
  XOR2_X1 U473 ( .A(G78GAT), .B(n404), .Z(n407) );
  XNOR2_X1 U474 ( .A(n405), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U476 ( .A(n454), .B(n408), .Z(n410) );
  NAND2_X1 U477 ( .A1(G231GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n411), .B(KEYINPUT12), .ZN(n414) );
  XOR2_X1 U480 ( .A(n412), .B(KEYINPUT82), .Z(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n416), .B(n415), .ZN(n489) );
  INV_X1 U483 ( .A(n489), .ZN(n590) );
  NOR2_X1 U484 ( .A1(n493), .A2(n590), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n417), .B(KEYINPUT103), .ZN(n418) );
  NOR2_X1 U486 ( .A1(n470), .A2(n418), .ZN(n421) );
  INV_X1 U487 ( .A(KEYINPUT37), .ZN(n419) );
  XOR2_X1 U488 ( .A(KEYINPUT30), .B(G15GAT), .Z(n423) );
  XNOR2_X1 U489 ( .A(G169GAT), .B(G197GAT), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U491 ( .A(KEYINPUT67), .B(G8GAT), .Z(n425) );
  XNOR2_X1 U492 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U494 ( .A(n427), .B(n426), .Z(n439) );
  XOR2_X1 U495 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n429) );
  XNOR2_X1 U496 ( .A(KEYINPUT71), .B(KEYINPUT65), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n437) );
  XOR2_X1 U498 ( .A(G22GAT), .B(G141GAT), .Z(n431) );
  XNOR2_X1 U499 ( .A(G50GAT), .B(G36GAT), .ZN(n430) );
  XNOR2_X1 U500 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U501 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U502 ( .A1(G229GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U504 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U505 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n441), .B(n440), .ZN(n582) );
  INV_X1 U507 ( .A(n582), .ZN(n557) );
  XNOR2_X1 U508 ( .A(n442), .B(KEYINPUT33), .ZN(n444) );
  AND2_X1 U509 ( .A1(G230GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U510 ( .A(n444), .B(n443), .ZN(n450) );
  XNOR2_X1 U511 ( .A(KEYINPUT75), .B(n445), .ZN(n448) );
  XNOR2_X1 U512 ( .A(G120GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U514 ( .A(n450), .B(n449), .ZN(n456) );
  XOR2_X1 U515 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n452) );
  XNOR2_X1 U516 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n451) );
  XNOR2_X1 U517 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n586) );
  NOR2_X1 U520 ( .A1(n557), .A2(n586), .ZN(n457) );
  XOR2_X1 U521 ( .A(KEYINPUT77), .B(n457), .Z(n494) );
  NAND2_X1 U522 ( .A1(n524), .A2(n494), .ZN(n458) );
  XNOR2_X1 U523 ( .A(n458), .B(KEYINPUT105), .ZN(n459) );
  XNOR2_X1 U524 ( .A(KEYINPUT38), .B(n459), .ZN(n511) );
  NAND2_X1 U525 ( .A1(n511), .A2(n538), .ZN(n462) );
  XOR2_X1 U526 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n460) );
  XNOR2_X1 U527 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U529 ( .A1(n568), .A2(n465), .ZN(n466) );
  NAND2_X1 U530 ( .A1(n489), .A2(n466), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n489), .A2(n470), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT45), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n557), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n586), .A2(n473), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT114), .B(n474), .ZN(n475) );
  NOR2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n537) );
  NOR2_X1 U538 ( .A1(n537), .A2(n479), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n481), .A2(n579), .ZN(n482) );
  XOR2_X1 U540 ( .A(n482), .B(KEYINPUT55), .Z(n483) );
  NAND2_X1 U541 ( .A1(n577), .A2(n568), .ZN(n488) );
  XOR2_X1 U542 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n486) );
  INV_X1 U543 ( .A(G190GAT), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n491) );
  OR2_X1 U545 ( .A1(n489), .A2(n568), .ZN(n490) );
  XNOR2_X1 U546 ( .A(n491), .B(n490), .ZN(n492) );
  NOR2_X1 U547 ( .A1(n493), .A2(n492), .ZN(n513) );
  NAND2_X1 U548 ( .A1(n513), .A2(n494), .ZN(n495) );
  XOR2_X1 U549 ( .A(KEYINPUT98), .B(n495), .Z(n505) );
  NAND2_X1 U550 ( .A1(n505), .A2(n527), .ZN(n499) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n497) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n496) );
  XNOR2_X1 U553 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U554 ( .A(n499), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n505), .A2(n529), .ZN(n500) );
  XNOR2_X1 U556 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n502) );
  NAND2_X1 U558 ( .A1(n505), .A2(n538), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n502), .B(n501), .ZN(n504) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT101), .Z(n503) );
  XNOR2_X1 U561 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  NAND2_X1 U562 ( .A1(n505), .A2(n532), .ZN(n506) );
  XNOR2_X1 U563 ( .A(n506), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .Z(n508) );
  NAND2_X1 U565 ( .A1(n511), .A2(n527), .ZN(n507) );
  XNOR2_X1 U566 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT106), .ZN(n510) );
  NAND2_X1 U568 ( .A1(n529), .A2(n511), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n510), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n511), .A2(n532), .ZN(n512) );
  XNOR2_X1 U571 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U572 ( .A(n561), .B(KEYINPUT108), .ZN(n572) );
  NAND2_X1 U573 ( .A1(n557), .A2(n572), .ZN(n525) );
  INV_X1 U574 ( .A(n513), .ZN(n514) );
  NOR2_X1 U575 ( .A1(n525), .A2(n514), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n521), .A2(n527), .ZN(n515) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n515), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  XOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT109), .Z(n518) );
  NAND2_X1 U580 ( .A1(n521), .A2(n529), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n538), .A2(n521), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(n520), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U586 ( .A1(n521), .A2(n532), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  INV_X1 U588 ( .A(n524), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n533), .A2(n529), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n538), .A2(n533), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n535) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n542) );
  BUF_X1 U601 ( .A(n537), .Z(n555) );
  NAND2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U603 ( .A1(n555), .A2(n540), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n551), .A2(n582), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U608 ( .A1(n551), .A2(n572), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n548) );
  NAND2_X1 U613 ( .A1(n551), .A2(n590), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n568), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n556), .A2(n580), .ZN(n560) );
  NOR2_X1 U621 ( .A1(n557), .A2(n560), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(n558), .Z(n559) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n563) );
  INV_X1 U625 ( .A(n560), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(n564), .B(KEYINPUT52), .Z(n566) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n590), .A2(n569), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U635 ( .A1(n582), .A2(n577), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT57), .Z(n574) );
  NAND2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U642 ( .A1(n590), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n584) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT125), .ZN(n592) );
  NAND2_X1 U647 ( .A1(n592), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U651 ( .A1(n592), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(n589), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n592), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U656 ( .A(n592), .ZN(n593) );
  NOR2_X1 U657 ( .A1(n470), .A2(n593), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

