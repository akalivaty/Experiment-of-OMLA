//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  AOI21_X1  g004(.A(KEYINPUT74), .B1(new_n190), .B2(G140), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(G140), .ZN(new_n192));
  OAI211_X1 g006(.A(KEYINPUT16), .B(new_n189), .C1(new_n191), .C2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT75), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G125), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n188), .A2(G125), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(KEYINPUT74), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n199), .A2(KEYINPUT75), .A3(KEYINPUT16), .A4(new_n189), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n196), .A2(new_n200), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT24), .B(G110), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(KEYINPUT72), .A3(KEYINPUT23), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G119), .A3(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n208), .A2(G119), .B1(KEYINPUT72), .B2(KEYINPUT23), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT73), .B1(new_n219), .B2(G110), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n213), .B2(new_n215), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n222));
  INV_X1    g036(.A(G110), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n212), .A3(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n192), .A2(new_n198), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n210), .A2(new_n211), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n202), .A2(new_n231), .A3(KEYINPUT76), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT76), .B1(new_n202), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G953), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(G221), .A3(G234), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT77), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT22), .B(G137), .Z(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT78), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n226), .B(new_n239), .C1(new_n232), .C2(new_n233), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n241), .A2(KEYINPUT25), .A3(new_n242), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G234), .ZN(new_n249));
  OAI21_X1  g063(.A(G217), .B1(new_n249), .B2(G902), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT79), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT79), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n254), .A3(new_n251), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n241), .A2(new_n243), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n251), .A2(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G113), .B(G122), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT88), .B(G104), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n203), .B1(new_n196), .B2(new_n200), .ZN(new_n264));
  NOR2_X1   g078(.A1(G237), .A2(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G214), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G143), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n266), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n199), .A2(new_n189), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(KEYINPUT19), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n264), .B(new_n271), .C1(new_n203), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT18), .A2(G131), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n269), .B(new_n276), .Z(new_n277));
  AOI21_X1  g091(.A(new_n228), .B1(new_n273), .B2(G146), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n263), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n269), .A2(KEYINPUT17), .A3(G131), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n202), .A2(new_n204), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT89), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n202), .A2(new_n286), .A3(new_n204), .A4(new_n281), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n279), .ZN(new_n289));
  INV_X1    g103(.A(new_n263), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G475), .A2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT20), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n290), .B1(new_n288), .B2(new_n289), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n242), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G475), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n292), .A2(KEYINPUT90), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n280), .A2(new_n291), .A3(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n302), .A2(KEYINPUT20), .A3(new_n293), .A4(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G128), .B(G143), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT13), .ZN(new_n307));
  INV_X1    g121(.A(G143), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G128), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n307), .B(G134), .C1(KEYINPUT13), .C2(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(G116), .B(G122), .Z(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G107), .ZN(new_n312));
  XNOR2_X1  g126(.A(G116), .B(G122), .ZN(new_n313));
  INV_X1    g127(.A(G107), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n306), .B(new_n317), .ZN(new_n320));
  INV_X1    g134(.A(G116), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT14), .A3(G122), .ZN(new_n322));
  OAI211_X1 g136(.A(G107), .B(new_n322), .C1(new_n311), .C2(KEYINPUT14), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT9), .B(G234), .Z(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(G217), .A3(new_n235), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n325), .A2(new_n327), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G478), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(KEYINPUT15), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT92), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n242), .A3(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(KEYINPUT93), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT91), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n330), .B2(G902), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT91), .B(new_n242), .C1(new_n328), .C2(new_n329), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n333), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(KEYINPUT93), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n301), .A2(new_n305), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G104), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n346), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n314), .A3(G104), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(G107), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n346), .A2(G107), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n314), .A2(G104), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G143), .B(G146), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n208), .A2(new_n203), .A3(G143), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n308), .B(G146), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n352), .A2(new_n355), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n352), .B2(new_n355), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT10), .B(new_n363), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G101), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT0), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n358), .B1(new_n374), .B2(new_n208), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT0), .B(G128), .Z(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n358), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n370), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT64), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n382), .A2(KEYINPUT11), .B1(new_n317), .B2(G137), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n384));
  INV_X1    g198(.A(G137), .ZN(new_n385));
  AND4_X1   g199(.A1(KEYINPUT64), .A2(new_n384), .A3(new_n385), .A4(G134), .ZN(new_n386));
  AOI22_X1  g200(.A1(KEYINPUT64), .A2(new_n384), .B1(new_n385), .B2(G134), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G131), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n270), .B(new_n383), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(KEYINPUT65), .A3(G131), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n393), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(new_n366), .A3(new_n380), .A4(new_n370), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(G110), .B(G140), .Z(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT80), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n235), .A2(G227), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n397), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(new_n402), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT82), .B1(new_n357), .B2(new_n363), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n356), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n411), .A3(new_n364), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n394), .A2(new_n412), .A3(KEYINPUT12), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT12), .B1(new_n394), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n398), .A2(KEYINPUT84), .A3(new_n402), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n405), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n242), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(new_n395), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n394), .A2(new_n412), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n406), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n402), .B1(new_n425), .B2(KEYINPUT83), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT83), .B(new_n397), .C1(new_n414), .C2(new_n415), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(G469), .B(new_n421), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G469), .A2(G902), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G221), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n326), .B2(new_n242), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT2), .B(G113), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(G116), .B(G119), .Z(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n373), .A2(new_n442), .A3(new_n379), .ZN(new_n443));
  XOR2_X1   g257(.A(G110), .B(G122), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n368), .A2(new_n369), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n206), .A3(G116), .ZN(new_n448));
  OAI211_X1 g262(.A(G113), .B(new_n448), .C1(new_n440), .C2(new_n447), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n439), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n443), .B(new_n445), .C1(new_n446), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n377), .A2(G125), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(G125), .B2(new_n409), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n235), .A2(G224), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT7), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT86), .B1(new_n450), .B2(new_n356), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n450), .A2(new_n356), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n457), .B(new_n458), .Z(new_n459));
  XNOR2_X1  g273(.A(new_n444), .B(KEYINPUT8), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n451), .B(new_n456), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n446), .A2(new_n450), .ZN(new_n462));
  INV_X1    g276(.A(new_n443), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n444), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n444), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n454), .B(KEYINPUT85), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n453), .B(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n461), .A2(new_n470), .A3(new_n242), .ZN(new_n471));
  OAI21_X1  g285(.A(G210), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n475), .A2(G952), .A3(new_n235), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(G902), .A3(G953), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT94), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n345), .A2(new_n435), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n392), .A2(new_n393), .A3(new_n377), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n385), .A2(G134), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n317), .A2(G137), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n363), .A2(new_n391), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n391), .A2(new_n490), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n391), .A2(KEYINPUT66), .A3(new_n490), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n363), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n487), .B1(new_n486), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n485), .B(new_n442), .C1(new_n492), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n442), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n392), .A2(new_n393), .A3(new_n377), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n496), .A2(new_n363), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT66), .B1(new_n391), .B2(new_n490), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT30), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n486), .A2(new_n497), .A3(new_n500), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT67), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n499), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n265), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n350), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT31), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT31), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n486), .A2(new_n491), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n442), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n522), .B2(new_n508), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n508), .A2(new_n524), .A3(new_n520), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n508), .B2(new_n520), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT69), .B1(new_n527), .B2(new_n515), .ZN(new_n528));
  INV_X1    g342(.A(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n508), .A2(new_n524), .A3(new_n520), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n522), .A2(new_n508), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n520), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n514), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n517), .A2(new_n519), .A3(new_n528), .A4(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G472), .A2(G902), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT32), .B1(new_n535), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n508), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n500), .B1(new_n486), .B2(new_n497), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT28), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n515), .A2(KEYINPUT29), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n529), .A3(new_n530), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n242), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT70), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n532), .A2(new_n515), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n510), .A2(new_n514), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT29), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G472), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT71), .B1(new_n539), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n535), .A2(new_n536), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n555));
  AND4_X1   g369(.A1(KEYINPUT71), .A2(new_n554), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n260), .B(new_n484), .C1(new_n551), .C2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(G101), .ZN(G3));
  NOR2_X1   g372(.A1(new_n259), .A2(new_n435), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n535), .A2(new_n242), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n560), .A2(G472), .B1(new_n536), .B2(new_n535), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n330), .A2(KEYINPUT33), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n330), .A2(KEYINPUT33), .ZN(new_n564));
  AND4_X1   g378(.A1(G478), .A2(new_n563), .A3(new_n242), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(G478), .B1(new_n338), .B2(new_n339), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n480), .B(new_n567), .C1(new_n301), .C2(new_n305), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n474), .A2(new_n569), .A3(new_n482), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n569), .B1(new_n474), .B2(new_n482), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n562), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT34), .B(G104), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G6));
  XOR2_X1   g390(.A(new_n300), .B(KEYINPUT96), .Z(new_n577));
  AND2_X1   g391(.A1(new_n302), .A2(new_n304), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n293), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n295), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n577), .A2(new_n580), .A3(new_n305), .A4(new_n343), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n480), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n562), .A2(new_n582), .A3(new_n573), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  AOI21_X1  g399(.A(new_n254), .B1(new_n248), .B2(new_n251), .ZN(new_n586));
  AOI211_X1 g400(.A(KEYINPUT79), .B(new_n250), .C1(new_n246), .C2(new_n247), .ZN(new_n587));
  OR3_X1    g401(.A1(new_n234), .A2(new_n240), .A3(KEYINPUT36), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n234), .B1(new_n240), .B2(KEYINPUT36), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n257), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT97), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n588), .A2(new_n592), .A3(new_n257), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n586), .A2(new_n587), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n435), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n345), .A2(new_n483), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n561), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n223), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n598), .B(new_n600), .ZN(G12));
  NAND3_X1  g415(.A1(new_n554), .A2(new_n550), .A3(new_n555), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT71), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n554), .A2(new_n550), .A3(KEYINPUT71), .A4(new_n555), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n474), .A2(new_n482), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT95), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n570), .ZN(new_n609));
  INV_X1    g423(.A(G900), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n476), .B1(new_n478), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n581), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(new_n596), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G128), .ZN(G30));
  AOI21_X1  g428(.A(new_n344), .B1(new_n301), .B2(new_n305), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n482), .ZN(new_n616));
  INV_X1    g430(.A(new_n595), .ZN(new_n617));
  OR3_X1    g431(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n554), .A2(new_n555), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n510), .A2(new_n514), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n540), .A2(new_n541), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n622), .B2(new_n514), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n474), .B(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT100), .B1(new_n616), .B2(new_n617), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n618), .A2(new_n625), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n611), .B(KEYINPUT39), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n435), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  AOI211_X1 g453(.A(new_n611), .B(new_n567), .C1(new_n301), .C2(new_n305), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n606), .A2(new_n573), .A3(new_n596), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT103), .B(G146), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G48));
  AOI21_X1  g457(.A(new_n259), .B1(new_n604), .B2(new_n605), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n418), .A2(new_n242), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G469), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n420), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n433), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n573), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n568), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  NAND4_X1  g467(.A1(new_n606), .A2(new_n260), .A3(new_n582), .A4(new_n650), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G116), .ZN(G18));
  NOR3_X1   g469(.A1(new_n649), .A2(new_n345), .A3(new_n595), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n606), .A3(new_n481), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G119), .ZN(G21));
  AND3_X1   g472(.A1(new_n542), .A2(new_n529), .A3(new_n530), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n517), .B(new_n519), .C1(new_n515), .C2(new_n659), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n560), .A2(G472), .B1(new_n536), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n260), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n615), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n609), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n663), .A2(new_n481), .A3(new_n648), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT104), .B(G122), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G24));
  AND2_X1   g482(.A1(new_n661), .A2(new_n617), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n650), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G125), .ZN(G27));
  XNOR2_X1  g485(.A(new_n430), .B(KEYINPUT105), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n420), .A2(new_n429), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n434), .A2(new_n482), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n474), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n606), .A2(new_n260), .A3(new_n640), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n602), .A2(KEYINPUT42), .A3(new_n260), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n640), .A4(new_n680), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n602), .A2(KEYINPUT42), .A3(new_n260), .A4(new_n640), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT108), .B1(new_n687), .B2(new_n679), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G131), .ZN(G33));
  NOR2_X1   g505(.A1(new_n581), .A2(new_n611), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n644), .A2(new_n692), .A3(new_n680), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G134), .ZN(G36));
  OR2_X1    g512(.A1(new_n565), .A2(new_n566), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n301), .A2(new_n305), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT43), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT43), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n561), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(KEYINPUT110), .A3(KEYINPUT44), .A4(new_n617), .ZN(new_n706));
  INV_X1    g520(.A(new_n482), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n474), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n704), .A3(new_n617), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n706), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n421), .B1(new_n426), .B2(new_n428), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(G469), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(KEYINPUT46), .A3(new_n673), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n420), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT46), .B1(new_n720), .B2(new_n673), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n434), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(new_n634), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n715), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G137), .ZN(G39));
  XOR2_X1   g541(.A(new_n724), .B(KEYINPUT47), .Z(new_n728));
  INV_X1    g542(.A(new_n606), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n640), .A2(new_n259), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n708), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G140), .ZN(G42));
  NOR3_X1   g546(.A1(new_n625), .A2(new_n259), .A3(new_n700), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n647), .A2(KEYINPUT49), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n677), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n647), .A2(KEYINPUT49), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n627), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n701), .A2(new_n476), .A3(new_n702), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT115), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n701), .A2(new_n740), .A3(new_n476), .A4(new_n702), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n662), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n707), .A3(new_n627), .A4(new_n648), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n647), .A2(new_n434), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n708), .B(new_n742), .C1(new_n728), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n739), .A2(new_n741), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n647), .A2(new_n474), .A3(new_n677), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n669), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n619), .A2(new_n624), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n260), .A2(new_n752), .A3(new_n476), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n301), .A2(new_n305), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n755), .A3(new_n567), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n745), .A2(new_n747), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n747), .A2(new_n751), .A3(new_n756), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n747), .B2(new_n758), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n745), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n259), .B1(new_n539), .B2(new_n550), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n750), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT48), .ZN(new_n769));
  INV_X1    g583(.A(G952), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n755), .A2(new_n567), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n770), .B(G953), .C1(new_n753), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n742), .A2(new_n650), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n766), .A2(new_n769), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n772), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n762), .B2(new_n765), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT117), .A3(new_n769), .A4(new_n773), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n657), .A2(new_n654), .A3(new_n666), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  INV_X1    g596(.A(new_n607), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n559), .A2(new_n561), .A3(new_n568), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n598), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n644), .B2(new_n484), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n343), .A2(new_n305), .A3(new_n296), .A4(new_n300), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n301), .A2(KEYINPUT111), .A3(new_n305), .A4(new_n343), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT112), .B1(new_n792), .B2(new_n483), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n794), .A3(new_n481), .A4(new_n783), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n562), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n782), .B1(new_n786), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n785), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n782), .A2(new_n557), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n651), .B(new_n781), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n606), .A2(new_n596), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n577), .A2(new_n305), .A3(new_n580), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n343), .A3(new_n611), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n708), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n680), .A2(new_n669), .A3(new_n640), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n690), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n609), .A2(new_n664), .A3(new_n433), .A4(new_n611), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n625), .A3(new_n595), .A4(new_n676), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n641), .A2(new_n613), .A3(new_n810), .A4(new_n670), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n641), .A2(new_n670), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .A3(new_n613), .A4(new_n810), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n808), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n806), .A2(new_n816), .A3(KEYINPUT53), .A4(new_n697), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  INV_X1    g632(.A(new_n807), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n683), .B2(new_n689), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n811), .A2(new_n812), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n811), .A2(new_n812), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n697), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n557), .A2(new_n796), .A3(new_n798), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT113), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n786), .A2(new_n782), .A3(new_n796), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n651), .A3(new_n804), .A4(new_n781), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n818), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n817), .A2(new_n829), .A3(KEYINPUT114), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n817), .A2(new_n829), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n817), .A2(new_n829), .A3(new_n830), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n780), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(G952), .A2(G953), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n737), .B1(new_n837), .B2(new_n838), .ZN(G75));
  AOI21_X1  g653(.A(new_n242), .B1(new_n817), .B2(new_n829), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT56), .B1(new_n840), .B2(G210), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n465), .A2(new_n467), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(new_n469), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT55), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n841), .A2(new_n844), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n235), .A2(G952), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G51));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n833), .A2(new_n849), .A3(new_n835), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n832), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n672), .B(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n418), .ZN(new_n854));
  INV_X1    g668(.A(new_n720), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n840), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n847), .B1(new_n854), .B2(new_n856), .ZN(G54));
  NAND2_X1  g671(.A1(KEYINPUT58), .A2(G475), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT119), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n840), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(new_n578), .Z(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n847), .ZN(G60));
  NAND2_X1  g676(.A1(G478), .A2(G902), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT59), .Z(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n836), .A2(new_n831), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n563), .A2(new_n564), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT120), .Z(new_n868));
  AOI21_X1  g682(.A(new_n847), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n864), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n850), .A2(new_n851), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n850), .A2(KEYINPUT121), .A3(new_n851), .A4(new_n870), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n869), .A2(new_n873), .A3(new_n874), .ZN(G63));
  INV_X1    g689(.A(new_n847), .ZN(new_n876));
  NAND2_X1  g690(.A1(G217), .A2(G902), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT60), .Z(new_n878));
  NAND4_X1  g692(.A1(new_n832), .A2(new_n588), .A3(new_n589), .A4(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n832), .A2(new_n878), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n876), .B(new_n879), .C1(new_n880), .C2(new_n256), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT61), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT61), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(G66));
  INV_X1    g700(.A(G224), .ZN(new_n887));
  OAI21_X1  g701(.A(G953), .B1(new_n479), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n800), .B(KEYINPUT123), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n842), .B1(G898), .B2(new_n235), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(G69));
  NOR2_X1   g706(.A1(new_n492), .A2(new_n498), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n274), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n792), .B1(new_n755), .B2(new_n567), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n644), .A2(new_n635), .A3(new_n708), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n726), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n814), .A2(new_n613), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n638), .ZN(new_n899));
  XOR2_X1   g713(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n900));
  OAI211_X1 g714(.A(new_n897), .B(new_n731), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n898), .B2(new_n638), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n235), .B(new_n894), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n235), .B1(G227), .B2(G900), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT126), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n767), .A2(new_n665), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n715), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n725), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n696), .B2(new_n695), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n898), .A2(new_n690), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n731), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT125), .A4(new_n731), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n235), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(G900), .A2(G953), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n904), .B(new_n906), .C1(new_n918), .C2(new_n894), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n905), .A2(KEYINPUT126), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G72));
  NAND2_X1  g735(.A1(G472), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT63), .Z(new_n923));
  AND4_X1   g737(.A1(new_n548), .A2(new_n832), .A3(new_n621), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n901), .A2(new_n903), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n889), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n621), .B1(new_n926), .B2(new_n923), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n914), .A2(new_n889), .A3(new_n915), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n923), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n928), .B(new_n876), .C1(new_n930), .C2(new_n548), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n548), .B1(new_n929), .B2(new_n923), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT127), .B1(new_n932), .B2(new_n847), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n924), .B(new_n927), .C1(new_n931), .C2(new_n933), .ZN(G57));
endmodule


