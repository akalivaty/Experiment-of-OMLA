

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769;

  INV_X1 U373 ( .A(n716), .ZN(n390) );
  AND2_X1 U374 ( .A1(n608), .A2(n353), .ZN(n381) );
  AND2_X1 U375 ( .A1(n567), .A2(n550), .ZN(n353) );
  INV_X1 U376 ( .A(G237), .ZN(n468) );
  XOR2_X1 U377 ( .A(G101), .B(G146), .Z(n408) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n481) );
  XNOR2_X1 U379 ( .A(G134), .B(G122), .ZN(n489) );
  BUF_X2 U380 ( .A(n668), .Z(n351) );
  OR2_X2 U381 ( .A1(n527), .A2(n695), .ZN(n566) );
  XNOR2_X2 U382 ( .A(n388), .B(n592), .ZN(n593) );
  XNOR2_X2 U383 ( .A(n352), .B(KEYINPUT45), .ZN(n743) );
  NAND2_X2 U384 ( .A1(n594), .A2(n593), .ZN(n352) );
  NAND2_X1 U385 ( .A1(n367), .A2(n385), .ZN(n388) );
  NOR2_X2 U386 ( .A1(n394), .A2(n702), .ZN(n530) );
  XNOR2_X2 U387 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X2 U388 ( .A1(n391), .A2(n389), .ZN(n572) );
  XNOR2_X2 U389 ( .A(n759), .B(n406), .ZN(n668) );
  NOR2_X2 U390 ( .A1(n668), .A2(G902), .ZN(n361) );
  XNOR2_X2 U391 ( .A(n370), .B(KEYINPUT33), .ZN(n716) );
  AND2_X4 U392 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  XOR2_X2 U393 ( .A(n470), .B(n469), .Z(n363) );
  XNOR2_X2 U394 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X2 U395 ( .A(n351), .B(n667), .ZN(n669) );
  XNOR2_X2 U396 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U397 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n460) );
  XNOR2_X1 U398 ( .A(KEYINPUT5), .B(KEYINPUT73), .ZN(n411) );
  XNOR2_X1 U399 ( .A(G131), .B(G143), .ZN(n479) );
  XNOR2_X1 U400 ( .A(G146), .B(G104), .ZN(n402) );
  INV_X1 U401 ( .A(G110), .ZN(n399) );
  INV_X1 U402 ( .A(G902), .ZN(n486) );
  XNOR2_X2 U403 ( .A(n636), .B(n635), .ZN(n355) );
  XNOR2_X2 U404 ( .A(n418), .B(n398), .ZN(n759) );
  NAND2_X2 U405 ( .A1(n547), .A2(n356), .ZN(n549) );
  XNOR2_X2 U406 ( .A(n522), .B(n521), .ZN(n547) );
  XNOR2_X2 U407 ( .A(n572), .B(n359), .ZN(n358) );
  NAND2_X2 U408 ( .A1(n674), .A2(n565), .ZN(n373) );
  XNOR2_X2 U409 ( .A(n373), .B(KEYINPUT89), .ZN(n579) );
  INV_X8 U410 ( .A(G953), .ZN(n752) );
  NAND2_X1 U411 ( .A1(n648), .A2(G953), .ZN(n681) );
  BUF_X4 U412 ( .A(G113), .Z(n369) );
  NOR2_X1 U413 ( .A1(n387), .A2(n386), .ZN(n385) );
  AND2_X1 U414 ( .A1(n383), .A2(n591), .ZN(n367) );
  NOR2_X1 U415 ( .A1(n358), .A2(n584), .ZN(n387) );
  XNOR2_X1 U416 ( .A(n560), .B(n559), .ZN(n596) );
  OR2_X1 U417 ( .A1(n558), .A2(n557), .ZN(n560) );
  AND2_X1 U418 ( .A1(n395), .A2(n392), .ZN(n391) );
  BUF_X1 U419 ( .A(n524), .Z(n693) );
  XNOR2_X2 U420 ( .A(KEYINPUT92), .B(G101), .ZN(n400) );
  NAND2_X2 U421 ( .A1(G234), .A2(G237), .ZN(n441) );
  XNOR2_X1 U422 ( .A(KEYINPUT24), .B(KEYINPUT77), .ZN(n427) );
  XOR2_X2 U423 ( .A(G137), .B(KEYINPUT98), .Z(n412) );
  XNOR2_X1 U424 ( .A(G128), .B(KEYINPUT23), .ZN(n428) );
  XNOR2_X2 U425 ( .A(G140), .B(G137), .ZN(n421) );
  XNOR2_X2 U426 ( .A(G116), .B(G107), .ZN(n495) );
  XNOR2_X2 U427 ( .A(KEYINPUT15), .B(G902), .ZN(n467) );
  XNOR2_X2 U428 ( .A(G110), .B(G119), .ZN(n420) );
  XNOR2_X2 U429 ( .A(G146), .B(G125), .ZN(n461) );
  XNOR2_X2 U430 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n426) );
  XNOR2_X2 U431 ( .A(n354), .B(n457), .ZN(n749) );
  XNOR2_X2 U432 ( .A(n483), .B(n456), .ZN(n354) );
  AND2_X1 U433 ( .A1(n584), .A2(KEYINPUT44), .ZN(n384) );
  XOR2_X1 U434 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n490) );
  XNOR2_X1 U435 ( .A(n495), .B(KEYINPUT103), .ZN(n368) );
  XNOR2_X1 U436 ( .A(G134), .B(G131), .ZN(n397) );
  XNOR2_X1 U437 ( .A(n369), .B(G116), .ZN(n407) );
  INV_X1 U438 ( .A(KEYINPUT71), .ZN(n574) );
  NOR2_X1 U439 ( .A1(n584), .A2(KEYINPUT44), .ZN(n386) );
  INV_X1 U440 ( .A(KEYINPUT86), .ZN(n592) );
  XNOR2_X1 U441 ( .A(n478), .B(n365), .ZN(n480) );
  XNOR2_X1 U442 ( .A(n479), .B(n366), .ZN(n365) );
  INV_X1 U443 ( .A(KEYINPUT101), .ZN(n366) );
  INV_X1 U444 ( .A(KEYINPUT106), .ZN(n372) );
  AND2_X1 U445 ( .A1(n393), .A2(n571), .ZN(n392) );
  NAND2_X1 U446 ( .A1(n394), .A2(KEYINPUT34), .ZN(n393) );
  NAND2_X1 U447 ( .A1(n390), .A2(KEYINPUT34), .ZN(n389) );
  NAND2_X1 U448 ( .A1(n375), .A2(n374), .ZN(n760) );
  INV_X1 U449 ( .A(n633), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U451 ( .A(KEYINPUT84), .ZN(n376) );
  XNOR2_X1 U452 ( .A(n542), .B(KEYINPUT39), .ZN(n558) );
  XNOR2_X1 U453 ( .A(n488), .B(n487), .ZN(n544) );
  NAND2_X1 U454 ( .A1(n380), .A2(n379), .ZN(n378) );
  XNOR2_X1 U455 ( .A(n494), .B(n368), .ZN(n496) );
  INV_X1 U456 ( .A(n358), .ZN(n583) );
  NOR2_X1 U457 ( .A1(n710), .A2(n546), .ZN(n356) );
  AND2_X1 U458 ( .A1(n523), .A2(n568), .ZN(n357) );
  INV_X1 U459 ( .A(n760), .ZN(n634) );
  XOR2_X1 U460 ( .A(KEYINPUT83), .B(KEYINPUT35), .Z(n359) );
  AND2_X2 U461 ( .A1(n639), .A2(n634), .ZN(n642) );
  NOR2_X2 U462 ( .A1(n355), .A2(n643), .ZN(n360) );
  NOR2_X1 U463 ( .A1(n355), .A2(n643), .ZN(n676) );
  NOR2_X2 U464 ( .A1(n642), .A2(n641), .ZN(n643) );
  INV_X1 U465 ( .A(n538), .ZN(n380) );
  XNOR2_X1 U466 ( .A(n566), .B(n372), .ZN(n371) );
  NOR2_X1 U467 ( .A1(n629), .A2(n628), .ZN(n630) );
  AND2_X1 U468 ( .A1(n561), .A2(n567), .ZN(n553) );
  XNOR2_X1 U469 ( .A(n362), .B(n363), .ZN(n513) );
  XNOR2_X2 U470 ( .A(n361), .B(G469), .ZN(n538) );
  NOR2_X1 U471 ( .A1(n658), .A2(n640), .ZN(n362) );
  XNOR2_X1 U472 ( .A(n364), .B(n657), .ZN(G60) );
  NAND2_X1 U473 ( .A1(n656), .A2(n681), .ZN(n364) );
  INV_X1 U474 ( .A(n523), .ZN(n394) );
  NAND2_X1 U475 ( .A1(n371), .A2(n506), .ZN(n370) );
  XNOR2_X2 U476 ( .A(n552), .B(KEYINPUT32), .ZN(n565) );
  NAND2_X1 U477 ( .A1(n564), .A2(n563), .ZN(n674) );
  XNOR2_X1 U478 ( .A(n579), .B(KEYINPUT88), .ZN(n573) );
  NAND2_X1 U479 ( .A1(n632), .A2(n631), .ZN(n377) );
  NOR2_X1 U480 ( .A1(n378), .A2(n698), .ZN(n585) );
  NOR2_X1 U481 ( .A1(n378), .A2(n539), .ZN(n541) );
  INV_X1 U482 ( .A(n695), .ZN(n379) );
  NAND2_X1 U483 ( .A1(n381), .A2(n561), .ZN(n552) );
  XNOR2_X2 U484 ( .A(n382), .B(G143), .ZN(n492) );
  XNOR2_X2 U485 ( .A(G128), .B(KEYINPUT78), .ZN(n382) );
  NAND2_X1 U486 ( .A1(n358), .A2(n384), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n716), .A2(n357), .ZN(n395) );
  XNOR2_X2 U488 ( .A(n455), .B(G104), .ZN(n483) );
  AND2_X1 U489 ( .A1(n396), .A2(n614), .ZN(n542) );
  XNOR2_X2 U490 ( .A(n409), .B(G119), .ZN(n456) );
  NOR2_X1 U491 ( .A1(n597), .A2(n537), .ZN(n396) );
  INV_X1 U492 ( .A(KEYINPUT87), .ZN(n584) );
  INV_X1 U493 ( .A(KEYINPUT44), .ZN(n576) );
  XNOR2_X1 U494 ( .A(n575), .B(n574), .ZN(n577) );
  INV_X1 U495 ( .A(KEYINPUT82), .ZN(n637) );
  INV_X1 U496 ( .A(KEYINPUT19), .ZN(n472) );
  INV_X1 U497 ( .A(n421), .ZN(n398) );
  INV_X1 U498 ( .A(KEYINPUT34), .ZN(n568) );
  BUF_X1 U499 ( .A(n676), .Z(n683) );
  XNOR2_X2 U500 ( .A(n492), .B(KEYINPUT4), .ZN(n458) );
  XNOR2_X2 U501 ( .A(n458), .B(n397), .ZN(n418) );
  XNOR2_X1 U502 ( .A(n400), .B(n399), .ZN(n751) );
  XNOR2_X1 U503 ( .A(n751), .B(KEYINPUT70), .ZN(n464) );
  INV_X1 U504 ( .A(n464), .ZN(n405) );
  NAND2_X1 U505 ( .A1(n752), .A2(G227), .ZN(n401) );
  XNOR2_X1 U506 ( .A(n401), .B(G107), .ZN(n403) );
  XNOR2_X1 U507 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U508 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U509 ( .A(n538), .B(KEYINPUT109), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X2 U511 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n409) );
  XNOR2_X1 U512 ( .A(n456), .B(n410), .ZN(n416) );
  XNOR2_X1 U513 ( .A(n412), .B(n411), .ZN(n414) );
  NAND2_X1 U514 ( .A1(n481), .A2(G210), .ZN(n413) );
  XNOR2_X1 U515 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U516 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U517 ( .A(n418), .B(n417), .ZN(n645) );
  OR2_X1 U518 ( .A1(n645), .A2(G902), .ZN(n419) );
  XNOR2_X2 U519 ( .A(n419), .B(G472), .ZN(n698) );
  INV_X1 U520 ( .A(n698), .ZN(n451) );
  XNOR2_X1 U521 ( .A(n420), .B(KEYINPUT95), .ZN(n422) );
  XNOR2_X1 U522 ( .A(n422), .B(n421), .ZN(n425) );
  NAND2_X1 U523 ( .A1(G234), .A2(n752), .ZN(n423) );
  XOR2_X1 U524 ( .A(KEYINPUT8), .B(n423), .Z(n493) );
  NAND2_X1 U525 ( .A1(n493), .A2(G221), .ZN(n424) );
  XNOR2_X1 U526 ( .A(n425), .B(n424), .ZN(n431) );
  XNOR2_X1 U527 ( .A(n461), .B(n426), .ZN(n758) );
  XNOR2_X1 U528 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U529 ( .A(n758), .B(n429), .ZN(n430) );
  XNOR2_X1 U530 ( .A(n431), .B(n430), .ZN(n678) );
  NAND2_X1 U531 ( .A1(n678), .A2(n486), .ZN(n440) );
  NAND2_X1 U532 ( .A1(n467), .A2(G234), .ZN(n433) );
  INV_X1 U533 ( .A(KEYINPUT20), .ZN(n432) );
  XNOR2_X1 U534 ( .A(n433), .B(n432), .ZN(n447) );
  INV_X1 U535 ( .A(G217), .ZN(n434) );
  OR2_X1 U536 ( .A1(n447), .A2(n434), .ZN(n438) );
  XNOR2_X1 U537 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n436) );
  XNOR2_X1 U538 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n435) );
  XNOR2_X1 U539 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U540 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U541 ( .A(n440), .B(n439), .ZN(n524) );
  XNOR2_X1 U542 ( .A(n441), .B(KEYINPUT94), .ZN(n442) );
  XNOR2_X1 U543 ( .A(KEYINPUT14), .B(n442), .ZN(n444) );
  AND2_X1 U544 ( .A1(n444), .A2(G953), .ZN(n443) );
  NAND2_X1 U545 ( .A1(G902), .A2(n443), .ZN(n516) );
  OR2_X1 U546 ( .A1(n516), .A2(G900), .ZN(n445) );
  NAND2_X1 U547 ( .A1(G952), .A2(n444), .ZN(n723) );
  OR2_X1 U548 ( .A1(n723), .A2(G953), .ZN(n517) );
  AND2_X1 U549 ( .A1(n445), .A2(n517), .ZN(n539) );
  INV_X1 U550 ( .A(G221), .ZN(n446) );
  OR2_X1 U551 ( .A1(n447), .A2(n446), .ZN(n448) );
  XNOR2_X1 U552 ( .A(n448), .B(KEYINPUT21), .ZN(n546) );
  NOR2_X1 U553 ( .A1(n539), .A2(n546), .ZN(n449) );
  XOR2_X1 U554 ( .A(KEYINPUT68), .B(n449), .Z(n450) );
  OR2_X1 U555 ( .A1(n693), .A2(n450), .ZN(n505) );
  NOR2_X1 U556 ( .A1(n451), .A2(n505), .ZN(n452) );
  XNOR2_X1 U557 ( .A(n452), .B(KEYINPUT28), .ZN(n453) );
  NAND2_X1 U558 ( .A1(n454), .A2(n453), .ZN(n599) );
  XNOR2_X2 U559 ( .A(G122), .B(G113), .ZN(n455) );
  XNOR2_X1 U560 ( .A(n495), .B(KEYINPUT16), .ZN(n457) );
  XNOR2_X1 U561 ( .A(n749), .B(n458), .ZN(n466) );
  NAND2_X1 U562 ( .A1(n752), .A2(G224), .ZN(n459) );
  XNOR2_X1 U563 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U565 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U566 ( .A(n466), .B(n465), .ZN(n658) );
  INV_X1 U567 ( .A(n467), .ZN(n640) );
  NAND2_X1 U568 ( .A1(n486), .A2(n468), .ZN(n471) );
  NAND2_X1 U569 ( .A1(n471), .A2(G210), .ZN(n470) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n469) );
  AND2_X1 U571 ( .A1(n471), .A2(G214), .ZN(n509) );
  NOR2_X2 U572 ( .A1(n513), .A2(n509), .ZN(n473) );
  XNOR2_X1 U573 ( .A(n473), .B(n472), .ZN(n520) );
  BUF_X1 U574 ( .A(n520), .Z(n474) );
  INV_X1 U575 ( .A(n474), .ZN(n475) );
  OR2_X1 U576 ( .A1(n599), .A2(n475), .ZN(n618) );
  INV_X1 U577 ( .A(n618), .ZN(n621) );
  XOR2_X1 U578 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n477) );
  XNOR2_X1 U579 ( .A(G140), .B(KEYINPUT12), .ZN(n476) );
  XNOR2_X1 U580 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U581 ( .A(n480), .B(n758), .ZN(n485) );
  NAND2_X1 U582 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U583 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n485), .B(n484), .ZN(n653) );
  NAND2_X1 U585 ( .A1(n653), .A2(n486), .ZN(n488) );
  XNOR2_X1 U586 ( .A(KEYINPUT13), .B(G475), .ZN(n487) );
  INV_X1 U587 ( .A(n544), .ZN(n569) );
  XNOR2_X1 U588 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n492), .B(n491), .ZN(n497) );
  NAND2_X1 U590 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n497), .B(n496), .ZN(n684) );
  NOR2_X1 U592 ( .A1(G902), .A2(n684), .ZN(n498) );
  XNOR2_X1 U593 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n499), .B(G478), .ZN(n545) );
  AND2_X1 U595 ( .A1(n569), .A2(n545), .ZN(n733) );
  NAND2_X1 U596 ( .A1(n621), .A2(n733), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n500), .B(G146), .ZN(G48) );
  XOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n502) );
  XNOR2_X1 U599 ( .A(G128), .B(KEYINPUT29), .ZN(n501) );
  XNOR2_X1 U600 ( .A(n502), .B(n501), .ZN(n504) );
  INV_X1 U601 ( .A(n545), .ZN(n570) );
  AND2_X1 U602 ( .A1(n570), .A2(n544), .ZN(n735) );
  NAND2_X1 U603 ( .A1(n621), .A2(n735), .ZN(n503) );
  XOR2_X1 U604 ( .A(n504), .B(n503), .Z(G30) );
  INV_X1 U605 ( .A(n733), .ZN(n557) );
  NOR2_X1 U606 ( .A1(n557), .A2(n505), .ZN(n507) );
  XNOR2_X1 U607 ( .A(n698), .B(KEYINPUT6), .ZN(n567) );
  INV_X1 U608 ( .A(n567), .ZN(n506) );
  NAND2_X1 U609 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U610 ( .A(n508), .B(KEYINPUT107), .ZN(n510) );
  INV_X1 U611 ( .A(n509), .ZN(n706) );
  AND2_X1 U612 ( .A1(n510), .A2(n706), .ZN(n605) );
  XNOR2_X1 U613 ( .A(KEYINPUT64), .B(KEYINPUT1), .ZN(n511) );
  XNOR2_X2 U614 ( .A(n538), .B(n511), .ZN(n527) );
  NAND2_X1 U615 ( .A1(n605), .A2(n527), .ZN(n512) );
  XNOR2_X1 U616 ( .A(n512), .B(KEYINPUT43), .ZN(n515) );
  BUF_X1 U617 ( .A(n513), .Z(n514) );
  NAND2_X1 U618 ( .A1(n515), .A2(n514), .ZN(n631) );
  XNOR2_X1 U619 ( .A(n631), .B(G140), .ZN(G42) );
  OR2_X1 U620 ( .A1(n516), .A2(G898), .ZN(n518) );
  NAND2_X1 U621 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U622 ( .A1(n520), .A2(n519), .ZN(n522) );
  INV_X1 U623 ( .A(KEYINPUT0), .ZN(n521) );
  BUF_X1 U624 ( .A(n547), .Z(n523) );
  INV_X1 U625 ( .A(n546), .ZN(n692) );
  NAND2_X1 U626 ( .A1(n524), .A2(n692), .ZN(n526) );
  INV_X1 U627 ( .A(KEYINPUT65), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n526), .B(n525), .ZN(n695) );
  INV_X1 U629 ( .A(n566), .ZN(n528) );
  NAND2_X1 U630 ( .A1(n528), .A2(n698), .ZN(n702) );
  XNOR2_X1 U631 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n529) );
  XNOR2_X1 U632 ( .A(n530), .B(n529), .ZN(n586) );
  NAND2_X1 U633 ( .A1(n586), .A2(n735), .ZN(n531) );
  XNOR2_X1 U634 ( .A(n531), .B(G116), .ZN(G18) );
  NAND2_X1 U635 ( .A1(n586), .A2(n733), .ZN(n532) );
  XNOR2_X1 U636 ( .A(n532), .B(n369), .ZN(G15) );
  INV_X1 U637 ( .A(KEYINPUT38), .ZN(n533) );
  XNOR2_X1 U638 ( .A(n514), .B(n533), .ZN(n597) );
  NAND2_X1 U639 ( .A1(n698), .A2(n706), .ZN(n536) );
  INV_X1 U640 ( .A(KEYINPUT108), .ZN(n534) );
  XNOR2_X1 U641 ( .A(n534), .B(KEYINPUT30), .ZN(n535) );
  XNOR2_X1 U642 ( .A(n536), .B(n535), .ZN(n612) );
  INV_X1 U643 ( .A(n612), .ZN(n537) );
  INV_X1 U644 ( .A(KEYINPUT75), .ZN(n540) );
  XNOR2_X1 U645 ( .A(n541), .B(n540), .ZN(n614) );
  INV_X1 U646 ( .A(n558), .ZN(n543) );
  AND2_X1 U647 ( .A1(n543), .A2(n735), .ZN(n633) );
  XOR2_X1 U648 ( .A(G134), .B(n633), .Z(G36) );
  NAND2_X1 U649 ( .A1(n545), .A2(n544), .ZN(n710) );
  INV_X1 U650 ( .A(KEYINPUT22), .ZN(n548) );
  XNOR2_X2 U651 ( .A(n549), .B(n548), .ZN(n561) );
  XNOR2_X1 U652 ( .A(n527), .B(KEYINPUT91), .ZN(n608) );
  INV_X1 U653 ( .A(n693), .ZN(n550) );
  XNOR2_X1 U654 ( .A(n565), .B(G119), .ZN(G21) );
  INV_X1 U655 ( .A(n553), .ZN(n554) );
  XOR2_X1 U656 ( .A(n554), .B(KEYINPUT85), .Z(n556) );
  NAND2_X1 U657 ( .A1(n527), .A2(n693), .ZN(n555) );
  NOR2_X1 U658 ( .A1(n556), .A2(n555), .ZN(n589) );
  XOR2_X1 U659 ( .A(G101), .B(n589), .Z(G3) );
  INV_X1 U660 ( .A(KEYINPUT40), .ZN(n559) );
  XOR2_X1 U661 ( .A(G131), .B(n596), .Z(G33) );
  NAND2_X1 U662 ( .A1(n561), .A2(n527), .ZN(n562) );
  XNOR2_X1 U663 ( .A(n562), .B(KEYINPUT105), .ZN(n564) );
  NOR2_X1 U664 ( .A1(n698), .A2(n693), .ZN(n563) );
  NAND2_X1 U665 ( .A1(n570), .A2(n569), .ZN(n610) );
  INV_X1 U666 ( .A(n610), .ZN(n571) );
  NAND2_X1 U667 ( .A1(n573), .A2(n583), .ZN(n575) );
  NAND2_X1 U668 ( .A1(n577), .A2(n576), .ZN(n582) );
  NOR2_X1 U669 ( .A1(n576), .A2(KEYINPUT71), .ZN(n578) );
  AND2_X1 U670 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U671 ( .A(n580), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n594) );
  AND2_X1 U673 ( .A1(n523), .A2(n585), .ZN(n736) );
  NOR2_X1 U674 ( .A1(n586), .A2(n736), .ZN(n587) );
  XNOR2_X1 U675 ( .A(n587), .B(KEYINPUT100), .ZN(n588) );
  NOR2_X1 U676 ( .A1(n735), .A2(n733), .ZN(n712) );
  NOR2_X1 U677 ( .A1(n588), .A2(n712), .ZN(n590) );
  NOR2_X1 U678 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U679 ( .A(n596), .ZN(n602) );
  INV_X1 U680 ( .A(n597), .ZN(n707) );
  NAND2_X1 U681 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U682 ( .A1(n710), .A2(n711), .ZN(n598) );
  XNOR2_X1 U683 ( .A(n598), .B(KEYINPUT41), .ZN(n725) );
  NOR2_X1 U684 ( .A1(n725), .A2(n599), .ZN(n600) );
  XNOR2_X1 U685 ( .A(n600), .B(KEYINPUT42), .ZN(n769) );
  INV_X1 U686 ( .A(n769), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U688 ( .A(n603), .B(KEYINPUT46), .ZN(n629) );
  INV_X1 U689 ( .A(n514), .ZN(n604) );
  NAND2_X1 U690 ( .A1(n605), .A2(n604), .ZN(n607) );
  INV_X1 U691 ( .A(KEYINPUT36), .ZN(n606) );
  XNOR2_X1 U692 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n609), .A2(n608), .ZN(n741) );
  NOR2_X1 U694 ( .A1(n610), .A2(n514), .ZN(n611) );
  AND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  AND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n740) );
  XNOR2_X1 U697 ( .A(n740), .B(KEYINPUT81), .ZN(n615) );
  AND2_X1 U698 ( .A1(n741), .A2(n615), .ZN(n627) );
  INV_X1 U699 ( .A(KEYINPUT66), .ZN(n616) );
  OR2_X1 U700 ( .A1(n712), .A2(n616), .ZN(n617) );
  NOR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT47), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(KEYINPUT72), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n712), .A2(KEYINPUT72), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n622) );
  OR2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT48), .ZN(n632) );
  AND2_X1 U710 ( .A1(n743), .A2(n634), .ZN(n688) );
  NAND2_X1 U711 ( .A1(n688), .A2(KEYINPUT2), .ZN(n636) );
  INV_X1 U712 ( .A(KEYINPUT74), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n743), .A2(n640), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n360), .A2(G472), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n644) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n649) );
  INV_X1 U718 ( .A(G952), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n681), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(G57) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n657) );
  NAND2_X1 U723 ( .A1(n360), .A2(G475), .ZN(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n676), .A2(G210), .ZN(n662) );
  BUF_X1 U727 ( .A(n658), .Z(n660) );
  XNOR2_X1 U728 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n663), .A2(n681), .ZN(n665) );
  INV_X1 U731 ( .A(KEYINPUT56), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(n664), .ZN(G51) );
  INV_X1 U733 ( .A(KEYINPUT120), .ZN(n673) );
  NAND2_X1 U734 ( .A1(n360), .A2(G469), .ZN(n670) );
  XNOR2_X1 U735 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n666) );
  XOR2_X1 U736 ( .A(n666), .B(KEYINPUT58), .Z(n667) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n671), .A2(n681), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(n673), .ZN(G54) );
  BUF_X1 U740 ( .A(n674), .Z(n675) );
  XNOR2_X1 U741 ( .A(n675), .B(G110), .ZN(G12) );
  XNOR2_X1 U742 ( .A(n583), .B(G122), .ZN(G24) );
  NAND2_X1 U743 ( .A1(n683), .A2(G217), .ZN(n680) );
  XNOR2_X1 U744 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(n682) );
  INV_X1 U747 ( .A(n681), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n682), .A2(n686), .ZN(G66) );
  NAND2_X1 U749 ( .A1(n683), .A2(G478), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(n684), .ZN(n687) );
  NOR2_X1 U751 ( .A1(n687), .A2(n686), .ZN(G63) );
  XNOR2_X1 U752 ( .A(KEYINPUT2), .B(KEYINPUT80), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n688), .A2(n689), .ZN(n690) );
  XOR2_X1 U754 ( .A(KEYINPUT79), .B(n690), .Z(n691) );
  NOR2_X1 U755 ( .A1(n691), .A2(n355), .ZN(n731) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U757 ( .A(n694), .B(KEYINPUT49), .ZN(n700) );
  NAND2_X1 U758 ( .A1(n527), .A2(n695), .ZN(n696) );
  XOR2_X1 U759 ( .A(KEYINPUT50), .B(n696), .Z(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U763 ( .A(n703), .B(KEYINPUT51), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n725), .A2(n704), .ZN(n705) );
  XOR2_X1 U765 ( .A(KEYINPUT113), .B(n705), .Z(n719) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n708), .B(KEYINPUT114), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U771 ( .A(KEYINPUT115), .B(n715), .Z(n717) );
  NOR2_X1 U772 ( .A1(n717), .A2(n390), .ZN(n718) );
  NOR2_X1 U773 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U774 ( .A(KEYINPUT116), .B(n720), .Z(n721) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n721), .Z(n722) );
  NOR2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U777 ( .A(KEYINPUT117), .B(n724), .Z(n727) );
  NOR2_X1 U778 ( .A1(n725), .A2(n390), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(KEYINPUT118), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(n752), .ZN(n730) );
  NOR2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n732), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U784 ( .A1(n736), .A2(n733), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n734), .B(G104), .ZN(G6) );
  XOR2_X1 U786 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n738) );
  NAND2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(G107), .B(n739), .ZN(G9) );
  XOR2_X1 U790 ( .A(G143), .B(n740), .Z(G45) );
  XOR2_X1 U791 ( .A(G125), .B(n741), .Z(n742) );
  XNOR2_X1 U792 ( .A(n742), .B(KEYINPUT37), .ZN(G27) );
  BUF_X1 U793 ( .A(n743), .Z(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(n752), .ZN(n748) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U797 ( .A1(n746), .A2(G898), .ZN(n747) );
  NAND2_X1 U798 ( .A1(n748), .A2(n747), .ZN(n756) );
  BUF_X1 U799 ( .A(n749), .Z(n750) );
  XNOR2_X1 U800 ( .A(n750), .B(n751), .ZN(n754) );
  NOR2_X1 U801 ( .A1(n752), .A2(G898), .ZN(n753) );
  NOR2_X1 U802 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U804 ( .A(KEYINPUT124), .B(n757), .ZN(G69) );
  XNOR2_X1 U805 ( .A(n759), .B(n758), .ZN(n763) );
  XNOR2_X1 U806 ( .A(n760), .B(n763), .ZN(n761) );
  NOR2_X1 U807 ( .A1(n761), .A2(G953), .ZN(n762) );
  XNOR2_X1 U808 ( .A(KEYINPUT125), .B(n762), .ZN(n768) );
  XOR2_X1 U809 ( .A(G227), .B(n763), .Z(n764) );
  NAND2_X1 U810 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U811 ( .A1(G953), .A2(n765), .ZN(n766) );
  XNOR2_X1 U812 ( .A(KEYINPUT126), .B(n766), .ZN(n767) );
  NAND2_X1 U813 ( .A1(n768), .A2(n767), .ZN(G72) );
  XOR2_X1 U814 ( .A(G137), .B(n769), .Z(G39) );
endmodule

