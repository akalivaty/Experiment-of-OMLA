

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n656), .A2(n655), .ZN(n657) );
  OR2_X1 U553 ( .A1(n549), .A2(G2105), .ZN(n550) );
  NAND2_X1 U554 ( .A1(n769), .A2(n768), .ZN(n771) );
  NOR2_X2 U555 ( .A1(G2104), .A2(n542), .ZN(n551) );
  INV_X1 U556 ( .A(KEYINPUT99), .ZN(n621) );
  XNOR2_X1 U557 ( .A(n622), .B(n621), .ZN(n627) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n670) );
  XNOR2_X1 U559 ( .A(n670), .B(KEYINPUT102), .ZN(n671) );
  XNOR2_X1 U560 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U561 ( .A1(n674), .A2(n673), .ZN(n686) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n714), .ZN(n688) );
  NOR2_X1 U563 ( .A1(G651), .A2(n586), .ZN(n814) );
  INV_X1 U564 ( .A(KEYINPUT40), .ZN(n770) );
  NOR2_X1 U565 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U566 ( .A(n561), .B(n560), .ZN(G160) );
  XNOR2_X1 U567 ( .A(G543), .B(KEYINPUT0), .ZN(n522) );
  XNOR2_X1 U568 ( .A(n522), .B(KEYINPUT69), .ZN(n586) );
  NAND2_X1 U569 ( .A1(G51), .A2(n814), .ZN(n525) );
  INV_X1 U570 ( .A(G651), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G543), .A2(n529), .ZN(n523) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n523), .Z(n810) );
  NAND2_X1 U573 ( .A1(n810), .A2(G63), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n526), .B(KEYINPUT6), .ZN(n527) );
  XOR2_X1 U576 ( .A(KEYINPUT81), .B(n527), .Z(n535) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n806) );
  NAND2_X1 U578 ( .A1(n806), .A2(G89), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  NOR2_X1 U580 ( .A1(n586), .A2(n529), .ZN(n807) );
  NAND2_X1 U581 ( .A1(G76), .A2(n807), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U583 ( .A(n532), .B(KEYINPUT80), .Z(n533) );
  XNOR2_X1 U584 ( .A(KEYINPUT5), .B(n533), .ZN(n534) );
  NOR2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U586 ( .A(KEYINPUT7), .B(n536), .Z(G168) );
  XOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U588 ( .A(KEYINPUT89), .ZN(n548) );
  INV_X1 U589 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U590 ( .A1(G126), .A2(n551), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XNOR2_X1 U592 ( .A(n537), .B(KEYINPUT67), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT68), .B(KEYINPUT17), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n539), .B(n538), .ZN(n555) );
  NAND2_X1 U595 ( .A1(G138), .A2(n555), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n546) );
  AND2_X1 U597 ( .A1(n542), .A2(G2104), .ZN(n897) );
  NAND2_X1 U598 ( .A1(G102), .A2(n897), .ZN(n544) );
  AND2_X1 U599 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U600 ( .A1(G114), .A2(n901), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n548), .B(n547), .ZN(G164) );
  NAND2_X1 U604 ( .A1(G101), .A2(G2104), .ZN(n549) );
  XOR2_X1 U605 ( .A(n550), .B(KEYINPUT23), .Z(n553) );
  NAND2_X1 U606 ( .A1(n551), .A2(G125), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U608 ( .A(n554), .B(KEYINPUT66), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G137), .A2(n555), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n901), .A2(G113), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U612 ( .A(KEYINPUT65), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n814), .A2(G53), .ZN(n568) );
  NAND2_X1 U614 ( .A1(G91), .A2(n806), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G65), .A2(n810), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n807), .A2(G78), .ZN(n564) );
  XOR2_X1 U618 ( .A(KEYINPUT74), .B(n564), .Z(n565) );
  NOR2_X1 U619 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U620 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U621 ( .A(KEYINPUT75), .B(n569), .Z(G299) );
  NAND2_X1 U622 ( .A1(n806), .A2(G90), .ZN(n570) );
  XNOR2_X1 U623 ( .A(n570), .B(KEYINPUT72), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G77), .A2(n807), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n573) );
  XNOR2_X1 U627 ( .A(n574), .B(n573), .ZN(n578) );
  NAND2_X1 U628 ( .A1(G64), .A2(n810), .ZN(n576) );
  NAND2_X1 U629 ( .A1(G52), .A2(n814), .ZN(n575) );
  AND2_X1 U630 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n578), .A2(n577), .ZN(G301) );
  NAND2_X1 U632 ( .A1(G75), .A2(n807), .ZN(n580) );
  NAND2_X1 U633 ( .A1(G50), .A2(n814), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U635 ( .A1(G88), .A2(n806), .ZN(n582) );
  NAND2_X1 U636 ( .A1(G62), .A2(n810), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U638 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U639 ( .A(n585), .B(KEYINPUT85), .Z(G166) );
  INV_X1 U640 ( .A(G166), .ZN(G303) );
  NAND2_X1 U641 ( .A1(G49), .A2(n814), .ZN(n588) );
  NAND2_X1 U642 ( .A1(G87), .A2(n586), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U644 ( .A1(n810), .A2(n589), .ZN(n591) );
  NAND2_X1 U645 ( .A1(G651), .A2(G74), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n591), .A2(n590), .ZN(G288) );
  NAND2_X1 U647 ( .A1(G86), .A2(n806), .ZN(n593) );
  NAND2_X1 U648 ( .A1(G61), .A2(n810), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U650 ( .A1(n807), .A2(G73), .ZN(n594) );
  XOR2_X1 U651 ( .A(KEYINPUT2), .B(n594), .Z(n595) );
  NOR2_X1 U652 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U653 ( .A1(n814), .A2(G48), .ZN(n597) );
  NAND2_X1 U654 ( .A1(n598), .A2(n597), .ZN(G305) );
  NAND2_X1 U655 ( .A1(n814), .A2(G47), .ZN(n605) );
  NAND2_X1 U656 ( .A1(G85), .A2(n806), .ZN(n600) );
  NAND2_X1 U657 ( .A1(G72), .A2(n807), .ZN(n599) );
  NAND2_X1 U658 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U659 ( .A1(n810), .A2(G60), .ZN(n601) );
  XOR2_X1 U660 ( .A(KEYINPUT70), .B(n601), .Z(n602) );
  NOR2_X1 U661 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U662 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U663 ( .A(KEYINPUT71), .B(n606), .Z(G290) );
  NOR2_X1 U664 ( .A1(G164), .A2(G1384), .ZN(n754) );
  INV_X1 U665 ( .A(n754), .ZN(n608) );
  NAND2_X1 U666 ( .A1(G40), .A2(G160), .ZN(n607) );
  XNOR2_X1 U667 ( .A(n607), .B(KEYINPUT90), .ZN(n755) );
  NOR2_X2 U668 ( .A1(n608), .A2(n755), .ZN(n623) );
  INV_X2 U669 ( .A(n623), .ZN(n675) );
  NAND2_X1 U670 ( .A1(G8), .A2(n675), .ZN(n714) );
  NAND2_X1 U671 ( .A1(n806), .A2(G92), .ZN(n609) );
  XOR2_X1 U672 ( .A(KEYINPUT77), .B(n609), .Z(n611) );
  NAND2_X1 U673 ( .A1(n810), .A2(G66), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U675 ( .A(KEYINPUT78), .B(n612), .ZN(n616) );
  NAND2_X1 U676 ( .A1(G79), .A2(n807), .ZN(n614) );
  NAND2_X1 U677 ( .A1(G54), .A2(n814), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U679 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U680 ( .A(KEYINPUT15), .B(n617), .Z(n618) );
  XOR2_X1 U681 ( .A(KEYINPUT79), .B(n618), .Z(n962) );
  INV_X1 U682 ( .A(n962), .ZN(n792) );
  NAND2_X1 U683 ( .A1(G1348), .A2(n675), .ZN(n620) );
  NAND2_X1 U684 ( .A1(n623), .A2(G2067), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n620), .A2(n619), .ZN(n630) );
  NOR2_X1 U686 ( .A1(n792), .A2(n630), .ZN(n629) );
  NAND2_X1 U687 ( .A1(G1956), .A2(n675), .ZN(n622) );
  XOR2_X1 U688 ( .A(KEYINPUT27), .B(KEYINPUT98), .Z(n625) );
  NAND2_X1 U689 ( .A1(G2072), .A2(n623), .ZN(n624) );
  XNOR2_X1 U690 ( .A(n625), .B(n624), .ZN(n626) );
  NAND2_X1 U691 ( .A1(n627), .A2(n626), .ZN(n653) );
  NOR2_X1 U692 ( .A1(n653), .A2(G299), .ZN(n628) );
  NOR2_X1 U693 ( .A1(n629), .A2(n628), .ZN(n651) );
  NAND2_X1 U694 ( .A1(n630), .A2(n792), .ZN(n649) );
  NAND2_X1 U695 ( .A1(n806), .A2(G81), .ZN(n631) );
  XNOR2_X1 U696 ( .A(n631), .B(KEYINPUT12), .ZN(n633) );
  NAND2_X1 U697 ( .A1(G68), .A2(n807), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U699 ( .A(n634), .B(KEYINPUT13), .ZN(n636) );
  NAND2_X1 U700 ( .A1(G43), .A2(n814), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U702 ( .A1(n810), .A2(G56), .ZN(n637) );
  XOR2_X1 U703 ( .A(KEYINPUT14), .B(n637), .Z(n638) );
  NOR2_X1 U704 ( .A1(n639), .A2(n638), .ZN(n955) );
  XNOR2_X1 U705 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n642) );
  OR2_X1 U706 ( .A1(n642), .A2(G1996), .ZN(n640) );
  NAND2_X1 U707 ( .A1(n955), .A2(n640), .ZN(n647) );
  INV_X1 U708 ( .A(G1341), .ZN(n956) );
  NAND2_X1 U709 ( .A1(n956), .A2(n642), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n641), .A2(n675), .ZN(n645) );
  INV_X1 U711 ( .A(G1996), .ZN(n870) );
  NOR2_X1 U712 ( .A1(n675), .A2(n870), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  AND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(KEYINPUT100), .B(n652), .ZN(n656) );
  NAND2_X1 U719 ( .A1(G299), .A2(n653), .ZN(n654) );
  XOR2_X1 U720 ( .A(KEYINPUT28), .B(n654), .Z(n655) );
  XNOR2_X1 U721 ( .A(n657), .B(KEYINPUT29), .ZN(n662) );
  XOR2_X1 U722 ( .A(KEYINPUT96), .B(G1961), .Z(n926) );
  NAND2_X1 U723 ( .A1(n926), .A2(n675), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n658), .B(KEYINPUT97), .ZN(n660) );
  XOR2_X1 U725 ( .A(G2078), .B(KEYINPUT25), .Z(n1014) );
  NOR2_X1 U726 ( .A1(n675), .A2(n1014), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n663) );
  OR2_X1 U728 ( .A1(G301), .A2(n663), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n674) );
  NAND2_X1 U730 ( .A1(n663), .A2(G301), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(KEYINPUT101), .ZN(n669) );
  NOR2_X1 U732 ( .A1(G2084), .A2(n675), .ZN(n685) );
  NOR2_X1 U733 ( .A1(n688), .A2(n685), .ZN(n665) );
  NAND2_X1 U734 ( .A1(G8), .A2(n665), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(KEYINPUT30), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n667), .A2(G168), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n686), .A2(G286), .ZN(n681) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n714), .ZN(n677) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n675), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n678), .A2(G303), .ZN(n679) );
  XOR2_X1 U743 ( .A(KEYINPUT103), .B(n679), .Z(n680) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n682), .B(KEYINPUT104), .ZN(n683) );
  NAND2_X1 U746 ( .A1(n683), .A2(G8), .ZN(n684) );
  XNOR2_X1 U747 ( .A(n684), .B(KEYINPUT32), .ZN(n709) );
  NAND2_X1 U748 ( .A1(G8), .A2(n685), .ZN(n690) );
  INV_X1 U749 ( .A(n686), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n710) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n951) );
  AND2_X1 U753 ( .A1(n710), .A2(n951), .ZN(n691) );
  NAND2_X1 U754 ( .A1(n709), .A2(n691), .ZN(n697) );
  INV_X1 U755 ( .A(n951), .ZN(n695) );
  NOR2_X1 U756 ( .A1(G288), .A2(G1976), .ZN(n692) );
  XOR2_X1 U757 ( .A(n692), .B(KEYINPUT105), .Z(n972) );
  NOR2_X1 U758 ( .A1(G1971), .A2(G303), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n972), .A2(n693), .ZN(n694) );
  OR2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  AND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n714), .A2(n698), .ZN(n699) );
  NOR2_X1 U763 ( .A1(KEYINPUT33), .A2(n699), .ZN(n704) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n959) );
  INV_X1 U765 ( .A(n972), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n714), .A2(n700), .ZN(n701) );
  NAND2_X1 U767 ( .A1(KEYINPUT33), .A2(n701), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n959), .A2(n702), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XOR2_X1 U771 ( .A(n705), .B(KEYINPUT24), .Z(n706) );
  NOR2_X1 U772 ( .A1(n714), .A2(n706), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n760) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U775 ( .A1(G2090), .A2(G303), .ZN(n711) );
  NAND2_X1 U776 ( .A1(G8), .A2(n711), .ZN(n712) );
  NAND2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n715) );
  NAND2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n758) );
  NAND2_X1 U779 ( .A1(G104), .A2(n897), .ZN(n717) );
  BUF_X1 U780 ( .A(n555), .Z(n898) );
  NAND2_X1 U781 ( .A1(G140), .A2(n898), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n718), .ZN(n723) );
  NAND2_X1 U784 ( .A1(G128), .A2(n551), .ZN(n720) );
  NAND2_X1 U785 ( .A1(G116), .A2(n901), .ZN(n719) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U787 ( .A(n721), .B(KEYINPUT35), .Z(n722) );
  NOR2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U789 ( .A(KEYINPUT36), .B(n724), .Z(n725) );
  XOR2_X1 U790 ( .A(KEYINPUT92), .B(n725), .Z(n913) );
  XNOR2_X1 U791 ( .A(G2067), .B(KEYINPUT37), .ZN(n726) );
  XOR2_X1 U792 ( .A(n726), .B(KEYINPUT91), .Z(n752) );
  OR2_X1 U793 ( .A1(n913), .A2(n752), .ZN(n727) );
  XNOR2_X1 U794 ( .A(n727), .B(KEYINPUT93), .ZN(n763) );
  NAND2_X1 U795 ( .A1(G129), .A2(n551), .ZN(n729) );
  NAND2_X1 U796 ( .A1(G141), .A2(n898), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U798 ( .A1(n897), .A2(G105), .ZN(n730) );
  XOR2_X1 U799 ( .A(KEYINPUT38), .B(n730), .Z(n731) );
  NOR2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U801 ( .A1(n901), .A2(G117), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n910) );
  NOR2_X1 U803 ( .A1(G1996), .A2(n910), .ZN(n981) );
  NOR2_X1 U804 ( .A1(G1986), .A2(G290), .ZN(n744) );
  NAND2_X1 U805 ( .A1(G119), .A2(n551), .ZN(n736) );
  NAND2_X1 U806 ( .A1(G107), .A2(n901), .ZN(n735) );
  NAND2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U808 ( .A(KEYINPUT94), .B(n737), .ZN(n740) );
  NAND2_X1 U809 ( .A1(G131), .A2(n898), .ZN(n738) );
  XNOR2_X1 U810 ( .A(KEYINPUT95), .B(n738), .ZN(n739) );
  NOR2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U812 ( .A1(n897), .A2(G95), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n742), .A2(n741), .ZN(n887) );
  NOR2_X1 U814 ( .A1(n887), .A2(G1991), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(KEYINPUT106), .ZN(n992) );
  NOR2_X1 U816 ( .A1(n744), .A2(n992), .ZN(n747) );
  NAND2_X1 U817 ( .A1(G1996), .A2(n910), .ZN(n746) );
  NAND2_X1 U818 ( .A1(G1991), .A2(n887), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n762) );
  NOR2_X1 U820 ( .A1(n747), .A2(n762), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n981), .A2(n748), .ZN(n749) );
  XOR2_X1 U822 ( .A(KEYINPUT39), .B(n749), .Z(n750) );
  NOR2_X1 U823 ( .A1(n763), .A2(n750), .ZN(n751) );
  XNOR2_X1 U824 ( .A(KEYINPUT107), .B(n751), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n913), .A2(n752), .ZN(n990) );
  NAND2_X1 U826 ( .A1(n753), .A2(n990), .ZN(n756) );
  NOR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n765) );
  NAND2_X1 U828 ( .A1(n756), .A2(n765), .ZN(n757) );
  XNOR2_X1 U829 ( .A(n757), .B(KEYINPUT108), .ZN(n761) );
  AND2_X1 U830 ( .A1(n758), .A2(n761), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n760), .A2(n759), .ZN(n769) );
  INV_X1 U832 ( .A(n761), .ZN(n767) );
  NOR2_X1 U833 ( .A1(n763), .A2(n762), .ZN(n998) );
  XOR2_X1 U834 ( .A(G1986), .B(G290), .Z(n957) );
  NAND2_X1 U835 ( .A1(n998), .A2(n957), .ZN(n764) );
  NAND2_X1 U836 ( .A1(n765), .A2(n764), .ZN(n766) );
  OR2_X1 U837 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U838 ( .A(n771), .B(n770), .ZN(G329) );
  XNOR2_X1 U839 ( .A(G2451), .B(G2427), .ZN(n781) );
  XOR2_X1 U840 ( .A(KEYINPUT109), .B(G2443), .Z(n773) );
  XNOR2_X1 U841 ( .A(G2435), .B(G2438), .ZN(n772) );
  XNOR2_X1 U842 ( .A(n773), .B(n772), .ZN(n777) );
  XOR2_X1 U843 ( .A(G2454), .B(G2430), .Z(n775) );
  XOR2_X1 U844 ( .A(G1348), .B(n956), .Z(n774) );
  XNOR2_X1 U845 ( .A(n775), .B(n774), .ZN(n776) );
  XOR2_X1 U846 ( .A(n777), .B(n776), .Z(n779) );
  XNOR2_X1 U847 ( .A(G2446), .B(KEYINPUT110), .ZN(n778) );
  XNOR2_X1 U848 ( .A(n779), .B(n778), .ZN(n780) );
  XNOR2_X1 U849 ( .A(n781), .B(n780), .ZN(n782) );
  AND2_X1 U850 ( .A1(n782), .A2(G14), .ZN(G401) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U852 ( .A(G57), .ZN(G237) );
  NAND2_X1 U853 ( .A1(G7), .A2(G661), .ZN(n783) );
  XNOR2_X1 U854 ( .A(n783), .B(KEYINPUT10), .ZN(n784) );
  XOR2_X1 U855 ( .A(KEYINPUT76), .B(n784), .Z(n925) );
  NAND2_X1 U856 ( .A1(n925), .A2(G567), .ZN(n785) );
  XOR2_X1 U857 ( .A(KEYINPUT11), .B(n785), .Z(G234) );
  NAND2_X1 U858 ( .A1(n955), .A2(G860), .ZN(G153) );
  NAND2_X1 U859 ( .A1(G868), .A2(G301), .ZN(n787) );
  INV_X1 U860 ( .A(G868), .ZN(n829) );
  NAND2_X1 U861 ( .A1(n792), .A2(n829), .ZN(n786) );
  NAND2_X1 U862 ( .A1(n787), .A2(n786), .ZN(G284) );
  NOR2_X1 U863 ( .A1(G868), .A2(G299), .ZN(n788) );
  XNOR2_X1 U864 ( .A(n788), .B(KEYINPUT82), .ZN(n790) );
  NOR2_X1 U865 ( .A1(n829), .A2(G286), .ZN(n789) );
  NOR2_X1 U866 ( .A1(n790), .A2(n789), .ZN(G297) );
  INV_X1 U867 ( .A(G860), .ZN(n791) );
  NAND2_X1 U868 ( .A1(n791), .A2(G559), .ZN(n793) );
  INV_X1 U869 ( .A(n792), .ZN(n817) );
  NAND2_X1 U870 ( .A1(n793), .A2(n817), .ZN(n794) );
  XNOR2_X1 U871 ( .A(n794), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U872 ( .A1(n817), .A2(G868), .ZN(n795) );
  NOR2_X1 U873 ( .A1(G559), .A2(n795), .ZN(n797) );
  AND2_X1 U874 ( .A1(n829), .A2(n955), .ZN(n796) );
  NOR2_X1 U875 ( .A1(n797), .A2(n796), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n551), .ZN(n798) );
  XNOR2_X1 U877 ( .A(n798), .B(KEYINPUT18), .ZN(n800) );
  NAND2_X1 U878 ( .A1(n897), .A2(G99), .ZN(n799) );
  NAND2_X1 U879 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U880 ( .A1(n901), .A2(G111), .ZN(n802) );
  NAND2_X1 U881 ( .A1(G135), .A2(n898), .ZN(n801) );
  NAND2_X1 U882 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U883 ( .A1(n804), .A2(n803), .ZN(n993) );
  XNOR2_X1 U884 ( .A(G2096), .B(n993), .ZN(n805) );
  INV_X1 U885 ( .A(G2100), .ZN(n862) );
  NAND2_X1 U886 ( .A1(n805), .A2(n862), .ZN(G156) );
  NAND2_X1 U887 ( .A1(G93), .A2(n806), .ZN(n809) );
  NAND2_X1 U888 ( .A1(G80), .A2(n807), .ZN(n808) );
  NAND2_X1 U889 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U890 ( .A1(n810), .A2(G67), .ZN(n811) );
  XOR2_X1 U891 ( .A(KEYINPUT84), .B(n811), .Z(n812) );
  NOR2_X1 U892 ( .A1(n813), .A2(n812), .ZN(n816) );
  NAND2_X1 U893 ( .A1(n814), .A2(G55), .ZN(n815) );
  NAND2_X1 U894 ( .A1(n816), .A2(n815), .ZN(n830) );
  NAND2_X1 U895 ( .A1(G559), .A2(n817), .ZN(n818) );
  XOR2_X1 U896 ( .A(n818), .B(n955), .Z(n827) );
  NOR2_X1 U897 ( .A1(n827), .A2(G860), .ZN(n819) );
  XNOR2_X1 U898 ( .A(n819), .B(KEYINPUT83), .ZN(n820) );
  XNOR2_X1 U899 ( .A(n830), .B(n820), .ZN(G145) );
  XNOR2_X1 U900 ( .A(KEYINPUT19), .B(G288), .ZN(n821) );
  XNOR2_X1 U901 ( .A(n821), .B(G290), .ZN(n824) );
  XOR2_X1 U902 ( .A(G303), .B(G305), .Z(n822) );
  XNOR2_X1 U903 ( .A(n822), .B(n830), .ZN(n823) );
  XNOR2_X1 U904 ( .A(n824), .B(n823), .ZN(n826) );
  XNOR2_X1 U905 ( .A(G299), .B(KEYINPUT86), .ZN(n825) );
  XNOR2_X1 U906 ( .A(n826), .B(n825), .ZN(n852) );
  XNOR2_X1 U907 ( .A(n852), .B(n827), .ZN(n828) );
  NOR2_X1 U908 ( .A1(n829), .A2(n828), .ZN(n832) );
  NOR2_X1 U909 ( .A1(G868), .A2(n830), .ZN(n831) );
  NOR2_X1 U910 ( .A1(n832), .A2(n831), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2084), .A2(G2078), .ZN(n833) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n833), .Z(n834) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n834), .ZN(n835) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n835), .ZN(n836) );
  NAND2_X1 U915 ( .A1(n836), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U916 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U917 ( .A1(G69), .A2(G120), .ZN(n837) );
  NOR2_X1 U918 ( .A1(G237), .A2(n837), .ZN(n838) );
  NAND2_X1 U919 ( .A1(G108), .A2(n838), .ZN(n850) );
  NAND2_X1 U920 ( .A1(n850), .A2(G567), .ZN(n845) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n840) );
  NAND2_X1 U922 ( .A1(G132), .A2(G82), .ZN(n839) );
  XNOR2_X1 U923 ( .A(n840), .B(n839), .ZN(n841) );
  NOR2_X1 U924 ( .A1(G218), .A2(n841), .ZN(n842) );
  NAND2_X1 U925 ( .A1(G96), .A2(n842), .ZN(n843) );
  XNOR2_X1 U926 ( .A(KEYINPUT88), .B(n843), .ZN(n851) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n851), .ZN(n844) );
  NAND2_X1 U928 ( .A1(n845), .A2(n844), .ZN(n924) );
  NAND2_X1 U929 ( .A1(G661), .A2(G483), .ZN(n846) );
  NOR2_X1 U930 ( .A1(n924), .A2(n846), .ZN(n849) );
  NAND2_X1 U931 ( .A1(n849), .A2(G36), .ZN(G176) );
  INV_X1 U932 ( .A(G301), .ZN(G171) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n925), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U935 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U937 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U939 ( .A(G132), .ZN(G219) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G82), .ZN(G220) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(n852), .B(G286), .Z(n854) );
  XOR2_X1 U947 ( .A(G301), .B(n955), .Z(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U949 ( .A(n855), .B(n962), .Z(n856) );
  NOR2_X1 U950 ( .A1(G37), .A2(n856), .ZN(G397) );
  XOR2_X1 U951 ( .A(KEYINPUT111), .B(G2090), .Z(n858) );
  XNOR2_X1 U952 ( .A(G2084), .B(G2078), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U954 ( .A(n859), .B(G2096), .Z(n861) );
  XNOR2_X1 U955 ( .A(G2072), .B(G2067), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n866) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n864) );
  XOR2_X1 U958 ( .A(G2678), .B(n862), .Z(n863) );
  XNOR2_X1 U959 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U960 ( .A(n866), .B(n865), .Z(G227) );
  XOR2_X1 U961 ( .A(G1981), .B(G1956), .Z(n868) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1961), .ZN(n867) );
  XNOR2_X1 U963 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U964 ( .A(n869), .B(G2474), .Z(n872) );
  XOR2_X1 U965 ( .A(n870), .B(G1991), .Z(n871) );
  XNOR2_X1 U966 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U967 ( .A(KEYINPUT41), .B(G1986), .Z(n874) );
  XNOR2_X1 U968 ( .A(G1971), .B(G1976), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U970 ( .A(n876), .B(n875), .ZN(G229) );
  XOR2_X1 U971 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n878) );
  NAND2_X1 U972 ( .A1(G124), .A2(n551), .ZN(n877) );
  XNOR2_X1 U973 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n879), .B(KEYINPUT112), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n897), .A2(G100), .ZN(n880) );
  NAND2_X1 U976 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U977 ( .A1(n901), .A2(G112), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G136), .A2(n898), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U980 ( .A1(n885), .A2(n884), .ZN(G162) );
  XOR2_X1 U981 ( .A(G160), .B(G162), .Z(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n896) );
  NAND2_X1 U983 ( .A1(G130), .A2(n551), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G118), .A2(n901), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G106), .A2(n897), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G142), .A2(n898), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  NOR2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U991 ( .A(n896), .B(n895), .Z(n908) );
  NAND2_X1 U992 ( .A1(G103), .A2(n897), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G139), .A2(n898), .ZN(n899) );
  NAND2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n906) );
  NAND2_X1 U995 ( .A1(G127), .A2(n551), .ZN(n903) );
  NAND2_X1 U996 ( .A1(G115), .A2(n901), .ZN(n902) );
  NAND2_X1 U997 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n986) );
  XNOR2_X1 U1000 ( .A(n993), .B(n986), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1004 ( .A(n912), .B(n911), .Z(n915) );
  XNOR2_X1 U1005 ( .A(G164), .B(n913), .ZN(n914) );
  XNOR2_X1 U1006 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1007 ( .A1(n916), .A2(G37), .ZN(n917) );
  XNOR2_X1 U1008 ( .A(n917), .B(KEYINPUT114), .ZN(G395) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n924), .ZN(n921) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G397), .A2(n919), .ZN(n920) );
  NAND2_X1 U1013 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(n922), .A2(G395), .ZN(n923) );
  XOR2_X1 U1015 ( .A(n923), .B(KEYINPUT115), .Z(G308) );
  INV_X1 U1016 ( .A(G308), .ZN(G225) );
  INV_X1 U1017 ( .A(n924), .ZN(G319) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  INV_X1 U1019 ( .A(n925), .ZN(G223) );
  XNOR2_X1 U1020 ( .A(n926), .B(G5), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(G1966), .B(G21), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(G1971), .B(G22), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(G23), .B(G1976), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1025 ( .A(G1986), .B(G24), .Z(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT58), .B(n931), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n946) );
  XOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .Z(n936) );
  XNOR2_X1 U1031 ( .A(G4), .B(n936), .ZN(n943) );
  XOR2_X1 U1032 ( .A(G19), .B(G1341), .Z(n940) );
  XNOR2_X1 U1033 ( .A(G1956), .B(G20), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(G6), .B(G1981), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT125), .B(n941), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT60), .B(n944), .Z(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n947), .Z(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT124), .B(G16), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n976) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(n950), .B(KEYINPUT123), .ZN(n974) );
  XOR2_X1 U1046 ( .A(G301), .B(G1961), .Z(n952) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G1956), .B(G299), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n970) );
  XOR2_X1 U1050 ( .A(n956), .B(n955), .Z(n958) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n968) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n961), .B(KEYINPUT57), .ZN(n966) );
  XOR2_X1 U1055 ( .A(n962), .B(G1348), .Z(n964) );
  XOR2_X1 U1056 ( .A(G166), .B(G1971), .Z(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1062 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1063 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(n977), .B(KEYINPUT126), .ZN(n978) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n978), .ZN(n1030) );
  XNOR2_X1 U1066 ( .A(G160), .B(G2084), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(n979), .B(KEYINPUT116), .ZN(n984) );
  XOR2_X1 U1068 ( .A(G2090), .B(G162), .Z(n980) );
  NOR2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1070 ( .A(KEYINPUT51), .B(n982), .Z(n983) );
  NAND2_X1 U1071 ( .A1(n984), .A2(n983), .ZN(n1000) );
  XOR2_X1 U1072 ( .A(G164), .B(G2078), .Z(n985) );
  XNOR2_X1 U1073 ( .A(KEYINPUT118), .B(n985), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G2072), .B(n986), .Z(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(n989), .B(KEYINPUT50), .ZN(n991) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n996) );
  NOR2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(KEYINPUT117), .B(n994), .ZN(n995) );
  NOR2_X1 U1080 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1081 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1082 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1083 ( .A(KEYINPUT52), .B(n1001), .ZN(n1002) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n1004) );
  NAND2_X1 U1085 ( .A1(n1002), .A2(n1004), .ZN(n1003) );
  NAND2_X1 U1086 ( .A1(n1003), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1087 ( .A(n1004), .B(KEYINPUT121), .ZN(n1024) );
  XNOR2_X1 U1088 ( .A(G2090), .B(G35), .ZN(n1019) );
  XNOR2_X1 U1089 ( .A(KEYINPUT119), .B(G2067), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1005), .B(G26), .ZN(n1013) );
  XNOR2_X1 U1091 ( .A(G2072), .B(G33), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G1991), .B(G25), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(G28), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT120), .B(G1996), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G32), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(G27), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(KEYINPUT53), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1103 ( .A(G2084), .B(G34), .Z(n1020) );
  XNOR2_X1 U1104 ( .A(KEYINPUT54), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NOR2_X1 U1107 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(KEYINPUT122), .B(n1026), .Z(n1027) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1110 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1031), .Z(n1032) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1032), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

