

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U322 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n416) );
  XOR2_X1 U323 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n290) );
  XOR2_X1 U324 ( .A(n352), .B(n351), .Z(n291) );
  XOR2_X1 U325 ( .A(n334), .B(n333), .Z(n292) );
  XOR2_X1 U326 ( .A(n347), .B(n390), .Z(n293) );
  XNOR2_X1 U327 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U328 ( .A(n421), .B(n420), .ZN(n424) );
  XNOR2_X1 U329 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n470) );
  NOR2_X1 U330 ( .A1(n516), .A2(n548), .ZN(n478) );
  XNOR2_X1 U331 ( .A(n471), .B(n470), .ZN(n476) );
  NOR2_X1 U332 ( .A1(n491), .A2(n481), .ZN(n483) );
  XNOR2_X1 U333 ( .A(n353), .B(n291), .ZN(n354) );
  XNOR2_X1 U334 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U335 ( .A(n381), .B(KEYINPUT99), .ZN(n382) );
  XNOR2_X1 U336 ( .A(n355), .B(n354), .ZN(n360) );
  XNOR2_X1 U337 ( .A(n439), .B(n438), .ZN(n465) );
  XNOR2_X1 U338 ( .A(n383), .B(n382), .ZN(n567) );
  XNOR2_X1 U339 ( .A(n417), .B(n416), .ZN(n535) );
  XNOR2_X1 U340 ( .A(n486), .B(n485), .ZN(n583) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n462) );
  XNOR2_X1 U342 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U343 ( .A(n462), .B(KEYINPUT40), .ZN(n463) );
  XNOR2_X1 U344 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n464), .B(n463), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n295), .B(n294), .ZN(n305) );
  XOR2_X1 U349 ( .A(G190GAT), .B(G99GAT), .Z(n297) );
  XOR2_X1 U350 ( .A(G71GAT), .B(G120GAT), .Z(n427) );
  XOR2_X1 U351 ( .A(G113GAT), .B(KEYINPUT0), .Z(n387) );
  XNOR2_X1 U352 ( .A(n427), .B(n387), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .Z(n323) );
  XOR2_X1 U355 ( .A(n298), .B(n323), .Z(n303) );
  XOR2_X1 U356 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n300) );
  NAND2_X1 U357 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U359 ( .A(KEYINPUT87), .B(n301), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U362 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(n308), .ZN(n369) );
  XNOR2_X1 U366 ( .A(n309), .B(n369), .ZN(n553) );
  XOR2_X1 U367 ( .A(KEYINPUT15), .B(G64GAT), .Z(n311) );
  XNOR2_X1 U368 ( .A(G183GAT), .B(G211GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U370 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n313) );
  XNOR2_X1 U371 ( .A(KEYINPUT14), .B(KEYINPUT81), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U373 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U374 ( .A(G8GAT), .B(KEYINPUT80), .Z(n368) );
  XOR2_X1 U375 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n317) );
  NAND2_X1 U376 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n368), .B(n318), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n329) );
  XOR2_X1 U380 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n322) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G78GAT), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G155GAT), .Z(n350) );
  XOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT13), .Z(n434) );
  XOR2_X1 U385 ( .A(n350), .B(n434), .Z(n325) );
  XOR2_X1 U386 ( .A(KEYINPUT68), .B(G1GAT), .Z(n451) );
  XNOR2_X1 U387 ( .A(n451), .B(n323), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U389 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n593) );
  INV_X1 U391 ( .A(n593), .ZN(n497) );
  XOR2_X1 U392 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n331) );
  XNOR2_X1 U393 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n334) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n290), .B(n332), .ZN(n333) );
  XOR2_X1 U397 ( .A(G134GAT), .B(KEYINPUT78), .Z(n386) );
  XOR2_X1 U398 ( .A(G36GAT), .B(G190GAT), .Z(n373) );
  XNOR2_X1 U399 ( .A(n386), .B(n373), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n292), .B(n335), .ZN(n339) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n347) );
  XOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .Z(n435) );
  XOR2_X1 U403 ( .A(n347), .B(n435), .Z(n337) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U406 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U407 ( .A(KEYINPUT67), .B(KEYINPUT8), .Z(n341) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G29GAT), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U410 ( .A(KEYINPUT7), .B(n342), .Z(n459) );
  XNOR2_X1 U411 ( .A(n459), .B(G92GAT), .ZN(n343) );
  XNOR2_X2 U412 ( .A(n344), .B(n343), .ZN(n575) );
  XOR2_X1 U413 ( .A(n575), .B(KEYINPUT104), .Z(n345) );
  XNOR2_X1 U414 ( .A(KEYINPUT36), .B(n345), .ZN(n493) );
  XNOR2_X1 U415 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n346), .B(KEYINPUT2), .ZN(n390) );
  NAND2_X1 U417 ( .A1(G228GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n293), .B(n348), .ZN(n349) );
  XOR2_X1 U419 ( .A(n349), .B(KEYINPUT22), .Z(n355) );
  XNOR2_X1 U420 ( .A(G204GAT), .B(n350), .ZN(n353) );
  XOR2_X1 U421 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n352) );
  XNOR2_X1 U422 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n351) );
  XOR2_X1 U423 ( .A(G211GAT), .B(KEYINPUT21), .Z(n357) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(G218GAT), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n367) );
  XNOR2_X1 U426 ( .A(G148GAT), .B(G106GAT), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n358), .B(G78GAT), .ZN(n430) );
  XNOR2_X1 U428 ( .A(n367), .B(n430), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n481) );
  INV_X1 U430 ( .A(G204GAT), .ZN(n361) );
  NAND2_X1 U431 ( .A1(n361), .A2(G64GAT), .ZN(n364) );
  INV_X1 U432 ( .A(G64GAT), .ZN(n362) );
  NAND2_X1 U433 ( .A1(n362), .A2(G204GAT), .ZN(n363) );
  NAND2_X1 U434 ( .A1(n364), .A2(n363), .ZN(n366) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G92GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n421) );
  XNOR2_X1 U437 ( .A(n367), .B(n421), .ZN(n377) );
  XOR2_X1 U438 ( .A(n368), .B(KEYINPUT97), .Z(n371) );
  XOR2_X1 U439 ( .A(n369), .B(KEYINPUT96), .Z(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U441 ( .A(n373), .B(n372), .Z(n375) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n516) );
  NOR2_X1 U445 ( .A1(n516), .A2(n553), .ZN(n378) );
  NOR2_X1 U446 ( .A1(n481), .A2(n378), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n379), .B(KEYINPUT101), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n380), .B(KEYINPUT25), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n516), .B(KEYINPUT27), .ZN(n410) );
  NAND2_X1 U450 ( .A1(n481), .A2(n553), .ZN(n383) );
  XOR2_X1 U451 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n381) );
  NOR2_X1 U452 ( .A1(n410), .A2(n567), .ZN(n384) );
  NOR2_X1 U453 ( .A1(n385), .A2(n384), .ZN(n409) );
  XOR2_X1 U454 ( .A(G85GAT), .B(G162GAT), .Z(n389) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n394) );
  XOR2_X1 U457 ( .A(n390), .B(KEYINPUT1), .Z(n392) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U460 ( .A(n394), .B(n393), .Z(n396) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(G127GAT), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U463 ( .A(G57GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(G120GAT), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U466 ( .A(n400), .B(n399), .Z(n408) );
  XOR2_X1 U467 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n402) );
  XNOR2_X1 U468 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U470 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n404) );
  XNOR2_X1 U471 ( .A(G148GAT), .B(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n512) );
  INV_X1 U475 ( .A(n512), .ZN(n536) );
  NOR2_X1 U476 ( .A1(n409), .A2(n536), .ZN(n414) );
  NOR2_X1 U477 ( .A1(n512), .A2(n410), .ZN(n411) );
  XOR2_X1 U478 ( .A(KEYINPUT98), .B(n411), .Z(n549) );
  XOR2_X1 U479 ( .A(n481), .B(KEYINPUT28), .Z(n520) );
  NAND2_X1 U480 ( .A1(n553), .A2(n520), .ZN(n412) );
  NOR2_X1 U481 ( .A1(n549), .A2(n412), .ZN(n413) );
  NOR2_X1 U482 ( .A1(n414), .A2(n413), .ZN(n499) );
  NOR2_X1 U483 ( .A1(n493), .A2(n499), .ZN(n415) );
  NAND2_X1 U484 ( .A1(n497), .A2(n415), .ZN(n417) );
  NAND2_X1 U485 ( .A1(G230GAT), .A2(G233GAT), .ZN(n419) );
  INV_X1 U486 ( .A(KEYINPUT74), .ZN(n418) );
  INV_X1 U487 ( .A(n424), .ZN(n423) );
  INV_X1 U488 ( .A(KEYINPUT75), .ZN(n422) );
  NAND2_X1 U489 ( .A1(n423), .A2(n422), .ZN(n426) );
  NAND2_X1 U490 ( .A1(n424), .A2(KEYINPUT75), .ZN(n425) );
  NAND2_X1 U491 ( .A1(n426), .A2(n425), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n427), .B(KEYINPUT33), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n439) );
  XOR2_X1 U495 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n433) );
  XNOR2_X1 U496 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n432) );
  XOR2_X1 U497 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U499 ( .A(KEYINPUT30), .B(G22GAT), .Z(n441) );
  XNOR2_X1 U500 ( .A(G8GAT), .B(G15GAT), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U502 ( .A(G113GAT), .B(G141GAT), .Z(n443) );
  XNOR2_X1 U503 ( .A(KEYINPUT71), .B(KEYINPUT65), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n457) );
  XOR2_X1 U506 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n447) );
  XNOR2_X1 U507 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n455) );
  XOR2_X1 U509 ( .A(G197GAT), .B(G36GAT), .Z(n449) );
  XNOR2_X1 U510 ( .A(G169GAT), .B(G50GAT), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U512 ( .A(n451), .B(n450), .Z(n453) );
  NAND2_X1 U513 ( .A1(G229GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(n585) );
  NAND2_X1 U518 ( .A1(n465), .A2(n585), .ZN(n502) );
  NOR2_X1 U519 ( .A1(n535), .A2(n502), .ZN(n460) );
  XOR2_X1 U520 ( .A(n460), .B(KEYINPUT38), .Z(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT106), .B(n461), .ZN(n519) );
  NOR2_X1 U522 ( .A1(n553), .A2(n519), .ZN(n464) );
  INV_X1 U523 ( .A(KEYINPUT125), .ZN(n486) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT41), .ZN(n579) );
  NAND2_X1 U525 ( .A1(n579), .A2(n585), .ZN(n467) );
  XOR2_X1 U526 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n593), .A2(n575), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n497), .A2(n493), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT45), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n465), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n585), .A2(n474), .ZN(n475) );
  NOR2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT48), .ZN(n548) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT54), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n512), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT64), .ZN(n491) );
  XNOR2_X1 U539 ( .A(KEYINPUT124), .B(KEYINPUT55), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n484), .A2(n553), .ZN(n485) );
  NAND2_X1 U542 ( .A1(n583), .A2(n575), .ZN(n490) );
  XOR2_X1 U543 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n488) );
  INV_X1 U544 ( .A(G190GAT), .ZN(n487) );
  INV_X1 U545 ( .A(G218GAT), .ZN(n496) );
  NOR2_X1 U546 ( .A1(n491), .A2(n567), .ZN(n492) );
  XOR2_X1 U547 ( .A(KEYINPUT127), .B(n492), .Z(n592) );
  INV_X1 U548 ( .A(n592), .ZN(n589) );
  NOR2_X1 U549 ( .A1(n493), .A2(n589), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT62), .B(n494), .ZN(n495) );
  XNOR2_X1 U551 ( .A(n496), .B(n495), .ZN(G1355GAT) );
  NOR2_X1 U552 ( .A1(n575), .A2(n497), .ZN(n498) );
  XNOR2_X1 U553 ( .A(n498), .B(KEYINPUT16), .ZN(n501) );
  INV_X1 U554 ( .A(n499), .ZN(n500) );
  NAND2_X1 U555 ( .A1(n501), .A2(n500), .ZN(n524) );
  NOR2_X1 U556 ( .A1(n502), .A2(n524), .ZN(n510) );
  NAND2_X1 U557 ( .A1(n536), .A2(n510), .ZN(n505) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n503) );
  XNOR2_X1 U559 ( .A(n503), .B(KEYINPUT102), .ZN(n504) );
  XNOR2_X1 U560 ( .A(n505), .B(n504), .ZN(G1324GAT) );
  INV_X1 U561 ( .A(n516), .ZN(n539) );
  NAND2_X1 U562 ( .A1(n539), .A2(n510), .ZN(n506) );
  XNOR2_X1 U563 ( .A(n506), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n508) );
  INV_X1 U565 ( .A(n553), .ZN(n542) );
  NAND2_X1 U566 ( .A1(n510), .A2(n542), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U568 ( .A(G15GAT), .B(n509), .Z(G1326GAT) );
  INV_X1 U569 ( .A(n520), .ZN(n551) );
  NAND2_X1 U570 ( .A1(n551), .A2(n510), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n511), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U572 ( .A1(n512), .A2(n519), .ZN(n514) );
  XNOR2_X1 U573 ( .A(KEYINPUT39), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U575 ( .A(G29GAT), .B(n515), .Z(G1328GAT) );
  NOR2_X1 U576 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(n517), .Z(n518) );
  XNOR2_X1 U578 ( .A(G36GAT), .B(n518), .ZN(G1329GAT) );
  NOR2_X1 U579 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U580 ( .A(G50GAT), .B(n521), .Z(G1331GAT) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n526) );
  INV_X1 U582 ( .A(n585), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n579), .A2(n522), .ZN(n523) );
  XOR2_X1 U584 ( .A(KEYINPUT109), .B(n523), .Z(n534) );
  NOR2_X1 U585 ( .A1(n534), .A2(n524), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n530), .A2(n536), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n526), .B(n525), .ZN(G1332GAT) );
  NAND2_X1 U588 ( .A1(n539), .A2(n530), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT110), .ZN(n528) );
  XNOR2_X1 U590 ( .A(G64GAT), .B(n528), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n530), .A2(n542), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n532) );
  NAND2_X1 U594 ( .A1(n530), .A2(n551), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U596 ( .A(G78GAT), .B(n533), .Z(G1335GAT) );
  NOR2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n536), .A2(n545), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n537), .B(KEYINPUT112), .ZN(n538) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n538), .ZN(G1336GAT) );
  XOR2_X1 U601 ( .A(G92GAT), .B(KEYINPUT113), .Z(n541) );
  NAND2_X1 U602 ( .A1(n545), .A2(n539), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(G1337GAT) );
  NAND2_X1 U604 ( .A1(n545), .A2(n542), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT114), .ZN(n544) );
  XNOR2_X1 U606 ( .A(G99GAT), .B(n544), .ZN(G1338GAT) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n545), .A2(n551), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(G1339GAT) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(KEYINPUT118), .ZN(n555) );
  NOR2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT117), .B(n550), .ZN(n566) );
  OR2_X1 U613 ( .A1(n566), .A2(n551), .ZN(n552) );
  NOR2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n562) );
  NAND2_X1 U615 ( .A1(n562), .A2(n585), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n555), .B(n554), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n557) );
  NAND2_X1 U618 ( .A1(n562), .A2(n579), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U620 ( .A(G120GAT), .B(n558), .Z(G1341GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n560) );
  NAND2_X1 U622 ( .A1(n562), .A2(n593), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(G127GAT), .B(n561), .Z(G1342GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT51), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U626 ( .A1(n562), .A2(n575), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U628 ( .A(G134GAT), .B(n565), .Z(G1343GAT) );
  NOR2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n576), .A2(n585), .ZN(n568) );
  XNOR2_X1 U631 ( .A(G141GAT), .B(n568), .ZN(G1344GAT) );
  XNOR2_X1 U632 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n570) );
  NAND2_X1 U634 ( .A1(n576), .A2(n579), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(G1345GAT) );
  XOR2_X1 U637 ( .A(G155GAT), .B(KEYINPUT123), .Z(n574) );
  NAND2_X1 U638 ( .A1(n576), .A2(n593), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1346GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U642 ( .A1(n585), .A2(n583), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U644 ( .A1(n583), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U648 ( .A1(n593), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n587) );
  NAND2_X1 U651 ( .A1(n592), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .Z(n591) );
  OR2_X1 U655 ( .A1(n589), .A2(n465), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
endmodule

