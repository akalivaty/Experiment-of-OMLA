//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(KEYINPUT64), .A3(G143), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(new_n188), .B2(G146), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n196), .B(new_n197), .C1(new_n199), .C2(new_n189), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT65), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT64), .B1(new_n190), .B2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n190), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n196), .A4(new_n197), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n194), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n212), .A3(KEYINPUT11), .A4(G134), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n209), .B2(G137), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n212), .A2(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n218), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n208), .B1(new_n217), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n217), .A2(new_n208), .A3(new_n224), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n207), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT2), .B(G113), .Z(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n203), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G128), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n189), .A2(new_n191), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n236), .B2(new_n237), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n204), .A3(new_n197), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n217), .A2(new_n208), .A3(new_n224), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n222), .A2(new_n210), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n250), .A3(G131), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n227), .A2(new_n233), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n257), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n233), .B1(new_n227), .B2(new_n253), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n227), .A2(KEYINPUT70), .A3(new_n233), .A4(new_n253), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n256), .B(new_n264), .C1(new_n269), .C2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n187), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n217), .A2(new_n224), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n246), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n241), .A2(new_n244), .B1(new_n249), .B2(new_n251), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n277), .A2(new_n207), .B1(new_n246), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT70), .B1(new_n279), .B2(new_n233), .ZN(new_n280));
  INV_X1    g094(.A(new_n268), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n227), .A2(KEYINPUT30), .A3(new_n253), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT30), .B1(new_n227), .B2(new_n253), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n283), .A2(new_n284), .A3(new_n233), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n263), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n270), .A2(new_n286), .A3(new_n271), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT73), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT74), .B(new_n187), .C1(new_n270), .C2(new_n271), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n270), .A2(new_n286), .A3(new_n290), .A4(new_n271), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n274), .A2(new_n288), .A3(new_n289), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G472), .ZN(new_n293));
  INV_X1    g107(.A(G472), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n279), .A2(KEYINPUT30), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n227), .A2(new_n253), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n298), .A3(new_n232), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n267), .A2(new_n268), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(new_n264), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT31), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n299), .A2(new_n300), .A3(new_n303), .A4(new_n264), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n265), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n280), .B2(new_n281), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n264), .B1(new_n308), .B2(new_n256), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n294), .B(new_n187), .C1(new_n305), .C2(new_n309), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n310), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT32), .B1(new_n310), .B2(KEYINPUT72), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n293), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G122), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G116), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(G116), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G107), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT89), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT14), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n315), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n321), .A2(KEYINPUT90), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n320), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n321), .B2(KEYINPUT90), .ZN(new_n324));
  OAI21_X1  g138(.A(G107), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n188), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n242), .A2(G143), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT88), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT88), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G134), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n209), .B1(new_n332), .B2(new_n328), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n319), .A2(new_n325), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n327), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n326), .A2(new_n336), .ZN(new_n339));
  OAI21_X1  g153(.A(G134), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n316), .A2(new_n317), .ZN(new_n341));
  INV_X1    g155(.A(G107), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n333), .B(new_n340), .C1(new_n343), .C2(new_n318), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT9), .B(G234), .Z(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G217), .A3(new_n259), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n347), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n187), .ZN(new_n352));
  INV_X1    g166(.A(G478), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(KEYINPUT15), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n352), .B(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G113), .B(G122), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G125), .B(G140), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT19), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n190), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT16), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(G125), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(G146), .B(new_n368), .C1(new_n372), .C2(new_n366), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n258), .A2(new_n259), .A3(G214), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(new_n188), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(G143), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n208), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n365), .A2(KEYINPUT86), .A3(new_n373), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT18), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n380), .B1(new_n385), .B2(new_n208), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n363), .B(new_n190), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n386), .B(new_n387), .C1(new_n385), .C2(new_n379), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n362), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n368), .B1(new_n372), .B2(new_n366), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n190), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n373), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n378), .A2(KEYINPUT17), .A3(G131), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n393), .B(new_n394), .C1(new_n382), .C2(KEYINPUT17), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n362), .A3(new_n388), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n359), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(new_n357), .C1(new_n389), .C2(new_n397), .ZN(new_n402));
  INV_X1    g216(.A(G234), .ZN(new_n403));
  OAI211_X1 g217(.A(G952), .B(new_n259), .C1(new_n403), .C2(new_n258), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(KEYINPUT91), .Z(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(G902), .B(G953), .C1(new_n403), .C2(new_n258), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT92), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT21), .B(G898), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n362), .B1(new_n395), .B2(new_n388), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n187), .B1(new_n397), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n414), .B2(G475), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n356), .A2(new_n401), .A3(new_n402), .A4(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n241), .A2(new_n370), .A3(new_n244), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n207), .B2(new_n370), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n259), .A2(G224), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT79), .B1(new_n342), .B2(G104), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n361), .A3(G107), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT3), .B1(new_n361), .B2(G107), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n342), .A3(G104), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G101), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n425), .ZN(new_n432));
  INV_X1    g246(.A(G101), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n427), .A4(new_n429), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(G101), .C1(new_n426), .C2(new_n430), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n232), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n342), .A2(G104), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n361), .A2(G107), .ZN(new_n440));
  OAI21_X1  g254(.A(G101), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G116), .ZN(new_n444));
  INV_X1    g258(.A(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n443), .A3(G116), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G113), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n231), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(G110), .B(G122), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n438), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT7), .B1(new_n420), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n457), .B2(new_n420), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n418), .B(new_n459), .C1(new_n207), .C2(new_n370), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n422), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n454), .B(KEYINPUT8), .Z(new_n462));
  AND2_X1   g276(.A1(new_n434), .A2(new_n441), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(new_n447), .B2(new_n448), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n229), .A2(new_n465), .A3(KEYINPUT5), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n464), .A2(G113), .A3(new_n466), .A4(new_n450), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n231), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n442), .A2(new_n452), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n468), .B2(KEYINPUT84), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n461), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n438), .A2(new_n453), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n454), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n478), .A3(new_n454), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n420), .B(KEYINPUT82), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n419), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n473), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n474), .B1(new_n473), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n417), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n416), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G221), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n346), .B2(new_n187), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n442), .A2(new_n241), .A3(new_n244), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n243), .A2(new_n204), .A3(new_n197), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n204), .A2(new_n197), .B1(G128), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n434), .B(new_n441), .C1(new_n491), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n277), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT12), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n207), .A2(new_n435), .A3(new_n437), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT10), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n226), .A2(new_n225), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n241), .B2(new_n244), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n463), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n495), .A2(new_n505), .A3(new_n277), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G140), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n259), .A2(G227), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n498), .A2(new_n500), .A3(new_n503), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT80), .B1(new_n226), .B2(new_n225), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n494), .A2(new_n499), .B1(new_n502), .B2(new_n463), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n514), .A3(new_n498), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n518), .A3(new_n510), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n512), .A2(G469), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(G469), .A2(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND4_X1   g336(.A1(new_n514), .A2(new_n498), .A3(new_n500), .A4(new_n503), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n514), .B1(new_n517), .B2(new_n498), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n511), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n497), .A2(new_n510), .A3(new_n504), .A4(new_n506), .ZN(new_n526));
  AOI211_X1 g340(.A(G469), .B(G902), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT81), .B(new_n489), .C1(new_n522), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G469), .ZN(new_n530));
  INV_X1    g344(.A(new_n526), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n510), .B1(new_n516), .B2(new_n518), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n530), .B(new_n187), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n521), .A3(new_n520), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT81), .B1(new_n534), .B2(new_n489), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n486), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT93), .ZN(new_n537));
  OAI21_X1  g351(.A(G217), .B1(new_n403), .B2(G902), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n487), .A2(new_n403), .A3(G953), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n242), .A2(G119), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n242), .A2(G119), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT23), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n242), .A3(G119), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT75), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G110), .B1(new_n548), .B2(KEYINPUT75), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT76), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n547), .ZN(new_n553));
  INV_X1    g367(.A(new_n543), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT75), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n549), .A4(G110), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n554), .A3(new_n544), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n552), .A2(new_n559), .A3(new_n561), .A4(new_n392), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n555), .A2(G110), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n554), .B2(new_n544), .ZN(new_n564));
  OAI221_X1 g378(.A(new_n373), .B1(G146), .B2(new_n372), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n562), .A2(KEYINPUT77), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT77), .B1(new_n562), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n542), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n565), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT77), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n541), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n187), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT78), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT25), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n538), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n568), .A2(new_n187), .A3(new_n571), .A4(new_n574), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n538), .A2(new_n187), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n568), .A2(new_n571), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n486), .B(new_n584), .C1(new_n529), .C2(new_n535), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n313), .A2(new_n537), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  OAI21_X1  g401(.A(new_n187), .B1(new_n305), .B2(new_n309), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n310), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n582), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n529), .A2(new_n535), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n473), .A2(new_n482), .A3(new_n474), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT94), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n417), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n483), .A2(new_n484), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(new_n594), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n412), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n414), .A2(G475), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n401), .A2(new_n402), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n351), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n348), .A2(KEYINPUT33), .A3(new_n350), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(G478), .A3(new_n187), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n352), .A2(new_n353), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n598), .A2(new_n599), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  XNOR2_X1  g426(.A(new_n600), .B(KEYINPUT95), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n352), .B(new_n354), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n401), .A2(new_n402), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n598), .A2(new_n599), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NOR2_X1   g433(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n569), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n580), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n576), .B2(new_n577), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n590), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n537), .A2(new_n625), .A3(new_n585), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G110), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G12));
  NAND2_X1  g443(.A1(new_n578), .A2(new_n622), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n597), .B(new_n630), .C1(new_n529), .C2(new_n535), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n406), .B1(new_n632), .B2(new_n409), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT97), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n616), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n313), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  XNOR2_X1  g452(.A(new_n596), .B(KEYINPUT38), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n624), .A2(new_n614), .A3(new_n417), .A4(new_n601), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n634), .B(KEYINPUT39), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n592), .A2(new_n641), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n639), .B(new_n640), .C1(new_n642), .C2(KEYINPUT40), .ZN(new_n643));
  INV_X1    g457(.A(new_n301), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n269), .A2(new_n264), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n187), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G472), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n311), .B2(new_n312), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT98), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n643), .A2(new_n652), .A3(new_n648), .A4(new_n649), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n188), .ZN(G45));
  AND3_X1   g469(.A1(new_n601), .A2(new_n607), .A3(new_n634), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n313), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT99), .B(G146), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G48));
  INV_X1    g475(.A(new_n597), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n525), .A2(new_n526), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n187), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G469), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n533), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n489), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n313), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n582), .A2(new_n412), .A3(new_n608), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND4_X1  g488(.A1(new_n613), .A2(new_n615), .A3(new_n614), .A4(new_n599), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n582), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT100), .B(G116), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G18));
  NOR2_X1   g493(.A1(new_n624), .A2(new_n416), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n313), .A2(new_n669), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  NAND2_X1  g496(.A1(new_n601), .A2(new_n614), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n601), .A2(KEYINPUT101), .A3(new_n614), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n597), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n668), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n591), .A2(new_n599), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  AND4_X1   g505(.A1(new_n310), .A2(new_n589), .A3(new_n630), .A4(new_n656), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n669), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(new_n484), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(new_n417), .A3(new_n593), .A4(new_n634), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(new_n608), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n521), .B(KEYINPUT102), .Z(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n519), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n519), .A2(new_n699), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n512), .A3(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n533), .B(new_n698), .C1(new_n702), .C2(new_n530), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n489), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n697), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT32), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n310), .B(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n293), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n706), .B(new_n583), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n310), .B(KEYINPUT32), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n582), .B1(new_n713), .B2(new_n293), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT105), .A3(new_n706), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n596), .A2(new_n417), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n704), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n313), .A2(new_n583), .A3(new_n656), .A4(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(KEYINPUT104), .A3(new_n705), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT104), .B1(new_n719), .B2(new_n705), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  INV_X1    g537(.A(new_n635), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n313), .A2(new_n583), .A3(new_n724), .A4(new_n718), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  INV_X1    g540(.A(new_n607), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n601), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT43), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n727), .B2(new_n601), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n624), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n590), .ZN(new_n733));
  INV_X1    g547(.A(new_n717), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT44), .B1(new_n732), .B2(new_n590), .ZN(new_n737));
  OR3_X1    g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n512), .A4(new_n701), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n740), .A2(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(KEYINPUT106), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT45), .B1(new_n512), .B2(new_n519), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n530), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n698), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n533), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n745), .B2(new_n698), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n489), .B(new_n641), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n738), .A2(new_n739), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  OAI21_X1  g566(.A(new_n489), .B1(new_n747), .B2(new_n748), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n313), .A2(new_n583), .A3(new_n697), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n405), .B1(new_n729), .B2(new_n731), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n591), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n717), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT111), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n755), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n667), .A2(new_n488), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n765), .B2(KEYINPUT112), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n760), .B(new_n764), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n648), .A2(new_n582), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n770), .A2(new_n405), .A3(new_n668), .A4(new_n717), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n615), .A3(new_n600), .A4(new_n727), .ZN(new_n772));
  INV_X1    g586(.A(new_n417), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n689), .A2(new_n773), .A3(new_n639), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n762), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT50), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(KEYINPUT50), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n761), .A2(new_n689), .A3(new_n734), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n776), .A2(new_n777), .B1(new_n625), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n769), .A2(new_n772), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n765), .A2(new_n767), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n764), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT113), .B1(new_n772), .B2(new_n779), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT51), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n778), .A2(new_n714), .ZN(new_n787));
  NOR2_X1   g601(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT114), .Z(new_n789));
  OR2_X1    g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n669), .ZN(new_n794));
  OAI211_X1 g608(.A(G952), .B(new_n259), .C1(new_n762), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n771), .B2(new_n609), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n786), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n608), .B1(new_n356), .B2(new_n601), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n599), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n485), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n591), .A3(new_n592), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n586), .A2(new_n626), .A3(new_n690), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n624), .A2(new_n696), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n613), .A2(new_n615), .A3(new_n356), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n803), .B(new_n804), .C1(new_n535), .C2(new_n529), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n806), .A2(new_n313), .B1(new_n692), .B2(new_n718), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n725), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n313), .B(new_n669), .C1(new_n671), .C2(new_n676), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n681), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n802), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n722), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT109), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n624), .A2(new_n703), .A3(new_n489), .A4(new_n634), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n687), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n648), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n637), .A2(new_n659), .A3(new_n816), .A4(new_n693), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n636), .A2(new_n313), .B1(new_n692), .B2(new_n669), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n659), .A4(new_n816), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n818), .A2(new_n821), .B1(new_n822), .B2(new_n817), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n817), .A2(new_n822), .A3(new_n820), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n722), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n813), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n818), .A2(new_n821), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n722), .A3(new_n811), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n811), .A2(new_n722), .A3(KEYINPUT53), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n825), .A2(new_n834), .B1(new_n831), .B2(new_n826), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n797), .A2(new_n838), .B1(G952), .B2(G953), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n728), .A2(new_n489), .A3(new_n417), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n666), .B2(KEYINPUT49), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n666), .A2(KEYINPUT49), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT108), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n841), .A2(new_n844), .A3(new_n639), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n770), .B2(new_n846), .ZN(G75));
  AND2_X1   g661(.A1(new_n477), .A2(new_n479), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT116), .Z(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n851));
  XNOR2_X1  g665(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n481), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n834), .A2(new_n825), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n818), .A2(new_n821), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n826), .B1(new_n812), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n187), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n851), .B(new_n853), .C1(new_n857), .C2(G210), .ZN(new_n858));
  INV_X1    g672(.A(new_n853), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n812), .A2(new_n823), .A3(new_n826), .A4(new_n824), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n719), .A2(new_n705), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT104), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n719), .A2(KEYINPUT104), .A3(new_n705), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n863), .A2(new_n864), .B1(new_n712), .B2(new_n715), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n586), .A2(new_n626), .A3(new_n690), .A4(new_n801), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n807), .A2(new_n725), .ZN(new_n867));
  INV_X1    g681(.A(new_n810), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT53), .B1(new_n870), .B2(new_n830), .ZN(new_n871));
  OAI211_X1 g685(.A(G210), .B(G902), .C1(new_n860), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n851), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n859), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n849), .B1(new_n858), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(G210), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n876), .B(new_n187), .C1(new_n854), .C2(new_n856), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n853), .B1(new_n877), .B2(new_n851), .ZN(new_n878));
  INV_X1    g692(.A(new_n849), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n873), .A3(new_n859), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n259), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n875), .A2(new_n881), .A3(new_n883), .ZN(G51));
  NAND2_X1  g698(.A1(new_n854), .A2(new_n856), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n837), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n698), .B(KEYINPUT57), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n663), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n857), .A2(new_n741), .A3(new_n742), .A4(new_n744), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(G54));
  NAND3_X1  g705(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n398), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n398), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n882), .ZN(G60));
  AND2_X1   g709(.A1(new_n603), .A2(new_n604), .ZN(new_n896));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n886), .B2(new_n837), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n883), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n838), .B2(new_n898), .ZN(new_n903));
  AOI211_X1 g717(.A(KEYINPUT119), .B(new_n899), .C1(new_n886), .C2(new_n837), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G63));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n568), .A2(new_n571), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n908));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n835), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n883), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n885), .A2(new_n621), .A3(new_n910), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n912), .B2(new_n883), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n906), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n912), .A2(new_n915), .A3(KEYINPUT61), .A4(new_n883), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n911), .B1(new_n854), .B2(new_n856), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n906), .B1(new_n922), .B2(new_n621), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(KEYINPUT122), .A3(new_n883), .A4(new_n912), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n918), .A2(new_n925), .ZN(G66));
  INV_X1    g740(.A(G224), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n411), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n802), .A2(new_n810), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n849), .B1(G898), .B2(new_n259), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(G69));
  AOI21_X1  g746(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n259), .A2(G900), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n819), .A2(new_n659), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n725), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n714), .A2(new_n688), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n750), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n722), .A3(new_n751), .A4(new_n758), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n940), .B2(new_n259), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n283), .A2(new_n284), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(new_n364), .Z(new_n943));
  OR2_X1    g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n313), .A2(new_n583), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n592), .A2(new_n641), .A3(new_n734), .A4(new_n798), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n751), .B(new_n758), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n651), .A2(new_n653), .A3(new_n936), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n651), .A2(KEYINPUT62), .A3(new_n653), .A4(new_n936), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n943), .B1(new_n954), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n944), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n946), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n944), .B(new_n955), .C1(new_n945), .C2(new_n933), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(G72));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  INV_X1    g775(.A(new_n929), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n940), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n961), .C1(new_n940), .C2(new_n962), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n282), .A2(new_n285), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n263), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n964), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(new_n883), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n970), .B2(new_n883), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n967), .A2(new_n263), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n954), .A2(new_n929), .ZN(new_n975));
  INV_X1    g789(.A(new_n961), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n286), .ZN(new_n978));
  OR3_X1    g792(.A1(new_n978), .A2(KEYINPUT127), .A3(new_n644), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n978), .B2(KEYINPUT127), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n829), .A2(new_n832), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n972), .A2(new_n973), .A3(new_n982), .ZN(G57));
endmodule


