

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730;

  NOR2_X1 U376 ( .A1(n372), .A2(n569), .ZN(n542) );
  BUF_X1 U377 ( .A(n640), .Z(n354) );
  XOR2_X1 U378 ( .A(G116), .B(G119), .Z(n353) );
  XNOR2_X1 U379 ( .A(n508), .B(KEYINPUT1), .ZN(n640) );
  NAND2_X2 U380 ( .A1(n368), .A2(n367), .ZN(n694) );
  AND2_X1 U381 ( .A1(n589), .A2(KEYINPUT2), .ZN(n637) );
  NOR2_X1 U382 ( .A1(n635), .A2(n590), .ZN(n366) );
  XNOR2_X1 U383 ( .A(n359), .B(n357), .ZN(n567) );
  NAND2_X1 U384 ( .A1(n360), .A2(n552), .ZN(n359) );
  XNOR2_X1 U385 ( .A(n550), .B(n549), .ZN(n553) );
  XNOR2_X1 U386 ( .A(n392), .B(G128), .ZN(n473) );
  INV_X1 U387 ( .A(G143), .ZN(n392) );
  XNOR2_X1 U388 ( .A(n473), .B(n393), .ZN(n415) );
  NAND2_X1 U389 ( .A1(n370), .A2(n656), .ZN(n511) );
  NOR2_X1 U390 ( .A1(n500), .A2(n493), .ZN(n494) );
  XNOR2_X1 U391 ( .A(n568), .B(KEYINPUT44), .ZN(n585) );
  AND2_X1 U392 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n404) );
  XNOR2_X1 U394 ( .A(G104), .B(G113), .ZN(n469) );
  XNOR2_X1 U395 ( .A(n415), .B(n414), .ZN(n715) );
  XNOR2_X1 U396 ( .A(n364), .B(n355), .ZN(n521) );
  NAND2_X1 U397 ( .A1(n686), .A2(n420), .ZN(n364) );
  OR2_X1 U398 ( .A1(n522), .A2(n521), .ZN(n659) );
  XNOR2_X1 U399 ( .A(KEYINPUT98), .B(KEYINPUT96), .ZN(n394) );
  INV_X1 U400 ( .A(KEYINPUT11), .ZN(n386) );
  XNOR2_X1 U401 ( .A(n414), .B(n376), .ZN(n380) );
  INV_X1 U402 ( .A(G953), .ZN(n455) );
  XNOR2_X1 U403 ( .A(n486), .B(KEYINPUT68), .ZN(n487) );
  NOR2_X1 U404 ( .A1(n664), .A2(n574), .ZN(n551) );
  XNOR2_X1 U405 ( .A(n511), .B(n510), .ZN(n548) );
  XNOR2_X1 U406 ( .A(n460), .B(G469), .ZN(n461) );
  XNOR2_X1 U407 ( .A(n434), .B(n433), .ZN(n435) );
  NAND2_X1 U408 ( .A1(n637), .A2(n369), .ZN(n367) );
  NAND2_X1 U409 ( .A1(n356), .A2(n366), .ZN(n368) );
  XNOR2_X1 U410 ( .A(n365), .B(KEYINPUT64), .ZN(n414) );
  INV_X1 U411 ( .A(G131), .ZN(n365) );
  XNOR2_X1 U412 ( .A(G143), .B(G122), .ZN(n376) );
  NAND2_X1 U413 ( .A1(n729), .A2(n727), .ZN(n498) );
  OR2_X1 U414 ( .A1(n588), .A2(KEYINPUT2), .ZN(n635) );
  NOR2_X1 U415 ( .A1(n625), .A2(n502), .ZN(n533) );
  OR2_X1 U416 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U417 ( .A(n471), .B(n470), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n469), .B(n468), .ZN(n471) );
  INV_X1 U419 ( .A(KEYINPUT72), .ZN(n541) );
  NOR2_X1 U420 ( .A1(n660), .A2(n659), .ZN(n496) );
  NOR2_X1 U421 ( .A1(n466), .A2(n465), .ZN(n519) );
  INV_X1 U422 ( .A(n521), .ZN(n515) );
  XNOR2_X1 U423 ( .A(n427), .B(n426), .ZN(n430) );
  XNOR2_X1 U424 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U425 ( .A(n389), .B(n388), .ZN(n686) );
  XNOR2_X1 U426 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U427 ( .A(n454), .B(n453), .ZN(n457) );
  NAND2_X1 U428 ( .A1(n694), .A2(G210), .ZN(n595) );
  XNOR2_X1 U429 ( .A(n363), .B(n361), .ZN(n727) );
  XNOR2_X1 U430 ( .A(n497), .B(n362), .ZN(n361) );
  OR2_X1 U431 ( .A1(n512), .A2(n655), .ZN(n363) );
  INV_X1 U432 ( .A(KEYINPUT104), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n551), .B(KEYINPUT34), .ZN(n360) );
  INV_X1 U434 ( .A(KEYINPUT77), .ZN(n513) );
  XNOR2_X1 U435 ( .A(n485), .B(n484), .ZN(n503) );
  INV_X1 U436 ( .A(n503), .ZN(n370) );
  XOR2_X1 U437 ( .A(KEYINPUT13), .B(G475), .Z(n355) );
  XOR2_X1 U438 ( .A(n717), .B(n541), .Z(n356) );
  XOR2_X1 U439 ( .A(KEYINPUT74), .B(KEYINPUT35), .Z(n357) );
  INV_X1 U440 ( .A(n590), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n358), .B(n478), .ZN(n480) );
  XNOR2_X1 U442 ( .A(n358), .B(n707), .ZN(n709) );
  INV_X1 U443 ( .A(n567), .ZN(n728) );
  INV_X1 U444 ( .A(n469), .ZN(n467) );
  NOR2_X1 U445 ( .A1(n642), .A2(n643), .ZN(n371) );
  XNOR2_X1 U446 ( .A(n648), .B(KEYINPUT6), .ZN(n372) );
  XOR2_X1 U447 ( .A(n558), .B(KEYINPUT76), .Z(n373) );
  AND2_X1 U448 ( .A1(n530), .A2(n529), .ZN(n374) );
  XOR2_X1 U449 ( .A(n498), .B(KEYINPUT46), .Z(n375) );
  INV_X1 U450 ( .A(n619), .ZN(n565) );
  INV_X1 U451 ( .A(G137), .ZN(n407) );
  XNOR2_X1 U452 ( .A(n408), .B(n407), .ZN(n409) );
  INV_X1 U453 ( .A(G134), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n410), .B(n409), .ZN(n413) );
  INV_X1 U455 ( .A(KEYINPUT24), .ZN(n424) );
  XNOR2_X1 U456 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U457 ( .A(n531), .B(KEYINPUT48), .ZN(n540) );
  XNOR2_X1 U458 ( .A(n425), .B(n424), .ZN(n427) );
  INV_X1 U459 ( .A(KEYINPUT66), .ZN(n460) );
  XNOR2_X1 U460 ( .A(n398), .B(KEYINPUT95), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U462 ( .A(n505), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U463 ( .A(n436), .B(n435), .ZN(n642) );
  XNOR2_X1 U464 ( .A(n488), .B(n487), .ZN(n532) );
  XNOR2_X1 U465 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n378) );
  XNOR2_X1 U467 ( .A(G140), .B(KEYINPUT12), .ZN(n377) );
  XNOR2_X1 U468 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U469 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U470 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n382) );
  NAND2_X1 U471 ( .A1(G214), .A2(n404), .ZN(n381) );
  XNOR2_X1 U472 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U473 ( .A(n384), .B(n383), .ZN(n389) );
  XNOR2_X1 U474 ( .A(G146), .B(G125), .ZN(n472) );
  INV_X1 U475 ( .A(KEYINPUT10), .ZN(n385) );
  XNOR2_X1 U476 ( .A(n472), .B(n385), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n467), .B(n423), .ZN(n387) );
  INV_X1 U478 ( .A(G902), .ZN(n420) );
  XOR2_X1 U479 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n391) );
  XNOR2_X1 U480 ( .A(G116), .B(KEYINPUT97), .ZN(n390) );
  XNOR2_X1 U481 ( .A(n391), .B(n390), .ZN(n396) );
  XNOR2_X1 U482 ( .A(n415), .B(n394), .ZN(n395) );
  XNOR2_X1 U483 ( .A(n396), .B(n395), .ZN(n400) );
  AND2_X1 U484 ( .A1(G234), .A2(n455), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n397), .B(KEYINPUT8), .ZN(n428) );
  AND2_X1 U486 ( .A1(G217), .A2(n428), .ZN(n398) );
  INV_X1 U487 ( .A(G122), .ZN(n401) );
  XNOR2_X1 U488 ( .A(n401), .B(G107), .ZN(n470) );
  XNOR2_X1 U489 ( .A(n402), .B(n470), .ZN(n692) );
  NAND2_X1 U490 ( .A1(n692), .A2(n420), .ZN(n403) );
  XNOR2_X1 U491 ( .A(n403), .B(G478), .ZN(n522) );
  OR2_X1 U492 ( .A1(n515), .A2(n522), .ZN(n625) );
  XNOR2_X1 U493 ( .A(KEYINPUT101), .B(KEYINPUT30), .ZN(n422) );
  XOR2_X1 U494 ( .A(KEYINPUT71), .B(KEYINPUT5), .Z(n406) );
  NAND2_X1 U495 ( .A1(n404), .A2(G210), .ZN(n405) );
  XNOR2_X1 U496 ( .A(n406), .B(n405), .ZN(n410) );
  XNOR2_X1 U497 ( .A(G113), .B(KEYINPUT90), .ZN(n408) );
  XNOR2_X1 U498 ( .A(KEYINPUT3), .B(KEYINPUT67), .ZN(n411) );
  XNOR2_X1 U499 ( .A(n353), .B(n411), .ZN(n706) );
  INV_X1 U500 ( .A(G101), .ZN(n412) );
  XNOR2_X1 U501 ( .A(n412), .B(KEYINPUT4), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n706), .B(n450), .ZN(n479) );
  XOR2_X1 U503 ( .A(n413), .B(n479), .Z(n416) );
  XNOR2_X1 U504 ( .A(G146), .B(n715), .ZN(n459) );
  XNOR2_X1 U505 ( .A(n416), .B(n459), .ZN(n605) );
  NOR2_X1 U506 ( .A1(n605), .A2(G902), .ZN(n418) );
  XNOR2_X1 U507 ( .A(G472), .B(KEYINPUT69), .ZN(n417) );
  XNOR2_X2 U508 ( .A(n418), .B(n417), .ZN(n648) );
  INV_X1 U509 ( .A(G237), .ZN(n419) );
  NAND2_X1 U510 ( .A1(n420), .A2(n419), .ZN(n481) );
  NAND2_X1 U511 ( .A1(n481), .A2(G214), .ZN(n656) );
  AND2_X1 U512 ( .A1(n648), .A2(n656), .ZN(n421) );
  XNOR2_X1 U513 ( .A(n422), .B(n421), .ZN(n466) );
  XOR2_X1 U514 ( .A(G137), .B(G140), .Z(n449) );
  XNOR2_X1 U515 ( .A(n449), .B(n423), .ZN(n713) );
  XNOR2_X1 U516 ( .A(G119), .B(G110), .ZN(n425) );
  XOR2_X1 U517 ( .A(G128), .B(KEYINPUT23), .Z(n426) );
  NAND2_X1 U518 ( .A1(n428), .A2(G221), .ZN(n429) );
  XNOR2_X1 U519 ( .A(n713), .B(n431), .ZN(n695) );
  NOR2_X1 U520 ( .A1(G902), .A2(n695), .ZN(n436) );
  XNOR2_X1 U521 ( .A(KEYINPUT15), .B(G902), .ZN(n590) );
  NAND2_X1 U522 ( .A1(G234), .A2(n590), .ZN(n432) );
  XNOR2_X1 U523 ( .A(KEYINPUT20), .B(n432), .ZN(n437) );
  NAND2_X1 U524 ( .A1(G217), .A2(n437), .ZN(n434) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(KEYINPUT88), .Z(n433) );
  NAND2_X1 U526 ( .A1(n437), .A2(G221), .ZN(n440) );
  INV_X1 U527 ( .A(KEYINPUT89), .ZN(n438) );
  XNOR2_X1 U528 ( .A(n438), .B(KEYINPUT21), .ZN(n439) );
  XNOR2_X1 U529 ( .A(n440), .B(n439), .ZN(n643) );
  NAND2_X1 U530 ( .A1(G234), .A2(G237), .ZN(n441) );
  XNOR2_X1 U531 ( .A(n441), .B(KEYINPUT14), .ZN(n443) );
  NAND2_X1 U532 ( .A1(G952), .A2(n443), .ZN(n442) );
  XNOR2_X1 U533 ( .A(KEYINPUT86), .B(n442), .ZN(n673) );
  NOR2_X1 U534 ( .A1(n673), .A2(G953), .ZN(n546) );
  INV_X1 U535 ( .A(n546), .ZN(n446) );
  NAND2_X1 U536 ( .A1(G902), .A2(n443), .ZN(n544) );
  NOR2_X1 U537 ( .A1(G900), .A2(n544), .ZN(n444) );
  NAND2_X1 U538 ( .A1(G953), .A2(n444), .ZN(n445) );
  NAND2_X1 U539 ( .A1(n446), .A2(n445), .ZN(n447) );
  XOR2_X1 U540 ( .A(KEYINPUT78), .B(n447), .Z(n448) );
  NOR2_X1 U541 ( .A1(n643), .A2(n448), .ZN(n491) );
  XNOR2_X1 U542 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U543 ( .A(G104), .B(G110), .Z(n452) );
  INV_X1 U544 ( .A(G107), .ZN(n451) );
  NAND2_X1 U545 ( .A1(G227), .A2(n455), .ZN(n456) );
  XNOR2_X1 U546 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U547 ( .A(n459), .B(n458), .ZN(n682) );
  NOR2_X1 U548 ( .A1(n682), .A2(G902), .ZN(n462) );
  XNOR2_X2 U549 ( .A(n462), .B(n461), .ZN(n508) );
  NAND2_X1 U550 ( .A1(n491), .A2(n508), .ZN(n463) );
  NOR2_X1 U551 ( .A1(n642), .A2(n463), .ZN(n464) );
  XNOR2_X1 U552 ( .A(n464), .B(KEYINPUT73), .ZN(n465) );
  XNOR2_X1 U553 ( .A(KEYINPUT16), .B(G110), .ZN(n468) );
  XNOR2_X1 U554 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U555 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n475) );
  NAND2_X1 U556 ( .A1(n455), .A2(G224), .ZN(n474) );
  XNOR2_X1 U557 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U558 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U559 ( .A(n480), .B(n479), .ZN(n593) );
  NAND2_X1 U560 ( .A1(n593), .A2(n590), .ZN(n485) );
  NAND2_X1 U561 ( .A1(n481), .A2(G210), .ZN(n483) );
  INV_X1 U562 ( .A(KEYINPUT85), .ZN(n482) );
  XNOR2_X1 U563 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT38), .ZN(n657) );
  NAND2_X1 U565 ( .A1(n519), .A2(n657), .ZN(n488) );
  XOR2_X1 U566 ( .A(KEYINPUT39), .B(KEYINPUT82), .Z(n486) );
  NOR2_X1 U567 ( .A1(n625), .A2(n532), .ZN(n490) );
  XNOR2_X1 U568 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U569 ( .A(n490), .B(n489), .ZN(n729) );
  INV_X1 U570 ( .A(n642), .ZN(n500) );
  XNOR2_X1 U571 ( .A(n491), .B(KEYINPUT65), .ZN(n499) );
  INV_X1 U572 ( .A(n499), .ZN(n492) );
  NAND2_X1 U573 ( .A1(n492), .A2(n648), .ZN(n493) );
  XNOR2_X1 U574 ( .A(KEYINPUT28), .B(n494), .ZN(n495) );
  NAND2_X1 U575 ( .A1(n508), .A2(n495), .ZN(n512) );
  NAND2_X1 U576 ( .A1(n657), .A2(n656), .ZN(n660) );
  XNOR2_X1 U577 ( .A(n496), .B(KEYINPUT41), .ZN(n655) );
  XNOR2_X1 U578 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n497) );
  INV_X1 U579 ( .A(n372), .ZN(n578) );
  NOR2_X1 U580 ( .A1(n500), .A2(n499), .ZN(n501) );
  NAND2_X1 U581 ( .A1(n578), .A2(n501), .ZN(n502) );
  XOR2_X1 U582 ( .A(n533), .B(KEYINPUT106), .Z(n504) );
  NOR2_X1 U583 ( .A1(n504), .A2(n511), .ZN(n507) );
  INV_X1 U584 ( .A(KEYINPUT36), .ZN(n505) );
  NAND2_X1 U585 ( .A1(n509), .A2(n354), .ZN(n632) );
  INV_X1 U586 ( .A(KEYINPUT19), .ZN(n510) );
  OR2_X1 U587 ( .A1(n512), .A2(n548), .ZN(n514) );
  XNOR2_X2 U588 ( .A(n514), .B(n513), .ZN(n623) );
  INV_X1 U589 ( .A(n623), .ZN(n517) );
  NAND2_X1 U590 ( .A1(n522), .A2(n515), .ZN(n629) );
  NAND2_X1 U591 ( .A1(n625), .A2(n629), .ZN(n576) );
  INV_X1 U592 ( .A(n576), .ZN(n661) );
  NOR2_X1 U593 ( .A1(KEYINPUT47), .A2(n661), .ZN(n516) );
  NAND2_X1 U594 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U595 ( .A1(n632), .A2(n518), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n661), .A2(KEYINPUT47), .ZN(n524) );
  NAND2_X1 U597 ( .A1(n519), .A2(n370), .ZN(n520) );
  XOR2_X1 U598 ( .A(KEYINPUT102), .B(n520), .Z(n523) );
  AND2_X1 U599 ( .A1(n522), .A2(n521), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n523), .A2(n552), .ZN(n622) );
  NAND2_X1 U601 ( .A1(n524), .A2(n622), .ZN(n525) );
  XNOR2_X1 U602 ( .A(KEYINPUT79), .B(n525), .ZN(n528) );
  NAND2_X1 U603 ( .A1(n623), .A2(KEYINPUT47), .ZN(n526) );
  XNOR2_X1 U604 ( .A(n526), .B(KEYINPUT80), .ZN(n527) );
  AND2_X1 U605 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U606 ( .A1(n375), .A2(n374), .ZN(n531) );
  OR2_X1 U607 ( .A1(n532), .A2(n629), .ZN(n633) );
  XOR2_X1 U608 ( .A(KEYINPUT100), .B(KEYINPUT43), .Z(n537) );
  NAND2_X1 U609 ( .A1(n533), .A2(n656), .ZN(n534) );
  XNOR2_X1 U610 ( .A(n534), .B(KEYINPUT99), .ZN(n535) );
  INV_X1 U611 ( .A(n354), .ZN(n562) );
  NAND2_X1 U612 ( .A1(n535), .A2(n562), .ZN(n536) );
  XNOR2_X1 U613 ( .A(n537), .B(n536), .ZN(n538) );
  OR2_X1 U614 ( .A1(n538), .A2(n370), .ZN(n603) );
  NAND2_X1 U615 ( .A1(n633), .A2(n603), .ZN(n539) );
  NOR2_X2 U616 ( .A1(n540), .A2(n539), .ZN(n717) );
  NAND2_X1 U617 ( .A1(n640), .A2(n371), .ZN(n569) );
  XNOR2_X1 U618 ( .A(KEYINPUT33), .B(n542), .ZN(n664) );
  NOR2_X1 U619 ( .A1(G898), .A2(n455), .ZN(n543) );
  XNOR2_X1 U620 ( .A(KEYINPUT87), .B(n543), .ZN(n708) );
  NOR2_X1 U621 ( .A1(n708), .A2(n544), .ZN(n545) );
  NOR2_X1 U622 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U623 ( .A(KEYINPUT0), .ZN(n549) );
  INV_X1 U624 ( .A(n553), .ZN(n574) );
  NOR2_X1 U625 ( .A1(n659), .A2(n643), .ZN(n554) );
  NAND2_X1 U626 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U627 ( .A(KEYINPUT70), .B(KEYINPUT22), .ZN(n555) );
  XNOR2_X1 U628 ( .A(n556), .B(n555), .ZN(n579) );
  INV_X1 U629 ( .A(n579), .ZN(n559) );
  AND2_X1 U630 ( .A1(n354), .A2(n372), .ZN(n557) );
  NAND2_X1 U631 ( .A1(n642), .A2(n557), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n373), .ZN(n561) );
  XNOR2_X1 U633 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n560) );
  XNOR2_X1 U634 ( .A(n561), .B(n560), .ZN(n602) );
  NOR2_X1 U635 ( .A1(n648), .A2(n354), .ZN(n563) );
  NAND2_X1 U636 ( .A1(n563), .A2(n642), .ZN(n564) );
  OR2_X1 U637 ( .A1(n579), .A2(n564), .ZN(n619) );
  NOR2_X1 U638 ( .A1(n602), .A2(n565), .ZN(n566) );
  INV_X1 U639 ( .A(n569), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n648), .A2(n570), .ZN(n651) );
  NOR2_X1 U641 ( .A1(n651), .A2(n574), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n571), .B(KEYINPUT31), .ZN(n628) );
  INV_X1 U643 ( .A(n648), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n572), .A2(n371), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n575), .A2(n508), .ZN(n614) );
  NAND2_X1 U647 ( .A1(n628), .A2(n614), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n583) );
  OR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT83), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n354), .A2(n642), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n611) );
  AND2_X1 U653 ( .A1(n583), .A2(n611), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U655 ( .A(KEYINPUT45), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n587), .B(n586), .ZN(n588) );
  INV_X1 U657 ( .A(n588), .ZN(n699) );
  NAND2_X1 U658 ( .A1(n699), .A2(n717), .ZN(n589) );
  XNOR2_X1 U659 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT84), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n595), .B(n594), .ZN(n597) );
  INV_X1 U663 ( .A(G952), .ZN(n596) );
  AND2_X1 U664 ( .A1(n596), .A2(G953), .ZN(n698) );
  NOR2_X2 U665 ( .A1(n597), .A2(n698), .ZN(n600) );
  INV_X1 U666 ( .A(KEYINPUT119), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT56), .ZN(n599) );
  XNOR2_X1 U668 ( .A(n600), .B(n599), .ZN(G51) );
  XOR2_X1 U669 ( .A(G119), .B(KEYINPUT126), .Z(n601) );
  XNOR2_X1 U670 ( .A(n602), .B(n601), .ZN(G21) );
  XNOR2_X1 U671 ( .A(n603), .B(G140), .ZN(G42) );
  NAND2_X1 U672 ( .A1(n694), .A2(G472), .ZN(n607) );
  XNOR2_X1 U673 ( .A(KEYINPUT108), .B(KEYINPUT62), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X2 U676 ( .A1(n608), .A2(n698), .ZN(n610) );
  XNOR2_X1 U677 ( .A(KEYINPUT109), .B(KEYINPUT63), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(G57) );
  XNOR2_X1 U679 ( .A(G101), .B(KEYINPUT110), .ZN(n612) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(G3) );
  NOR2_X1 U681 ( .A1(n625), .A2(n614), .ZN(n613) );
  XOR2_X1 U682 ( .A(G104), .B(n613), .Z(G6) );
  NOR2_X1 U683 ( .A1(n614), .A2(n629), .ZN(n618) );
  XOR2_X1 U684 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n616) );
  XNOR2_X1 U685 ( .A(G107), .B(KEYINPUT26), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(G9) );
  XNOR2_X1 U688 ( .A(G110), .B(n619), .ZN(G12) );
  XOR2_X1 U689 ( .A(G128), .B(KEYINPUT29), .Z(n621) );
  OR2_X1 U690 ( .A1(n623), .A2(n629), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G30) );
  XNOR2_X1 U692 ( .A(G143), .B(n622), .ZN(G45) );
  NOR2_X1 U693 ( .A1(n625), .A2(n623), .ZN(n624) );
  XOR2_X1 U694 ( .A(G146), .B(n624), .Z(G48) );
  NOR2_X1 U695 ( .A1(n625), .A2(n628), .ZN(n626) );
  XOR2_X1 U696 ( .A(KEYINPUT112), .B(n626), .Z(n627) );
  XNOR2_X1 U697 ( .A(G113), .B(n627), .ZN(G15) );
  NOR2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U699 ( .A(G116), .B(n630), .Z(G18) );
  XOR2_X1 U700 ( .A(G125), .B(KEYINPUT37), .Z(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(G27) );
  XNOR2_X1 U702 ( .A(G134), .B(n633), .ZN(G36) );
  NOR2_X1 U703 ( .A1(KEYINPUT2), .A2(n717), .ZN(n634) );
  XOR2_X1 U704 ( .A(KEYINPUT81), .B(n634), .Z(n639) );
  INV_X1 U705 ( .A(n635), .ZN(n636) );
  NOR2_X1 U706 ( .A1(n637), .A2(n636), .ZN(n638) );
  OR2_X1 U707 ( .A1(n639), .A2(n638), .ZN(n677) );
  NOR2_X1 U708 ( .A1(n664), .A2(n655), .ZN(n675) );
  XOR2_X1 U709 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n671) );
  OR2_X1 U710 ( .A1(n354), .A2(n371), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT50), .ZN(n650) );
  XOR2_X1 U712 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n645) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(KEYINPUT113), .ZN(n647) );
  NOR2_X1 U716 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U719 ( .A(KEYINPUT51), .B(n653), .ZN(n654) );
  NOR2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n668) );
  NOR2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n663) );
  NOR2_X1 U723 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U724 ( .A1(n663), .A2(n662), .ZN(n665) );
  NOR2_X1 U725 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U726 ( .A(KEYINPUT115), .B(n666), .Z(n667) );
  NOR2_X1 U727 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U728 ( .A(n669), .B(KEYINPUT116), .ZN(n670) );
  XNOR2_X1 U729 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U730 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U732 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U733 ( .A(KEYINPUT118), .B(n678), .ZN(n679) );
  NOR2_X1 U734 ( .A1(n679), .A2(G953), .ZN(n680) );
  XNOR2_X1 U735 ( .A(n680), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U736 ( .A1(n694), .A2(G469), .ZN(n684) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  XNOR2_X1 U738 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U739 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U740 ( .A1(n698), .A2(n685), .ZN(G54) );
  NAND2_X1 U741 ( .A1(n694), .A2(G475), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n686), .B(KEYINPUT59), .ZN(n687) );
  XNOR2_X1 U743 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X2 U744 ( .A1(n689), .A2(n698), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n694), .A2(G478), .ZN(n691) );
  XOR2_X1 U747 ( .A(n692), .B(n691), .Z(n693) );
  NOR2_X1 U748 ( .A1(n698), .A2(n693), .ZN(G63) );
  NAND2_X1 U749 ( .A1(n694), .A2(G217), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U751 ( .A1(n698), .A2(n697), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n699), .A2(n455), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n700), .B(KEYINPUT120), .ZN(n704) );
  NAND2_X1 U754 ( .A1(G953), .A2(G224), .ZN(n701) );
  XNOR2_X1 U755 ( .A(KEYINPUT61), .B(n701), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n702), .A2(G898), .ZN(n703) );
  NAND2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT121), .ZN(n711) );
  XNOR2_X1 U759 ( .A(n706), .B(G101), .ZN(n707) );
  NAND2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U762 ( .A(KEYINPUT122), .B(n712), .ZN(G69) );
  XOR2_X1 U763 ( .A(n713), .B(KEYINPUT123), .Z(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U765 ( .A(KEYINPUT4), .B(n716), .ZN(n721) );
  INV_X1 U766 ( .A(n721), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(n455), .ZN(n720) );
  XNOR2_X1 U769 ( .A(KEYINPUT124), .B(n720), .ZN(n726) );
  XNOR2_X1 U770 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U772 ( .A1(G953), .A2(n723), .ZN(n724) );
  XOR2_X1 U773 ( .A(KEYINPUT125), .B(n724), .Z(n725) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(G72) );
  XNOR2_X1 U775 ( .A(n727), .B(G137), .ZN(G39) );
  XOR2_X1 U776 ( .A(n728), .B(G122), .Z(G24) );
  XOR2_X1 U777 ( .A(n729), .B(G131), .Z(n730) );
  XNOR2_X1 U778 ( .A(KEYINPUT127), .B(n730), .ZN(G33) );
endmodule

