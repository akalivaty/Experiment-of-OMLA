//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  OR2_X1    g0000(.A1(KEYINPUT64), .A2(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(KEYINPUT64), .A2(G50), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  OR3_X1    g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n208), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n222), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n217), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT67), .B(G223), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n253), .A3(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n254), .B(new_n256), .C1(new_n257), .C2(new_n252), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n260), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n259), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(G226), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n262), .A2(G190), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n226), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n216), .A2(KEYINPUT8), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT68), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(KEYINPUT68), .A3(G58), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n225), .A3(G33), .A4(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n277), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n210), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n268), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n226), .A3(new_n275), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n290), .B1(new_n210), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n274), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n273), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n262), .A2(new_n272), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n287), .A2(new_n293), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(G200), .B1(new_n297), .B2(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n297), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n305), .B(new_n306), .C1(G179), .C2(new_n296), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT70), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT69), .B(G107), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G232), .A2(G1698), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n255), .A2(G238), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n252), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n315), .A2(new_n318), .A3(new_n261), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n271), .A2(G244), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n266), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n309), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(new_n318), .A3(new_n261), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n323), .A2(KEYINPUT70), .A3(new_n266), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G190), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  INV_X1    g0127(.A(new_n278), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n327), .A2(new_n328), .B1(new_n225), .B2(new_n257), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n225), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n276), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n289), .A2(new_n257), .ZN(new_n334));
  INV_X1    g0134(.A(new_n292), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G77), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n326), .B(new_n338), .C1(new_n339), .C2(new_n325), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n325), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n322), .A2(new_n324), .A3(new_n304), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n308), .A2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT71), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n328), .A2(new_n210), .B1(new_n225), .B2(G68), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n331), .A2(new_n257), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n276), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT74), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n288), .A2(KEYINPUT12), .A3(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT12), .B1(new_n288), .B2(G68), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n354), .A2(new_n355), .B1(new_n335), .B2(G68), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n211), .A2(new_n255), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n217), .A2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n312), .C2(new_n313), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n261), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(G274), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n270), .B2(new_n259), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n271), .A2(G238), .B1(new_n367), .B2(new_n265), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n260), .B1(new_n361), .B2(new_n362), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n260), .A2(G238), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n266), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT13), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(KEYINPUT72), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n364), .A2(new_n368), .A3(new_n376), .A4(new_n365), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(G169), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n369), .A2(KEYINPUT73), .A3(new_n374), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(KEYINPUT13), .C1(new_n370), .C2(new_n373), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G179), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n375), .A2(new_n385), .A3(G169), .A4(new_n377), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT75), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n379), .A2(new_n384), .A3(KEYINPUT75), .A4(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n358), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n375), .A2(G200), .A3(new_n377), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n380), .B2(new_n382), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n357), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n314), .B2(new_n225), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n251), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G68), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n216), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n202), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n278), .A2(G159), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n277), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n250), .A2(new_n225), .A3(new_n251), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n401), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n403), .A2(new_n404), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT76), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n284), .A2(new_n292), .A3(new_n285), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n289), .B1(new_n284), .B2(new_n285), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n284), .A2(new_n292), .A3(new_n285), .ZN(new_n419));
  INV_X1    g0219(.A(new_n285), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n283), .B2(new_n327), .ZN(new_n421));
  OAI211_X1 g0221(.A(KEYINPUT76), .B(new_n419), .C1(new_n421), .C2(new_n289), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n407), .A2(new_n414), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n424));
  INV_X1    g0224(.A(G223), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n255), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n211), .A2(G1698), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n312), .C2(new_n313), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n261), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n260), .A2(G232), .A3(new_n371), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n266), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT78), .B(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT79), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n260), .B1(new_n428), .B2(new_n429), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n266), .A2(new_n432), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT79), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n434), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n431), .A2(new_n433), .A3(KEYINPUT77), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n437), .B2(new_n438), .ZN(new_n445));
  AOI21_X1  g0245(.A(G200), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n423), .B(new_n424), .C1(new_n442), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OR2_X1    g0248(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT77), .B1(new_n431), .B2(new_n433), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n437), .A2(new_n438), .A3(new_n444), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n339), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n436), .A3(new_n441), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n449), .B1(new_n453), .B2(new_n423), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n418), .A2(new_n422), .ZN(new_n456));
  INV_X1    g0256(.A(new_n413), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT16), .B1(new_n400), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n276), .B1(new_n412), .B2(new_n405), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n439), .A2(new_n341), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n304), .B1(new_n450), .B2(new_n451), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT18), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT18), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n443), .A2(new_n445), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(new_n304), .B1(new_n341), .B2(new_n439), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(new_n460), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n455), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n346), .B2(KEYINPUT71), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n347), .A2(new_n396), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G107), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n289), .B2(new_n473), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n268), .A2(G33), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n277), .A2(new_n288), .A3(new_n476), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n473), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n225), .B(G87), .C1(new_n312), .C2(new_n313), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n252), .A2(KEYINPUT22), .A3(new_n225), .A4(G87), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT23), .B1(new_n310), .B2(new_n225), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n225), .A2(KEYINPUT23), .A3(G107), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(G20), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n225), .A2(KEYINPUT84), .A3(G33), .A4(G116), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT85), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n493), .A2(new_n276), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n490), .A2(new_n491), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n490), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n478), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n499));
  OAI211_X1 g0299(.A(G250), .B(new_n255), .C1(new_n312), .C2(new_n313), .ZN(new_n500));
  INV_X1    g0300(.A(G294), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(new_n500), .C1(new_n249), .C2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n264), .A2(G1), .ZN(new_n503));
  AND2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n506), .A2(new_n260), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n502), .A2(new_n261), .B1(new_n507), .B2(G264), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT5), .B(G41), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n367), .A2(new_n503), .A3(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n508), .A2(KEYINPUT86), .A3(new_n393), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n502), .A2(new_n261), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(G264), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n512), .B1(new_n515), .B2(new_n339), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(G190), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n498), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n330), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n288), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n288), .A2(new_n476), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n522), .A2(new_n523), .A3(new_n276), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n225), .B1(new_n362), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n218), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n310), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n252), .A2(new_n225), .A3(G68), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n525), .B1(new_n331), .B2(new_n218), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n521), .B(new_n524), .C1(new_n531), .C2(new_n276), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n268), .A2(G45), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n260), .A2(G250), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n260), .A2(G274), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n533), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n537));
  OAI211_X1 g0337(.A(G238), .B(new_n255), .C1(new_n312), .C2(new_n313), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(new_n486), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n539), .B2(new_n261), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G190), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n532), .B(new_n541), .C1(new_n339), .C2(new_n540), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n531), .A2(new_n276), .ZN(new_n543));
  INV_X1    g0343(.A(new_n521), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n522), .A2(new_n276), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n520), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n341), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(G169), .C2(new_n540), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(new_n255), .C1(new_n312), .C2(new_n313), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G283), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n261), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n506), .A2(new_n260), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n510), .B1(new_n559), .B2(new_n219), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G169), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n557), .B2(new_n261), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G179), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n218), .A2(new_n473), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT81), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(KEYINPUT6), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n567), .A2(new_n568), .ZN(new_n571));
  MUX2_X1   g0371(.A(new_n569), .B(G97), .S(KEYINPUT6), .Z(new_n572));
  OAI211_X1 g0372(.A(G20), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n278), .A2(G77), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n311), .B1(new_n411), .B2(new_n398), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(KEYINPUT82), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(KEYINPUT82), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n276), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n288), .A2(G97), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n545), .B2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n566), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n562), .A2(G190), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n564), .A2(G200), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n578), .B(new_n580), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n550), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n515), .A2(new_n304), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G179), .B2(new_n515), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n494), .A2(new_n497), .ZN(new_n589));
  INV_X1    g0389(.A(new_n478), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n592));
  OAI211_X1 g0392(.A(G257), .B(new_n255), .C1(new_n312), .C2(new_n313), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n250), .A2(G303), .A3(new_n251), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT83), .A4(new_n594), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n261), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n510), .B1(new_n559), .B2(new_n213), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n434), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n260), .B1(new_n595), .B2(new_n596), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n604), .B2(new_n598), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n339), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n275), .A2(new_n226), .B1(G20), .B2(new_n212), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n555), .B(new_n225), .C1(G33), .C2(new_n218), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT20), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n608), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n288), .A2(G116), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n545), .B2(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n603), .A2(new_n606), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n608), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n609), .ZN(new_n619));
  INV_X1    g0419(.A(new_n613), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n477), .B2(new_n212), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n617), .B1(new_n605), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n304), .B1(new_n612), .B2(new_n614), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n602), .A2(new_n624), .A3(KEYINPUT21), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n605), .A2(G179), .A3(new_n615), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n591), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n472), .A2(new_n519), .A3(new_n586), .A4(new_n628), .ZN(G372));
  NOR2_X1   g0429(.A1(new_n395), .A2(new_n344), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n455), .B1(new_n391), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n469), .B1(new_n300), .B2(new_n302), .ZN(new_n632));
  INV_X1    g0432(.A(new_n307), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT89), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n632), .A2(KEYINPUT89), .A3(new_n633), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n566), .A2(new_n638), .B1(new_n578), .B2(new_n580), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n563), .A2(KEYINPUT88), .A3(new_n565), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n550), .A4(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n549), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n566), .A2(new_n581), .A3(new_n549), .A4(new_n542), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n627), .A2(KEYINPUT87), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n623), .A2(new_n625), .A3(new_n626), .A4(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n591), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n519), .A2(new_n582), .A3(new_n585), .A4(new_n550), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n642), .B(new_n645), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n472), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n637), .A2(new_n652), .ZN(G369));
  NAND3_X1  g0453(.A1(new_n268), .A2(new_n225), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n615), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n646), .B2(new_n648), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n616), .B(new_n661), .C1(new_n627), .C2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n589), .A2(new_n590), .ZN(new_n663));
  INV_X1    g0463(.A(new_n588), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n659), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n519), .ZN(new_n666));
  INV_X1    g0466(.A(new_n591), .ZN(new_n667));
  INV_X1    g0467(.A(new_n659), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n662), .A2(G330), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n627), .A2(new_n668), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n665), .A3(new_n519), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT90), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n659), .B(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n591), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n672), .A2(KEYINPUT91), .A3(new_n676), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n670), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n228), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G1), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n310), .A2(G116), .A3(new_n527), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n223), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n651), .A2(new_n675), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n566), .A2(new_n638), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n641), .A3(new_n581), .ZN(new_n694));
  INV_X1    g0494(.A(new_n550), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT26), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n549), .B(KEYINPUT93), .Z(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n627), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n650), .B1(new_n700), .B2(new_n667), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT29), .B(new_n668), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n692), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n628), .A2(new_n586), .A3(new_n519), .A4(new_n675), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n540), .A2(G179), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n602), .A2(new_n562), .A3(new_n706), .A4(new_n515), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n508), .A2(new_n540), .A3(KEYINPUT92), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT92), .B1(new_n508), .B2(new_n540), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n605), .A2(G179), .A3(new_n564), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n508), .A2(new_n540), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT92), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n508), .A2(new_n540), .A3(KEYINPUT92), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n711), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n707), .B1(new_n712), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  INV_X1    g0523(.A(new_n707), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT30), .B1(new_n710), .B2(new_n711), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n718), .A2(new_n719), .A3(new_n713), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n723), .B1(new_n727), .B2(new_n668), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n705), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n704), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n689), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(G13), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n268), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n684), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n226), .B1(G20), .B2(new_n304), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n393), .A2(G179), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n225), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n225), .A2(new_n341), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n434), .ZN(new_n747));
  AOI22_X1  g0547(.A1(G294), .A2(new_n744), .B1(new_n747), .B2(G326), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n339), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n434), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G322), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n225), .A2(G179), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n393), .A3(new_n339), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n252), .B1(new_n755), .B2(G329), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n746), .A2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(KEYINPUT33), .B(G317), .Z(new_n759));
  NOR2_X1   g0559(.A1(new_n750), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n753), .A2(new_n393), .A3(G200), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(G303), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n749), .A2(new_n752), .A3(new_n756), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n751), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n771), .A2(new_n216), .B1(new_n761), .B2(new_n257), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n758), .A2(new_n401), .B1(new_n473), .B2(new_n765), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n766), .A2(new_n523), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n314), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n754), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n743), .A2(new_n218), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G50), .B2(new_n747), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n774), .A2(new_n777), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n741), .B1(new_n770), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n740), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n683), .A2(new_n314), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G355), .B1(new_n212), .B2(new_n683), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n243), .A2(G45), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n683), .A2(new_n252), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n224), .B2(G45), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n739), .B(new_n784), .C1(new_n788), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n787), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n662), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n662), .A2(G330), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n739), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n662), .A2(G330), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(G396));
  NOR2_X1   g0603(.A1(new_n740), .A2(new_n785), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n739), .B1(new_n257), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n252), .B1(new_n754), .B2(new_n806), .C1(new_n743), .C2(new_n216), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n210), .A2(new_n766), .B1(new_n765), .B2(new_n401), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n747), .A2(G137), .B1(new_n760), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G143), .ZN(new_n810));
  INV_X1    g0610(.A(G150), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n771), .C1(new_n811), .C2(new_n758), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT34), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n807), .B(new_n808), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n765), .A2(new_n523), .B1(new_n754), .B2(new_n762), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  AOI22_X1  g0617(.A1(new_n747), .A2(G303), .B1(new_n760), .B2(G116), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n764), .B2(new_n758), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n771), .A2(new_n501), .B1(new_n473), .B2(new_n766), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n819), .A2(new_n820), .A3(new_n252), .A4(new_n781), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n814), .A2(new_n815), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n337), .A2(new_n659), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n340), .A2(new_n824), .B1(new_n343), .B2(new_n342), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n344), .A2(new_n659), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n805), .B1(new_n741), .B2(new_n822), .C1(new_n827), .C2(new_n786), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n825), .A2(new_n826), .A3(new_n674), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n651), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n690), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n827), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n738), .B1(new_n832), .B2(new_n730), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n730), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(G384));
  NOR3_X1   g0636(.A1(new_n226), .A2(new_n225), .A3(new_n212), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT35), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT36), .Z(new_n842));
  NAND2_X1  g0642(.A1(new_n201), .A2(new_n203), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n401), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n402), .A2(new_n223), .A3(new_n257), .ZN(new_n845));
  OAI211_X1 g0645(.A(G1), .B(new_n734), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT100), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n705), .A2(new_n850), .A3(new_n728), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n389), .A2(new_n390), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n357), .B(new_n659), .C1(new_n852), .C2(new_n395), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n358), .A2(new_n668), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n391), .A2(new_n395), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n827), .B(new_n851), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n657), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n460), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n455), .B2(new_n469), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n859), .B2(KEYINPUT101), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n423), .B1(new_n442), .B2(new_n446), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(new_n463), .A3(new_n863), .A4(new_n859), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n463), .A3(new_n859), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n407), .A2(new_n414), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n657), .B1(new_n866), .B2(new_n456), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n860), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n865), .B(new_n862), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n436), .A2(new_n441), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n460), .B1(new_n875), .B2(new_n452), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n447), .B1(new_n876), .B2(new_n449), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n463), .A2(KEYINPUT18), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n467), .A2(new_n465), .A3(new_n460), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n867), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n849), .B1(new_n857), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n851), .A2(new_n827), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n865), .A2(new_n861), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n863), .A2(new_n463), .A3(KEYINPUT37), .A4(new_n859), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT102), .B1(new_n448), .B2(new_n454), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n447), .C1(new_n876), .C2(new_n449), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n469), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n893), .B2(new_n867), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n886), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n341), .B1(new_n380), .B2(new_n382), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n375), .A2(G169), .A3(new_n377), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n385), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT75), .B1(new_n898), .B2(new_n379), .ZN(new_n899));
  INV_X1    g0699(.A(new_n390), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n357), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n395), .ZN(new_n902));
  INV_X1    g0702(.A(new_n855), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n853), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n885), .A2(new_n895), .A3(KEYINPUT40), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n884), .A2(G330), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n472), .A2(G330), .A3(new_n851), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n884), .A2(new_n906), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n472), .A2(new_n851), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n911), .B(new_n912), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n703), .A2(new_n472), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n637), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n901), .A2(new_n659), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n886), .C1(new_n894), .C2(KEYINPUT38), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT39), .B1(new_n873), .B2(new_n882), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n919), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n883), .ZN(new_n928));
  INV_X1    g0728(.A(new_n826), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n830), .A2(new_n929), .B1(new_n904), .B2(new_n853), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n928), .A2(new_n930), .B1(new_n880), .B2(new_n657), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n918), .B(new_n932), .Z(new_n933));
  OAI22_X1  g0733(.A1(new_n916), .A2(new_n933), .B1(new_n268), .B2(new_n735), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n916), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n848), .B1(new_n934), .B2(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n581), .A2(new_n674), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n582), .A2(new_n585), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT106), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n639), .A2(new_n641), .A3(new_n674), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n672), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT42), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n582), .B1(new_n941), .B2(new_n667), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n675), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n550), .B1(new_n532), .B2(new_n668), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n549), .A2(new_n532), .A3(new_n668), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n670), .A2(new_n941), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n943), .A2(new_n951), .A3(new_n950), .A4(new_n945), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n684), .B(KEYINPUT41), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n939), .A2(new_n940), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n681), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT45), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n681), .A2(new_n961), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n670), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n799), .B(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n731), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n963), .A2(new_n965), .A3(new_n670), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n960), .B1(new_n973), .B2(new_n732), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n959), .B1(new_n974), .B2(new_n737), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n751), .A2(G150), .B1(new_n760), .B2(new_n843), .ZN(new_n976));
  INV_X1    g0776(.A(G137), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n252), .B1(new_n754), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n766), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(G58), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G68), .A2(new_n744), .B1(new_n757), .B2(G159), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n765), .A2(new_n257), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n747), .B2(G143), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n976), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n765), .A2(new_n218), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n252), .B(new_n985), .C1(G317), .C2(new_n755), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n744), .A2(new_n310), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n751), .A2(G303), .B1(new_n757), .B2(G294), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT108), .B(G311), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n747), .A2(new_n989), .B1(new_n760), .B2(G283), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT109), .B1(new_n979), .B2(G116), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT46), .Z(new_n993));
  OAI21_X1  g0793(.A(new_n984), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT110), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT47), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n741), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n996), .B2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n793), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n788), .B1(new_n228), .B2(new_n330), .C1(new_n239), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n738), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT107), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n998), .B(new_n1002), .C1(new_n797), .C2(new_n949), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT111), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n975), .A2(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n970), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n737), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n747), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n210), .A2(new_n771), .B1(new_n1009), .B2(new_n778), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G68), .B2(new_n760), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n421), .A2(new_n757), .ZN(new_n1012));
  XOR2_X1   g0812(.A(KEYINPUT112), .B(G150), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n252), .B1(new_n1013), .B2(new_n754), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n985), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n744), .A2(new_n520), .B1(new_n979), .B2(G77), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G303), .A2(new_n760), .B1(new_n757), .B2(new_n989), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n751), .A2(G317), .ZN(new_n1019));
  XOR2_X1   g0819(.A(KEYINPUT113), .B(G322), .Z(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1019), .C1(new_n1009), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n743), .A2(new_n764), .B1(new_n766), .B2(new_n501), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n252), .B1(new_n755), .B2(G326), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n212), .C2(new_n765), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1017), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n740), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n236), .A2(new_n264), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(new_n793), .B1(new_n687), .B2(new_n790), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n327), .A2(G50), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT50), .Z(new_n1035));
  OAI21_X1  g0835(.A(new_n264), .B1(new_n401), .B2(new_n257), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1035), .A2(new_n687), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1033), .A2(new_n1037), .B1(G107), .B2(new_n228), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n739), .B1(new_n1038), .B2(new_n788), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1031), .B(new_n1039), .C1(new_n669), .C2(new_n797), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1008), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n971), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n684), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n732), .A2(new_n1007), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G393));
  INV_X1    g0845(.A(new_n972), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n670), .B1(new_n963), .B2(new_n965), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n973), .A3(new_n684), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n968), .A2(new_n737), .A3(new_n972), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n246), .A2(new_n793), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n740), .B(new_n787), .C1(G97), .C2(new_n683), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n739), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G311), .A2(new_n751), .B1(new_n747), .B2(G317), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  AOI22_X1  g0855(.A1(G116), .A2(new_n744), .B1(new_n760), .B2(G294), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n767), .B2(new_n758), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n754), .A2(new_n1020), .B1(new_n766), .B2(new_n764), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n314), .B1(new_n765), .B2(new_n473), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G150), .A2(new_n747), .B1(new_n751), .B2(G159), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT51), .Z(new_n1063));
  OAI22_X1  g0863(.A1(new_n761), .A2(new_n327), .B1(new_n766), .B2(new_n401), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n757), .A2(new_n843), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n257), .B2(new_n743), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n252), .B1(new_n754), .B2(new_n810), .C1(new_n523), .C2(new_n765), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1055), .A2(new_n1061), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1053), .B1(new_n741), .B2(new_n1069), .C1(new_n961), .C2(new_n797), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1049), .A2(new_n1050), .A3(new_n1070), .ZN(G390));
  NAND2_X1  g0871(.A1(new_n921), .A2(new_n922), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT103), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n919), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n905), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n826), .B1(new_n651), .B2(new_n829), .ZN(new_n1076));
  OAI211_X1 g0876(.A(KEYINPUT116), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT116), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n930), .B2(new_n919), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n924), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n895), .A2(new_n1074), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT115), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n905), .B(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n825), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n668), .B(new_n1084), .C1(new_n699), .C2(new_n701), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n929), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1080), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n885), .A2(G330), .A3(new_n905), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n729), .A2(G330), .A3(new_n827), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n905), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1080), .A2(new_n1095), .A3(new_n1088), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1076), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1075), .A2(new_n1093), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1090), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1086), .B1(new_n1094), .B2(new_n905), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n851), .A2(G330), .A3(new_n827), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n905), .A2(new_n1082), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT115), .B1(new_n904), .B2(new_n853), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1098), .A2(new_n1100), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n908), .B(new_n917), .C1(new_n635), .C2(new_n636), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1097), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1092), .A2(new_n1108), .A3(new_n1096), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n684), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1073), .A2(new_n785), .A3(new_n924), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n804), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n738), .B1(new_n421), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1013), .A2(new_n766), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n843), .A2(new_n393), .A3(G200), .A4(new_n753), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n314), .B1(new_n755), .B2(G125), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G137), .A2(new_n757), .B1(new_n760), .B2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1125), .A2(KEYINPUT117), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(KEYINPUT117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n747), .A2(G128), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G159), .A2(new_n744), .B1(new_n751), .B2(G132), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n252), .B(new_n775), .C1(G294), .C2(new_n755), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n401), .B2(new_n765), .C1(new_n257), .C2(new_n743), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n751), .A2(G116), .B1(new_n757), .B2(new_n310), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n218), .B2(new_n761), .C1(new_n764), .C2(new_n1009), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1122), .A2(new_n1130), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1115), .B1(new_n1135), .B2(new_n740), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT119), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1080), .A2(new_n1095), .A3(new_n1088), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1090), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1138), .B1(new_n1141), .B2(new_n737), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1112), .A2(new_n1142), .ZN(G378));
  AOI21_X1  g0943(.A(new_n1107), .B1(new_n1141), .B2(new_n1108), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n297), .A2(new_n657), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n308), .B(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n907), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1148), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1150), .A2(new_n884), .A3(G330), .A4(new_n906), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n927), .A3(new_n931), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1149), .A2(new_n1151), .B1(new_n927), .B2(new_n931), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT122), .B1(new_n1144), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1107), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1111), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT122), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1152), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .A4(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1111), .A2(new_n1157), .B1(new_n1160), .B2(new_n1152), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n684), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n736), .B1(new_n1160), .B2(new_n1152), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n738), .B1(new_n843), .B2(new_n1114), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1150), .A2(new_n786), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n314), .B2(new_n263), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n263), .B(new_n314), .C1(new_n754), .C2(new_n764), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G68), .B2(new_n744), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n765), .A2(new_n216), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n747), .B2(G116), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n751), .A2(G107), .B1(new_n757), .B2(G97), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n760), .A2(new_n520), .B1(new_n979), .B2(G77), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1171), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n755), .C2(G124), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n747), .A2(G125), .B1(new_n760), .B2(G137), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n806), .B2(new_n758), .C1(new_n811), .C2(new_n743), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n751), .A2(G128), .B1(new_n979), .B2(new_n1124), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT59), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1181), .B1(new_n778), .B2(new_n765), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1180), .B1(new_n1179), .B2(new_n1178), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1168), .B(new_n1169), .C1(new_n740), .C2(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT121), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT121), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1167), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1166), .A2(new_n1196), .ZN(G375));
  INV_X1    g0997(.A(new_n960), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1109), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1083), .A2(new_n785), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n738), .B1(G68), .B2(new_n1114), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n751), .A2(G283), .B1(new_n760), .B2(new_n310), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n212), .B2(new_n758), .C1(new_n501), .C2(new_n1009), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n252), .B(new_n982), .C1(G303), .C2(new_n755), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n218), .B2(new_n766), .C1(new_n330), .C2(new_n743), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n314), .B(new_n1174), .C1(G128), .C2(new_n755), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n806), .B2(new_n1009), .C1(new_n758), .C2(new_n1123), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n760), .A2(G150), .B1(new_n979), .B2(G159), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n210), .B2(new_n743), .C1(new_n977), .C2(new_n771), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1204), .A2(new_n1206), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1202), .B1(new_n1211), .B2(new_n740), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n1201), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1106), .B2(new_n736), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1200), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT124), .ZN(G381));
  INV_X1    g1018(.A(G375), .ZN(new_n1219));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  INV_X1    g1020(.A(G390), .ZN(new_n1221));
  INV_X1    g1021(.A(G384), .ZN(new_n1222));
  INV_X1    g1022(.A(G396), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n1041), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1222), .A3(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1226), .A2(G381), .A3(G387), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1219), .A2(new_n1220), .A3(new_n1227), .ZN(G407));
  NAND2_X1  g1028(.A1(new_n658), .A2(G213), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1219), .A2(new_n1220), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(new_n1231), .A3(G213), .ZN(G409));
  OAI211_X1 g1032(.A(G378), .B(new_n1196), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1164), .A2(new_n1198), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1167), .A2(new_n1193), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1220), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1199), .B1(new_n1108), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT60), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n684), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1216), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1222), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(G384), .A3(new_n1216), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1237), .A2(new_n1229), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT62), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1237), .A2(new_n1229), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(G2897), .A3(new_n1230), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1230), .A2(G2897), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1243), .A2(new_n1244), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1230), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1246), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1248), .A2(new_n1255), .A3(new_n1256), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1224), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT125), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n975), .A2(new_n1005), .A3(G390), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n975), .B2(new_n1005), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G387), .A2(new_n1221), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n975), .A2(G390), .A3(new_n1005), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1261), .A2(new_n1269), .A3(new_n1224), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1260), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1273), .B(new_n1256), .C1(new_n1257), .C2(new_n1253), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1247), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1247), .B2(new_n1278), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1257), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1246), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1277), .A2(new_n1279), .A3(new_n1281), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1275), .A2(new_n1283), .ZN(G405));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1166), .B2(new_n1196), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1233), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1246), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1273), .A2(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1286), .A2(new_n1287), .A3(new_n1246), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1285), .B(new_n1274), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1286), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1233), .A3(new_n1245), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1274), .A2(new_n1285), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1289), .A4(new_n1288), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(G402));
endmodule


