//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n644,
    new_n645, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  AOI22_X1  g031(.A1(new_n451), .A2(G567), .B1(new_n453), .B2(G2106), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n473), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G124), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(G136), .A3(new_n466), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n483), .A3(KEYINPUT69), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT68), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(new_n476), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n485), .B1(new_n489), .B2(new_n482), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n484), .A2(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G138), .B(new_n466), .C1(new_n459), .C2(new_n460), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT70), .A2(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT70), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(G2104), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n474), .A2(KEYINPUT4), .A3(G138), .A4(new_n466), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n474), .A2(G126), .A3(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n494), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n505), .A2(new_n507), .A3(G50), .A4(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G50), .A4(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n505), .B(new_n507), .C1(new_n515), .C2(new_n516), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n513), .A2(new_n520), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n510), .A2(G51), .A3(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n521), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT72), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(G168));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n528), .B2(new_n529), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g123(.A(KEYINPUT73), .B(new_n546), .C1(new_n517), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT74), .B(G90), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n505), .A2(new_n507), .A3(G543), .ZN(new_n552));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n521), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G171));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT76), .B(G43), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n521), .A2(new_n558), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n504), .ZN(new_n563));
  OAI21_X1  g138(.A(G56), .B1(new_n515), .B2(new_n516), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n566), .A2(KEYINPUT75), .A3(G651), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n560), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND4_X1  g149(.A1(new_n505), .A2(new_n507), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n510), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n522), .A2(G91), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n504), .C2(new_n581), .ZN(G299));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n550), .A2(new_n583), .A3(new_n555), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n583), .B1(new_n550), .B2(new_n555), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G301));
  NAND3_X1  g162(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(G286));
  NAND2_X1  g163(.A1(new_n522), .A2(G87), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n590));
  INV_X1    g165(.A(new_n552), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n528), .B2(new_n529), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G86), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT80), .B1(new_n521), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n591), .A2(G48), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n530), .A2(new_n510), .A3(new_n603), .A4(G86), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n604), .ZN(G305));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  INV_X1    g181(.A(G47), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT81), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G47), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n521), .A2(new_n606), .B1(new_n552), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(G60), .B1(new_n515), .B2(new_n516), .ZN(new_n613));
  NAND2_X1  g188(.A1(G72), .A2(G543), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n504), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G60), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n528), .B2(new_n529), .ZN(new_n618));
  INV_X1    g193(.A(new_n614), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n530), .A2(new_n510), .A3(G85), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n510), .A2(G543), .A3(new_n608), .A4(new_n610), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n624), .ZN(G290));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n629));
  INV_X1    g204(.A(G92), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n521), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n628), .A2(new_n631), .B1(G54), .B2(new_n591), .ZN(new_n632));
  INV_X1    g207(.A(G66), .ZN(new_n633));
  INV_X1    g208(.A(G79), .ZN(new_n634));
  OAI22_X1  g209(.A1(new_n517), .A2(new_n633), .B1(new_n634), .B2(new_n527), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI221_X1 g212(.A(KEYINPUT84), .B1(new_n634), .B2(new_n527), .C1(new_n517), .C2(new_n633), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G651), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n626), .A2(KEYINPUT83), .B1(new_n627), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(KEYINPUT83), .B2(new_n626), .ZN(G284));
  OAI21_X1  g217(.A(new_n641), .B1(KEYINPUT83), .B2(new_n626), .ZN(G321));
  NOR2_X1   g218(.A1(G286), .A2(new_n627), .ZN(new_n644));
  XOR2_X1   g219(.A(G299), .B(KEYINPUT85), .Z(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(new_n627), .ZN(G297));
  AOI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n627), .ZN(G280));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(G860), .ZN(G148));
  INV_X1    g225(.A(new_n560), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT75), .B1(new_n566), .B2(G651), .ZN(new_n652));
  AOI211_X1 g227(.A(new_n561), .B(new_n504), .C1(new_n564), .C2(new_n565), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n627), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n640), .A2(G559), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n655), .B1(new_n656), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g232(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g233(.A1(new_n474), .A2(new_n466), .ZN(new_n659));
  INV_X1    g234(.A(G2104), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n659), .A2(KEYINPUT12), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(KEYINPUT12), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT13), .ZN(new_n664));
  INV_X1    g239(.A(G2100), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n488), .A2(new_n476), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G123), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n461), .A2(G2105), .ZN(new_n670));
  OR2_X1    g245(.A1(G99), .A2(G2105), .ZN(new_n671));
  INV_X1    g246(.A(G111), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n660), .B1(new_n672), .B2(G2105), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n670), .A2(G135), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n666), .A2(new_n667), .A3(new_n677), .ZN(G156));
  INV_X1    g253(.A(G14), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT15), .B(G2435), .ZN(new_n680));
  INV_X1    g255(.A(G2438), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2427), .B(G2430), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT87), .B(KEYINPUT14), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G2443), .B(G2446), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2451), .B(G2454), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n687), .A2(new_n688), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n687), .A2(new_n688), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1341), .B(G1348), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT88), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n679), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n699), .B2(new_n702), .ZN(new_n706));
  AOI211_X1 g281(.A(KEYINPUT89), .B(new_n703), .C1(new_n694), .C2(new_n698), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G401));
  XNOR2_X1  g284(.A(G2072), .B(G2078), .ZN(new_n710));
  XNOR2_X1  g285(.A(G2067), .B(G2678), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n713));
  XOR2_X1   g288(.A(G2084), .B(G2090), .Z(new_n714));
  OR3_X1    g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(new_n711), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n710), .B(KEYINPUT17), .Z(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n714), .A2(new_n710), .A3(new_n711), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT18), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n714), .A3(new_n717), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(new_n676), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G2100), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(G2096), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(new_n665), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(G227));
  XNOR2_X1  g303(.A(G1991), .B(G1996), .ZN(new_n729));
  INV_X1    g304(.A(G1981), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(G1971), .B(G1976), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT19), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(G1956), .B(G2474), .Z(new_n736));
  XOR2_X1   g311(.A(G1961), .B(G1966), .Z(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT20), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n736), .A2(new_n737), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n735), .A2(new_n738), .A3(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G1986), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n739), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n742), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G1986), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n745), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n753), .B1(new_n745), .B2(new_n751), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n732), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n745), .A2(new_n751), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(new_n752), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n759), .A2(new_n731), .A3(new_n754), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(G229));
  INV_X1    g336(.A(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G23), .ZN(new_n763));
  INV_X1    g338(.A(G288), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n762), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT33), .B(G1976), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n762), .A2(G22), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G166), .B2(new_n762), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(G1971), .B2(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G6), .B(G305), .S(G16), .Z(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n773), .C1(G1971), .C2(new_n769), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT34), .ZN(new_n776));
  INV_X1    g351(.A(G290), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G16), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G16), .B2(G24), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(new_n750), .ZN(new_n780));
  INV_X1    g355(.A(G29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G25), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n668), .A2(G119), .ZN(new_n783));
  OR2_X1    g358(.A1(G95), .A2(G2105), .ZN(new_n784));
  INV_X1    g359(.A(G107), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n660), .B1(new_n785), .B2(G2105), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n670), .A2(G131), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n782), .B1(new_n789), .B2(new_n781), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n790), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n779), .A2(new_n750), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n780), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n775), .A2(new_n776), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT36), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(G28), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n781), .B1(new_n798), .B2(G28), .ZN(new_n800));
  AND2_X1   g375(.A1(KEYINPUT31), .A2(G11), .ZN(new_n801));
  NOR2_X1   g376(.A1(KEYINPUT31), .A2(G11), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n675), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G29), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n781), .A2(G32), .ZN(new_n808));
  INV_X1    g383(.A(G129), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n488), .B2(new_n476), .ZN(new_n810));
  NAND3_X1  g385(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n474), .A2(G141), .A3(new_n466), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n808), .B1(new_n817), .B2(new_n781), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT27), .B(G1996), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n670), .A2(G139), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT93), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n466), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT25), .Z(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n781), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n781), .B2(G33), .ZN(new_n830));
  INV_X1    g405(.A(G2072), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n807), .B(new_n820), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n762), .A2(G5), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G171), .B2(new_n762), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(G1961), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n762), .A2(G21), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G168), .B2(new_n762), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G1966), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(G1961), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(G1966), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n805), .A2(new_n806), .ZN(new_n842));
  AND2_X1   g417(.A1(KEYINPUT24), .A2(G34), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n781), .B1(KEYINPUT24), .B2(G34), .ZN(new_n844));
  OAI22_X1  g419(.A1(G160), .A2(new_n781), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(G2084), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G2084), .B2(new_n845), .ZN(new_n847));
  NOR4_X1   g422(.A1(new_n832), .A2(new_n840), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n830), .A2(new_n831), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT94), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n781), .A2(G27), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G164), .B2(new_n781), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(G2078), .Z(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n848), .A2(KEYINPUT97), .A3(new_n850), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(G29), .A2(G35), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G162), .B2(G29), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT29), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G2090), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n762), .A2(G4), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n648), .B2(new_n762), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT91), .B(G1348), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT92), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n864), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n762), .A2(G20), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT23), .ZN(new_n869));
  INV_X1    g444(.A(G299), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n762), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G1956), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n762), .A2(G19), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n568), .B2(new_n762), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G1341), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n781), .A2(G26), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT28), .ZN(new_n877));
  INV_X1    g452(.A(G128), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n488), .B2(new_n476), .ZN(new_n879));
  INV_X1    g454(.A(G116), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n660), .B1(new_n880), .B2(G2105), .ZN(new_n881));
  OR2_X1    g456(.A1(G104), .A2(G2105), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G140), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n659), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n877), .B1(new_n886), .B2(new_n781), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G2067), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n872), .A2(new_n875), .A3(new_n888), .ZN(new_n889));
  AND4_X1   g464(.A1(new_n857), .A2(new_n862), .A3(new_n867), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n848), .A2(new_n850), .A3(new_n856), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n797), .A2(new_n890), .A3(new_n893), .ZN(G150));
  INV_X1    g469(.A(G150), .ZN(G311));
  NAND4_X1  g470(.A1(new_n505), .A2(new_n507), .A3(G55), .A4(G543), .ZN(new_n896));
  XOR2_X1   g471(.A(KEYINPUT98), .B(G93), .Z(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n521), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(G67), .B1(new_n515), .B2(new_n516), .ZN(new_n899));
  NAND2_X1  g474(.A1(G80), .A2(G543), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n504), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G860), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n648), .A2(G559), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT38), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n898), .B2(new_n901), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT100), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n902), .A2(KEYINPUT99), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n908), .B(new_n912), .C1(new_n898), .C2(new_n901), .ZN(new_n913));
  AND4_X1   g488(.A1(new_n568), .A2(new_n910), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n910), .A2(new_n913), .B1(new_n568), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n907), .B(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n903), .B1(new_n918), .B2(KEYINPUT39), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n905), .B1(new_n919), .B2(new_n920), .ZN(G145));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n923));
  OAI21_X1  g498(.A(G129), .B1(new_n475), .B2(new_n477), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n923), .B(new_n924), .C1(new_n879), .C2(new_n885), .ZN(new_n925));
  OAI21_X1  g500(.A(G128), .B1(new_n475), .B2(new_n477), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n670), .A2(G140), .B1(new_n882), .B2(new_n881), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n926), .B(new_n927), .C1(new_n810), .C2(new_n816), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n928), .A3(G164), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G164), .B1(new_n925), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n828), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT102), .B(new_n828), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n925), .A2(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n502), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n827), .A3(new_n929), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT103), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n937), .A2(new_n940), .A3(new_n827), .A4(new_n929), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n934), .A2(new_n935), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G142), .ZN(new_n943));
  NOR2_X1   g518(.A1(G106), .A2(G2105), .ZN(new_n944));
  OAI21_X1  g519(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n659), .A2(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(G130), .B2(new_n668), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(new_n663), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(new_n788), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n484), .A2(new_n490), .A3(new_n471), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n471), .B1(new_n484), .B2(new_n490), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT101), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT69), .B1(new_n478), .B2(new_n483), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n489), .A2(new_n485), .A3(new_n482), .ZN(new_n954));
  OAI21_X1  g529(.A(G160), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n484), .A2(new_n490), .A3(new_n471), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n952), .A2(new_n804), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n804), .B1(new_n952), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n949), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n948), .B(new_n789), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT101), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n675), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n952), .A2(new_n804), .A3(new_n958), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n942), .A2(new_n961), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT104), .B(G37), .Z(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n942), .B1(new_n961), .B2(new_n967), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n922), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n961), .A2(new_n967), .ZN(new_n973));
  INV_X1    g548(.A(new_n942), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(KEYINPUT105), .A3(new_n969), .A4(new_n968), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g553(.A1(G303), .A2(G305), .ZN(new_n979));
  NOR2_X1   g554(.A1(G303), .A2(G305), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n616), .A2(new_n983), .A3(new_n624), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n616), .B2(new_n624), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n984), .A2(new_n985), .A3(G288), .ZN(new_n986));
  NAND2_X1  g561(.A1(G290), .A2(KEYINPUT107), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n616), .A2(new_n983), .A3(new_n624), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n764), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n982), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(G288), .B1(new_n984), .B2(new_n985), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n987), .A2(new_n764), .A3(new_n988), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(KEYINPUT108), .A3(new_n982), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n993), .A2(new_n994), .A3(new_n999), .A4(new_n981), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n992), .A2(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(KEYINPUT110), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(KEYINPUT110), .B2(new_n1002), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n916), .B(new_n656), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n640), .A2(new_n870), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G299), .B1(new_n639), .B2(new_n632), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT106), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n632), .A2(G299), .A3(new_n639), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n1009), .B2(KEYINPUT106), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n640), .A2(KEYINPUT106), .A3(new_n870), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT41), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT41), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1008), .A2(new_n1010), .A3(new_n1018), .A4(new_n1011), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1014), .B1(new_n1021), .B2(new_n1005), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n998), .A2(new_n1000), .ZN(new_n1023));
  INV_X1    g598(.A(new_n996), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT108), .B1(new_n995), .B2(new_n982), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n1026), .A2(KEYINPUT110), .A3(new_n1002), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1004), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n1004), .B2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g604(.A(G868), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(G868), .B2(new_n902), .ZN(G295));
  OAI21_X1  g606(.A(new_n1030), .B1(G868), .B2(new_n902), .ZN(G331));
  OAI21_X1  g607(.A(G168), .B1(new_n585), .B2(new_n586), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G286), .A2(new_n556), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1033), .B(new_n1034), .C1(new_n914), .C2(new_n915), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n910), .A2(new_n568), .A3(new_n911), .A4(new_n913), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT98), .B(G93), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n530), .A2(new_n510), .A3(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n899), .A2(new_n900), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n896), .B(new_n1038), .C1(new_n1039), .C2(new_n504), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n912), .B1(new_n1040), .B2(new_n908), .ZN(new_n1041));
  INV_X1    g616(.A(new_n913), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n908), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1041), .A2(new_n1042), .B1(new_n1043), .B2(new_n654), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n556), .A2(KEYINPUT78), .ZN(new_n1045));
  AOI21_X1  g620(.A(G286), .B1(new_n1045), .B2(new_n584), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1034), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1036), .B(new_n1044), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1035), .A2(new_n1012), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1035), .A2(new_n1048), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1021), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1023), .B(new_n1052), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1035), .A2(new_n1048), .A3(new_n1012), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1035), .A2(new_n1048), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(new_n1020), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n1001), .A3(new_n1052), .ZN(new_n1058));
  INV_X1    g633(.A(G37), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n969), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1051), .A2(new_n1001), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1057), .A2(new_n1026), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT43), .B1(new_n1067), .B2(KEYINPUT114), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1069), .B(new_n1064), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT44), .B(new_n1063), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1051), .A2(new_n1001), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1057), .A2(new_n1026), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n969), .B(new_n1061), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT44), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1072), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(G397));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  AND3_X1   g657(.A1(G299), .A2(new_n1082), .A3(KEYINPUT57), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(G299), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1384), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n502), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT50), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n465), .A2(new_n470), .A3(G40), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n502), .A2(new_n1090), .A3(new_n1086), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT45), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1086), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1096), .A2(new_n1089), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1085), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  INV_X1    g676(.A(G2067), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n465), .A2(new_n470), .A3(G40), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1087), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1092), .A2(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(new_n640), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1094), .A2(new_n1085), .A3(new_n1099), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1100), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n648), .B1(new_n1105), .B2(KEYINPUT60), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1105), .B2(KEYINPUT60), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1105), .A2(new_n1111), .A3(KEYINPUT60), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1109), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1100), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1107), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1100), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1096), .A2(new_n1089), .A3(new_n1097), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1124), .A2(G1996), .B1(new_n1104), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(KEYINPUT59), .A3(new_n568), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n568), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1120), .A2(new_n1123), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1108), .B1(new_n1118), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  INV_X1    g708(.A(G2084), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1088), .A2(new_n1134), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1135));
  INV_X1    g710(.A(G1966), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1133), .A2(new_n1135), .B1(new_n1124), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(KEYINPUT120), .A3(new_n1134), .A4(new_n1088), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(G168), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(G8), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1135), .A2(new_n1133), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1124), .A2(new_n1136), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1139), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G168), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1137), .A2(G286), .A3(new_n1139), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G8), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1142), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1104), .A2(new_n1150), .ZN(new_n1153));
  INV_X1    g728(.A(G1976), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT52), .B1(G288), .B2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1153), .B(new_n1155), .C1(new_n1154), .C2(G288), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT49), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n599), .A2(new_n602), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n521), .A2(new_n600), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n730), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G305), .A2(G1981), .ZN(new_n1162));
  OAI211_X1 g737(.A(KEYINPUT119), .B(new_n1157), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1162), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n599), .A2(new_n602), .ZN(new_n1165));
  OAI21_X1  g740(.A(G1981), .B1(new_n1165), .B2(new_n1159), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1157), .A2(KEYINPUT119), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1163), .A2(new_n1168), .A3(new_n1153), .ZN(new_n1169));
  OAI221_X1 g744(.A(G8), .B1(G288), .B2(new_n1154), .C1(new_n1087), .C2(new_n1103), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1170), .A2(new_n1171), .A3(KEYINPUT52), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1170), .B2(KEYINPUT52), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1156), .B(new_n1169), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1124), .A2(KEYINPUT117), .ZN(new_n1175));
  INV_X1    g750(.A(G1971), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1096), .A2(new_n1177), .A3(new_n1089), .A4(new_n1097), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1092), .A2(G2090), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1150), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(G303), .A2(G8), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT55), .Z(new_n1183));
  AOI21_X1  g758(.A(new_n1174), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(G8), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AND4_X1   g763(.A1(new_n1143), .A2(new_n1152), .A3(new_n1184), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT54), .ZN(new_n1190));
  INV_X1    g765(.A(G1961), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1092), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT53), .ZN(new_n1193));
  OR3_X1    g768(.A1(new_n1124), .A2(new_n1193), .A3(G2078), .ZN(new_n1194));
  AOI21_X1  g769(.A(G2078), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1192), .B(new_n1194), .C1(new_n1195), .C2(KEYINPUT53), .ZN(new_n1196));
  INV_X1    g771(.A(G301), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n470), .B(KEYINPUT124), .Z(new_n1199));
  INV_X1    g774(.A(G40), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1193), .A2(new_n1200), .A3(G2078), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n465), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1199), .A2(new_n1096), .A3(new_n1097), .A4(new_n1202), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1192), .B(new_n1203), .C1(new_n1195), .C2(KEYINPUT53), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(G171), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1190), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1190), .B1(new_n1204), .B2(new_n1197), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1132), .B(new_n1189), .C1(new_n1206), .C2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1152), .A2(KEYINPUT62), .A3(new_n1143), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(KEYINPUT125), .ZN(new_n1211));
  AND4_X1   g786(.A1(new_n1197), .A2(new_n1184), .A3(new_n1188), .A4(new_n1196), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1152), .A2(new_n1143), .A3(new_n1213), .A4(KEYINPUT62), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n1215));
  AOI211_X1 g790(.A(new_n1142), .B(new_n1150), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT51), .B1(new_n1140), .B2(G8), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1184), .A2(new_n1188), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1221), .A2(KEYINPUT121), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(KEYINPUT121), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1184), .A2(new_n1188), .A3(new_n1224), .A4(new_n1220), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NOR3_X1   g801(.A1(new_n1186), .A2(new_n1174), .A3(new_n1187), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1169), .A2(new_n1154), .A3(new_n764), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1164), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1227), .B1(new_n1153), .B2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g805(.A1(new_n1209), .A2(new_n1219), .A3(new_n1226), .A4(new_n1230), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n777), .A2(new_n750), .ZN(new_n1234));
  AOI21_X1  g809(.A(new_n1233), .B1(new_n1234), .B2(KEYINPUT115), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1235), .B1(KEYINPUT115), .B2(new_n1234), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1232), .A2(G1986), .A3(G290), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT116), .ZN(new_n1239));
  XNOR2_X1  g814(.A(new_n886), .B(G2067), .ZN(new_n1240));
  NOR2_X1   g815(.A1(new_n817), .A2(G1996), .ZN(new_n1241));
  INV_X1    g816(.A(G1996), .ZN(new_n1242));
  NOR3_X1   g817(.A1(new_n810), .A2(new_n816), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1240), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n788), .B(new_n791), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1245), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1232), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  AND2_X1   g822(.A1(new_n1239), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1231), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1233), .B1(new_n1240), .B2(new_n817), .ZN(new_n1250));
  INV_X1    g825(.A(KEYINPUT46), .ZN(new_n1251));
  NOR3_X1   g826(.A1(new_n1233), .A2(new_n1251), .A3(G1996), .ZN(new_n1252));
  AOI21_X1  g827(.A(KEYINPUT46), .B1(new_n1232), .B2(new_n1242), .ZN(new_n1253));
  OR3_X1    g828(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g829(.A(KEYINPUT47), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n886), .A2(new_n1102), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n789), .A2(new_n791), .ZN(new_n1257));
  OAI21_X1  g832(.A(new_n1256), .B1(new_n1244), .B2(new_n1257), .ZN(new_n1258));
  AOI22_X1  g833(.A1(new_n1254), .A2(new_n1255), .B1(new_n1232), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g834(.A(KEYINPUT48), .ZN(new_n1260));
  NOR2_X1   g835(.A1(new_n1236), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1236), .A2(new_n1260), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1262), .A2(new_n1247), .ZN(new_n1263));
  OAI221_X1 g838(.A(new_n1259), .B1(new_n1255), .B2(new_n1254), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g839(.A(new_n1264), .B(KEYINPUT126), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1249), .A2(new_n1265), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g841(.A1(new_n725), .A2(new_n727), .A3(G319), .ZN(new_n1268));
  AOI21_X1  g842(.A(new_n1268), .B1(new_n757), .B2(new_n760), .ZN(new_n1269));
  NAND2_X1  g843(.A1(new_n708), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g844(.A(new_n1270), .B1(new_n972), .B2(new_n976), .ZN(new_n1271));
  AND3_X1   g845(.A1(new_n1077), .A2(new_n1271), .A3(KEYINPUT127), .ZN(new_n1272));
  AOI21_X1  g846(.A(KEYINPUT127), .B1(new_n1077), .B2(new_n1271), .ZN(new_n1273));
  NOR2_X1   g847(.A1(new_n1272), .A2(new_n1273), .ZN(G308));
  NAND2_X1  g848(.A1(new_n1077), .A2(new_n1271), .ZN(G225));
endmodule


