

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744;

  XNOR2_X1 U374 ( .A(n471), .B(KEYINPUT4), .ZN(n485) );
  INV_X1 U375 ( .A(KEYINPUT16), .ZN(n358) );
  INV_X2 U376 ( .A(G953), .ZN(n735) );
  XOR2_X2 U377 ( .A(KEYINPUT31), .B(n526), .Z(n711) );
  NAND2_X2 U378 ( .A1(n352), .A2(n408), .ZN(n515) );
  INV_X2 U379 ( .A(n659), .ZN(n372) );
  OR2_X2 U380 ( .A1(n363), .A2(G902), .ZN(n503) );
  INV_X1 U381 ( .A(G140), .ZN(n498) );
  NOR2_X2 U382 ( .A1(n617), .A2(n647), .ZN(n619) );
  XNOR2_X2 U383 ( .A(n430), .B(KEYINPUT33), .ZN(n683) );
  XNOR2_X2 U384 ( .A(n385), .B(KEYINPUT1), .ZN(n554) );
  INV_X1 U385 ( .A(n658), .ZN(n353) );
  INV_X2 U386 ( .A(G125), .ZN(n401) );
  NOR2_X1 U387 ( .A1(n634), .A2(n647), .ZN(n635) );
  NOR2_X1 U388 ( .A1(n623), .A2(n647), .ZN(n624) );
  AND2_X2 U389 ( .A1(n613), .A2(n612), .ZN(n373) );
  AND2_X1 U390 ( .A1(n357), .A2(n584), .ZN(n356) );
  OR2_X1 U391 ( .A1(n682), .A2(n589), .ZN(n361) );
  XNOR2_X1 U392 ( .A(n376), .B(KEYINPUT22), .ZN(n521) );
  NAND2_X1 U393 ( .A1(n379), .A2(n599), .ZN(n734) );
  XNOR2_X1 U394 ( .A(n359), .B(n591), .ZN(n379) );
  NAND2_X1 U395 ( .A1(n356), .A2(n360), .ZN(n359) );
  AND2_X1 U396 ( .A1(n583), .A2(n582), .ZN(n357) );
  XNOR2_X1 U397 ( .A(n590), .B(n371), .ZN(n360) );
  XNOR2_X1 U398 ( .A(n588), .B(n587), .ZN(n636) );
  XNOR2_X1 U399 ( .A(n354), .B(KEYINPUT47), .ZN(n563) );
  XNOR2_X1 U400 ( .A(n361), .B(KEYINPUT42), .ZN(n744) );
  XNOR2_X1 U401 ( .A(n355), .B(KEYINPUT76), .ZN(n704) );
  NOR2_X1 U402 ( .A1(n589), .A2(n560), .ZN(n355) );
  XNOR2_X1 U403 ( .A(n362), .B(KEYINPUT41), .ZN(n682) );
  INV_X1 U404 ( .A(n521), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n572), .B(KEYINPUT75), .ZN(n411) );
  NOR2_X1 U406 ( .A1(n671), .A2(n670), .ZN(n362) );
  NAND2_X1 U407 ( .A1(n437), .A2(n571), .ZN(n572) );
  XNOR2_X1 U408 ( .A(n529), .B(n528), .ZN(n707) );
  XNOR2_X1 U409 ( .A(n519), .B(KEYINPUT6), .ZN(n409) );
  XNOR2_X1 U410 ( .A(n494), .B(n493), .ZN(n519) );
  XNOR2_X1 U411 ( .A(n377), .B(n364), .ZN(n363) );
  XNOR2_X1 U412 ( .A(n498), .B(KEYINPUT10), .ZN(n429) );
  XNOR2_X1 U413 ( .A(n358), .B(G110), .ZN(n393) );
  XNOR2_X1 U414 ( .A(KEYINPUT15), .B(G902), .ZN(n606) );
  NAND2_X1 U415 ( .A1(n704), .A2(n561), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n363), .B(n644), .ZN(n645) );
  NOR2_X1 U417 ( .A1(n629), .A2(n647), .ZN(n630) );
  NOR2_X2 U418 ( .A1(n525), .A2(n663), .ZN(n526) );
  XNOR2_X2 U419 ( .A(n721), .B(n496), .ZN(n492) );
  INV_X1 U420 ( .A(n507), .ZN(n378) );
  NOR2_X1 U421 ( .A1(n530), .A2(n527), .ZN(n580) );
  NOR2_X1 U422 ( .A1(n397), .A2(n547), .ZN(n570) );
  XNOR2_X1 U423 ( .A(n546), .B(KEYINPUT101), .ZN(n397) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n488) );
  INV_X1 U425 ( .A(G134), .ZN(n483) );
  XNOR2_X1 U426 ( .A(KEYINPUT69), .B(G137), .ZN(n507) );
  INV_X1 U427 ( .A(KEYINPUT45), .ZN(n541) );
  XNOR2_X1 U428 ( .A(n419), .B(n417), .ZN(n504) );
  XNOR2_X1 U429 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n419) );
  NOR2_X1 U430 ( .A1(n418), .A2(G953), .ZN(n417) );
  INV_X1 U431 ( .A(G234), .ZN(n418) );
  XNOR2_X1 U432 ( .A(n507), .B(n505), .ZN(n416) );
  XNOR2_X1 U433 ( .A(G128), .B(KEYINPUT79), .ZN(n505) );
  XNOR2_X1 U434 ( .A(n506), .B(n508), .ZN(n414) );
  XNOR2_X1 U435 ( .A(KEYINPUT66), .B(G101), .ZN(n496) );
  NAND2_X1 U436 ( .A1(n550), .A2(n405), .ZN(n551) );
  AND2_X1 U437 ( .A1(n707), .A2(n557), .ZN(n550) );
  XNOR2_X1 U438 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U439 ( .A(KEYINPUT34), .ZN(n403) );
  OR2_X1 U440 ( .A1(n670), .A2(n548), .ZN(n461) );
  XNOR2_X1 U441 ( .A(n559), .B(n558), .ZN(n394) );
  XNOR2_X1 U442 ( .A(n444), .B(n422), .ZN(n530) );
  XNOR2_X1 U443 ( .A(n445), .B(G475), .ZN(n422) );
  XNOR2_X1 U444 ( .A(n455), .B(n421), .ZN(n527) );
  XNOR2_X1 U445 ( .A(n456), .B(n457), .ZN(n421) );
  XNOR2_X1 U446 ( .A(n427), .B(n423), .ZN(n631) );
  XNOR2_X1 U447 ( .A(n426), .B(n424), .ZN(n423) );
  XNOR2_X1 U448 ( .A(n733), .B(n428), .ZN(n427) );
  XNOR2_X1 U449 ( .A(n442), .B(n425), .ZN(n424) );
  NOR2_X1 U450 ( .A1(n735), .A2(G952), .ZN(n647) );
  NAND2_X1 U451 ( .A1(n598), .A2(n707), .ZN(n588) );
  OR2_X1 U452 ( .A1(G237), .A2(G902), .ZN(n476) );
  INV_X1 U453 ( .A(KEYINPUT104), .ZN(n432) );
  INV_X1 U454 ( .A(G902), .ZN(n509) );
  XNOR2_X1 U455 ( .A(G146), .B(G116), .ZN(n486) );
  XOR2_X1 U456 ( .A(KEYINPUT5), .B(G137), .Z(n487) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n477) );
  NAND2_X1 U458 ( .A1(G237), .A2(G234), .ZN(n398) );
  XNOR2_X1 U459 ( .A(KEYINPUT72), .B(KEYINPUT14), .ZN(n399) );
  NOR2_X1 U460 ( .A1(n658), .A2(n409), .ZN(n431) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n549) );
  INV_X1 U462 ( .A(KEYINPUT70), .ZN(n395) );
  NOR2_X1 U463 ( .A1(n570), .A2(n548), .ZN(n396) );
  NAND2_X1 U464 ( .A1(n380), .A2(n653), .ZN(n658) );
  XNOR2_X1 U465 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n447) );
  XNOR2_X1 U466 ( .A(G134), .B(G122), .ZN(n449) );
  XOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n450) );
  XNOR2_X1 U468 ( .A(n446), .B(G107), .ZN(n462) );
  INV_X1 U469 ( .A(G116), .ZN(n446) );
  XNOR2_X1 U470 ( .A(G113), .B(G143), .ZN(n442) );
  INV_X1 U471 ( .A(KEYINPUT92), .ZN(n425) );
  XNOR2_X1 U472 ( .A(n443), .B(n441), .ZN(n428) );
  XNOR2_X1 U473 ( .A(n463), .B(n440), .ZN(n426) );
  XNOR2_X1 U474 ( .A(KEYINPUT86), .B(KEYINPUT18), .ZN(n466) );
  XOR2_X1 U475 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n467) );
  XNOR2_X1 U476 ( .A(n407), .B(n406), .ZN(n719) );
  INV_X1 U477 ( .A(n462), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n393), .B(n439), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n412), .B(KEYINPUT39), .ZN(n598) );
  NAND2_X1 U480 ( .A1(n352), .A2(n367), .ZN(n388) );
  INV_X1 U481 ( .A(KEYINPUT3), .ZN(n464) );
  XNOR2_X1 U482 ( .A(n415), .B(n413), .ZN(n637) );
  XNOR2_X1 U483 ( .A(n434), .B(n414), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n733), .B(n416), .ZN(n415) );
  NAND2_X1 U485 ( .A1(n402), .A2(n580), .ZN(n518) );
  AND2_X1 U486 ( .A1(n514), .A2(n409), .ZN(n408) );
  INV_X1 U487 ( .A(n527), .ZN(n531) );
  INV_X1 U488 ( .A(n388), .ZN(n699) );
  NAND2_X1 U489 ( .A1(n527), .A2(n420), .ZN(n529) );
  INV_X1 U490 ( .A(n530), .ZN(n420) );
  XNOR2_X1 U491 ( .A(n524), .B(n387), .ZN(n534) );
  INV_X1 U492 ( .A(KEYINPUT100), .ZN(n387) );
  XOR2_X1 U493 ( .A(KEYINPUT121), .B(n620), .Z(n621) );
  XOR2_X1 U494 ( .A(KEYINPUT59), .B(n631), .Z(n632) );
  XNOR2_X1 U495 ( .A(n534), .B(n386), .ZN(G3) );
  INV_X1 U496 ( .A(G101), .ZN(n386) );
  XOR2_X1 U497 ( .A(n502), .B(n501), .Z(n364) );
  XNOR2_X1 U498 ( .A(n512), .B(n511), .ZN(n365) );
  OR2_X1 U499 ( .A1(n433), .A2(n656), .ZN(n366) );
  AND2_X1 U500 ( .A1(n659), .A2(n520), .ZN(n367) );
  AND2_X1 U501 ( .A1(n575), .A2(n668), .ZN(n368) );
  AND2_X1 U502 ( .A1(n353), .A2(n656), .ZN(n369) );
  XNOR2_X1 U503 ( .A(KEYINPUT65), .B(KEYINPUT0), .ZN(n370) );
  XOR2_X1 U504 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n371) );
  XNOR2_X1 U505 ( .A(n433), .B(n432), .ZN(n437) );
  AND2_X1 U506 ( .A1(n613), .A2(n612), .ZN(n641) );
  INV_X1 U507 ( .A(n373), .ZN(n374) );
  INV_X1 U508 ( .A(n374), .ZN(n375) );
  XNOR2_X1 U509 ( .A(n491), .B(n492), .ZN(n382) );
  XNOR2_X1 U510 ( .A(n719), .B(n492), .ZN(n392) );
  NAND2_X1 U511 ( .A1(n372), .A2(n369), .ZN(n663) );
  NAND2_X1 U512 ( .A1(n683), .A2(n381), .ZN(n404) );
  NAND2_X1 U513 ( .A1(n482), .A2(n381), .ZN(n376) );
  XNOR2_X2 U514 ( .A(n384), .B(n378), .ZN(n377) );
  XNOR2_X1 U515 ( .A(n377), .B(n733), .ZN(n737) );
  INV_X1 U516 ( .A(n380), .ZN(n522) );
  XNOR2_X2 U517 ( .A(n513), .B(n365), .ZN(n380) );
  AND2_X1 U518 ( .A1(n522), .A2(n548), .ZN(n654) );
  NOR2_X1 U519 ( .A1(n549), .A2(n380), .ZN(n557) );
  NOR2_X1 U520 ( .A1(n656), .A2(n380), .ZN(n520) );
  NOR2_X1 U521 ( .A1(n659), .A2(n380), .ZN(n514) );
  XNOR2_X2 U522 ( .A(n481), .B(n370), .ZN(n381) );
  INV_X1 U523 ( .A(n381), .ZN(n525) );
  NOR2_X1 U524 ( .A1(n525), .A2(n366), .ZN(n694) );
  XNOR2_X1 U525 ( .A(n384), .B(n382), .ZN(n614) );
  XNOR2_X2 U526 ( .A(n485), .B(n484), .ZN(n384) );
  AND2_X2 U527 ( .A1(n383), .A2(n388), .ZN(n390) );
  AND2_X1 U528 ( .A1(n383), .A2(n742), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n383), .B(G122), .ZN(G24) );
  XNOR2_X2 U530 ( .A(n518), .B(n517), .ZN(n383) );
  NAND2_X1 U531 ( .A1(n353), .A2(n385), .ZN(n433) );
  NAND2_X1 U532 ( .A1(n394), .A2(n385), .ZN(n589) );
  XNOR2_X2 U533 ( .A(n503), .B(G469), .ZN(n385) );
  NAND2_X1 U534 ( .A1(n389), .A2(KEYINPUT44), .ZN(n536) );
  NAND2_X1 U535 ( .A1(n390), .A2(n742), .ZN(n389) );
  XNOR2_X2 U536 ( .A(n515), .B(KEYINPUT32), .ZN(n742) );
  XNOR2_X1 U537 ( .A(n392), .B(n473), .ZN(n626) );
  BUF_X1 U538 ( .A(n683), .Z(n391) );
  XNOR2_X1 U539 ( .A(n400), .B(n470), .ZN(n472) );
  NAND2_X1 U540 ( .A1(n556), .A2(n480), .ZN(n481) );
  XNOR2_X2 U541 ( .A(n552), .B(KEYINPUT19), .ZN(n556) );
  XNOR2_X1 U542 ( .A(n468), .B(n469), .ZN(n400) );
  XNOR2_X2 U543 ( .A(n401), .B(G146), .ZN(n468) );
  INV_X1 U544 ( .A(n554), .ZN(n659) );
  NOR2_X1 U545 ( .A1(n521), .A2(n405), .ZN(n410) );
  INV_X1 U546 ( .A(n409), .ZN(n405) );
  INV_X1 U547 ( .A(n439), .ZN(n463) );
  NAND2_X1 U548 ( .A1(n410), .A2(n523), .ZN(n524) );
  AND2_X1 U549 ( .A1(n411), .A2(n575), .ZN(n586) );
  NAND2_X1 U550 ( .A1(n411), .A2(n368), .ZN(n412) );
  NAND2_X1 U551 ( .A1(n431), .A2(n554), .ZN(n430) );
  NAND2_X1 U552 ( .A1(n527), .A2(n530), .ZN(n670) );
  XNOR2_X2 U553 ( .A(n468), .B(n429), .ZN(n733) );
  NAND2_X1 U554 ( .A1(n504), .A2(G221), .ZN(n434) );
  XNOR2_X1 U555 ( .A(n542), .B(n541), .ZN(n608) );
  XNOR2_X1 U556 ( .A(n734), .B(n600), .ZN(n601) );
  XOR2_X1 U557 ( .A(KEYINPUT36), .B(KEYINPUT109), .Z(n435) );
  OR2_X1 U558 ( .A1(n606), .A2(n605), .ZN(n436) );
  INV_X1 U559 ( .A(KEYINPUT73), .ZN(n600) );
  INV_X1 U560 ( .A(KEYINPUT80), .ZN(n603) );
  XNOR2_X1 U561 ( .A(KEYINPUT93), .B(KEYINPUT13), .ZN(n445) );
  XNOR2_X2 U562 ( .A(G122), .B(G104), .ZN(n439) );
  XOR2_X1 U563 ( .A(KEYINPUT11), .B(KEYINPUT91), .Z(n441) );
  NAND2_X1 U564 ( .A1(G214), .A2(n488), .ZN(n440) );
  XOR2_X1 U565 ( .A(KEYINPUT12), .B(G131), .Z(n443) );
  NOR2_X1 U566 ( .A1(G902), .A2(n631), .ZN(n444) );
  XNOR2_X1 U567 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n456) );
  XNOR2_X2 U568 ( .A(G143), .B(G128), .ZN(n471) );
  XOR2_X1 U569 ( .A(n471), .B(n447), .Z(n448) );
  XNOR2_X1 U570 ( .A(n462), .B(n448), .ZN(n454) );
  NAND2_X1 U571 ( .A1(G217), .A2(n504), .ZN(n452) );
  XNOR2_X1 U572 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U573 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U574 ( .A(n454), .B(n453), .ZN(n620) );
  NOR2_X1 U575 ( .A1(G902), .A2(n620), .ZN(n455) );
  INV_X1 U576 ( .A(G478), .ZN(n457) );
  NAND2_X1 U577 ( .A1(n606), .A2(G234), .ZN(n458) );
  XNOR2_X1 U578 ( .A(n458), .B(KEYINPUT20), .ZN(n510) );
  NAND2_X1 U579 ( .A1(n510), .A2(G221), .ZN(n460) );
  INV_X1 U580 ( .A(KEYINPUT21), .ZN(n459) );
  XNOR2_X1 U581 ( .A(n460), .B(n459), .ZN(n653) );
  INV_X1 U582 ( .A(n653), .ZN(n548) );
  XNOR2_X1 U583 ( .A(n461), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X2 U584 ( .A(G119), .B(G113), .ZN(n465) );
  XNOR2_X2 U585 ( .A(n465), .B(n464), .ZN(n721) );
  XNOR2_X1 U586 ( .A(n467), .B(n466), .ZN(n470) );
  NAND2_X1 U587 ( .A1(G224), .A2(n735), .ZN(n469) );
  XNOR2_X1 U588 ( .A(n485), .B(n472), .ZN(n473) );
  NAND2_X1 U589 ( .A1(n626), .A2(n606), .ZN(n475) );
  AND2_X1 U590 ( .A1(G210), .A2(n476), .ZN(n474) );
  XNOR2_X2 U591 ( .A(n475), .B(n474), .ZN(n576) );
  NAND2_X1 U592 ( .A1(G214), .A2(n476), .ZN(n667) );
  NAND2_X2 U593 ( .A1(n576), .A2(n667), .ZN(n552) );
  AND2_X1 U594 ( .A1(n477), .A2(G952), .ZN(n680) );
  AND2_X1 U595 ( .A1(n680), .A2(n735), .ZN(n547) );
  XOR2_X1 U596 ( .A(G898), .B(KEYINPUT88), .Z(n728) );
  NAND2_X1 U597 ( .A1(G953), .A2(n728), .ZN(n723) );
  NAND2_X1 U598 ( .A1(G902), .A2(n477), .ZN(n544) );
  NOR2_X1 U599 ( .A1(n723), .A2(n544), .ZN(n478) );
  NOR2_X1 U600 ( .A1(n547), .A2(n478), .ZN(n479) );
  XNOR2_X1 U601 ( .A(KEYINPUT89), .B(n479), .ZN(n480) );
  XNOR2_X1 U602 ( .A(n483), .B(G131), .ZN(n484) );
  XNOR2_X1 U603 ( .A(n487), .B(n486), .ZN(n490) );
  NAND2_X1 U604 ( .A1(n488), .A2(G210), .ZN(n489) );
  XNOR2_X1 U605 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U606 ( .A1(n614), .A2(n509), .ZN(n494) );
  XOR2_X1 U607 ( .A(G472), .B(KEYINPUT71), .Z(n493) );
  NAND2_X1 U608 ( .A1(n735), .A2(G227), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n495), .B(G146), .ZN(n497) );
  XNOR2_X1 U610 ( .A(n497), .B(n496), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n498), .B(G107), .ZN(n500) );
  XNOR2_X1 U612 ( .A(G104), .B(G110), .ZN(n499) );
  XNOR2_X1 U613 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U614 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n506) );
  XNOR2_X1 U615 ( .A(G119), .B(G110), .ZN(n508) );
  NAND2_X1 U616 ( .A1(n637), .A2(n509), .ZN(n513) );
  XOR2_X1 U617 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n512) );
  NAND2_X1 U618 ( .A1(n510), .A2(G217), .ZN(n511) );
  INV_X1 U619 ( .A(KEYINPUT82), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n516), .B(KEYINPUT35), .ZN(n517) );
  BUF_X2 U621 ( .A(n519), .Z(n656) );
  NOR2_X1 U622 ( .A1(n372), .A2(n522), .ZN(n523) );
  NOR2_X1 U623 ( .A1(n711), .A2(n694), .ZN(n532) );
  INV_X1 U624 ( .A(KEYINPUT98), .ZN(n528) );
  AND2_X1 U625 ( .A1(n531), .A2(n530), .ZN(n710) );
  OR2_X1 U626 ( .A1(n707), .A2(n710), .ZN(n565) );
  INV_X1 U627 ( .A(n565), .ZN(n672) );
  NOR2_X1 U628 ( .A1(n532), .A2(n672), .ZN(n533) );
  NOR2_X1 U629 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U631 ( .A(n537), .B(KEYINPUT85), .ZN(n540) );
  NOR2_X1 U632 ( .A1(n699), .A2(KEYINPUT44), .ZN(n538) );
  NAND2_X1 U633 ( .A1(n438), .A2(n538), .ZN(n539) );
  NAND2_X1 U634 ( .A1(n540), .A2(n539), .ZN(n542) );
  NOR2_X1 U635 ( .A1(n608), .A2(n606), .ZN(n543) );
  XNOR2_X1 U636 ( .A(n543), .B(KEYINPUT81), .ZN(n602) );
  NOR2_X1 U637 ( .A1(G900), .A2(n544), .ZN(n545) );
  NAND2_X1 U638 ( .A1(G953), .A2(n545), .ZN(n546) );
  XNOR2_X1 U639 ( .A(n551), .B(KEYINPUT102), .ZN(n593) );
  NOR2_X1 U640 ( .A1(n593), .A2(n552), .ZN(n553) );
  XNOR2_X1 U641 ( .A(n553), .B(n435), .ZN(n555) );
  NAND2_X1 U642 ( .A1(n555), .A2(n372), .ZN(n713) );
  XNOR2_X1 U643 ( .A(n713), .B(KEYINPUT84), .ZN(n584) );
  NOR2_X1 U644 ( .A1(n672), .A2(KEYINPUT67), .ZN(n561) );
  INV_X1 U645 ( .A(n556), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n557), .A2(n656), .ZN(n559) );
  XNOR2_X1 U647 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n558) );
  INV_X1 U648 ( .A(KEYINPUT77), .ZN(n562) );
  NAND2_X1 U649 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U650 ( .A1(KEYINPUT47), .A2(n704), .ZN(n564) );
  NAND2_X1 U651 ( .A1(n564), .A2(KEYINPUT77), .ZN(n567) );
  NAND2_X1 U652 ( .A1(n565), .A2(KEYINPUT77), .ZN(n566) );
  AND2_X1 U653 ( .A1(n567), .A2(n566), .ZN(n568) );
  AND2_X1 U654 ( .A1(n569), .A2(n568), .ZN(n583) );
  INV_X1 U655 ( .A(n570), .ZN(n571) );
  NAND2_X1 U656 ( .A1(n656), .A2(n667), .ZN(n574) );
  XNOR2_X1 U657 ( .A(KEYINPUT105), .B(KEYINPUT30), .ZN(n573) );
  XNOR2_X1 U658 ( .A(n574), .B(n573), .ZN(n575) );
  BUF_X1 U659 ( .A(n576), .Z(n577) );
  NAND2_X1 U660 ( .A1(n586), .A2(n577), .ZN(n579) );
  INV_X1 U661 ( .A(KEYINPUT106), .ZN(n578) );
  XNOR2_X1 U662 ( .A(n579), .B(n578), .ZN(n581) );
  NAND2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n702) );
  XNOR2_X1 U664 ( .A(n702), .B(KEYINPUT78), .ZN(n582) );
  XNOR2_X1 U665 ( .A(n577), .B(KEYINPUT38), .ZN(n585) );
  INV_X1 U666 ( .A(n585), .ZN(n668) );
  XNOR2_X1 U667 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n668), .A2(n667), .ZN(n671) );
  NAND2_X1 U669 ( .A1(n636), .A2(n744), .ZN(n590) );
  XNOR2_X1 U670 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n659), .A2(n667), .ZN(n592) );
  NOR2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U673 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n594) );
  XNOR2_X1 U674 ( .A(n595), .B(n594), .ZN(n597) );
  INV_X1 U675 ( .A(n577), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n718) );
  NAND2_X1 U677 ( .A1(n598), .A2(n710), .ZN(n716) );
  AND2_X1 U678 ( .A1(n718), .A2(n716), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n604), .B(n603), .ZN(n607) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n607), .A2(n436), .ZN(n613) );
  BUF_X1 U683 ( .A(n608), .Z(n649) );
  INV_X1 U684 ( .A(n734), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n609), .A2(KEYINPUT2), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n649), .A2(n610), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT74), .ZN(n652) );
  INV_X1 U688 ( .A(n652), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n641), .A2(G472), .ZN(n616) );
  XOR2_X1 U690 ( .A(KEYINPUT62), .B(n614), .Z(n615) );
  XNOR2_X1 U691 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U692 ( .A(KEYINPUT63), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(G57) );
  NAND2_X1 U694 ( .A1(n373), .A2(G478), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U697 ( .A1(n641), .A2(G210), .ZN(n628) );
  XNOR2_X1 U698 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U702 ( .A1(n373), .A2(G475), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U705 ( .A(n636), .B(G131), .ZN(G33) );
  NAND2_X1 U706 ( .A1(n375), .A2(G217), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT123), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U709 ( .A1(n640), .A2(n647), .ZN(G66) );
  NAND2_X1 U710 ( .A1(n375), .A2(G469), .ZN(n646) );
  XNOR2_X1 U711 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n643) );
  XNOR2_X1 U712 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(n648) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(G54) );
  NOR2_X1 U716 ( .A1(n649), .A2(n734), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n690) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(n654), .Z(n655) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U721 ( .A(KEYINPUT117), .B(n657), .Z(n662) );
  NAND2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT50), .ZN(n661) );
  NAND2_X1 U724 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U726 ( .A(KEYINPUT51), .B(n665), .ZN(n666) );
  NOR2_X1 U727 ( .A1(n682), .A2(n666), .ZN(n678) );
  NOR2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U731 ( .A1(n674), .A2(n673), .ZN(n676) );
  INV_X1 U732 ( .A(n391), .ZN(n675) );
  NOR2_X1 U733 ( .A1(n676), .A2(n675), .ZN(n677) );
  OR2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n679), .B(KEYINPUT52), .ZN(n681) );
  NAND2_X1 U736 ( .A1(n681), .A2(n680), .ZN(n688) );
  INV_X1 U737 ( .A(n682), .ZN(n684) );
  NAND2_X1 U738 ( .A1(n684), .A2(n391), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n685), .B(KEYINPUT118), .ZN(n686) );
  AND2_X1 U740 ( .A1(n686), .A2(n735), .ZN(n687) );
  NAND2_X1 U741 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U742 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n691), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U744 ( .A1(n707), .A2(n694), .ZN(n692) );
  XNOR2_X1 U745 ( .A(n692), .B(KEYINPUT110), .ZN(n693) );
  XNOR2_X1 U746 ( .A(G104), .B(n693), .ZN(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT26), .B(KEYINPUT111), .Z(n696) );
  NAND2_X1 U748 ( .A1(n694), .A2(n710), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n696), .B(n695), .ZN(n698) );
  XOR2_X1 U750 ( .A(G107), .B(KEYINPUT27), .Z(n697) );
  XNOR2_X1 U751 ( .A(n698), .B(n697), .ZN(G9) );
  XOR2_X1 U752 ( .A(G110), .B(n699), .Z(G12) );
  XOR2_X1 U753 ( .A(G128), .B(KEYINPUT29), .Z(n701) );
  NAND2_X1 U754 ( .A1(n710), .A2(n704), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(G30) );
  XNOR2_X1 U756 ( .A(G143), .B(KEYINPUT112), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(G45) );
  XOR2_X1 U758 ( .A(G146), .B(KEYINPUT113), .Z(n706) );
  NAND2_X1 U759 ( .A1(n704), .A2(n707), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(G48) );
  NAND2_X1 U761 ( .A1(n707), .A2(n711), .ZN(n708) );
  XNOR2_X1 U762 ( .A(n708), .B(KEYINPUT114), .ZN(n709) );
  XNOR2_X1 U763 ( .A(G113), .B(n709), .ZN(G15) );
  NAND2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n712), .B(G116), .ZN(G18) );
  XOR2_X1 U766 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n715) );
  XOR2_X1 U767 ( .A(n713), .B(G125), .Z(n714) );
  XNOR2_X1 U768 ( .A(n715), .B(n714), .ZN(G27) );
  XNOR2_X1 U769 ( .A(n716), .B(G134), .ZN(n717) );
  XNOR2_X1 U770 ( .A(KEYINPUT116), .B(n717), .ZN(G36) );
  XNOR2_X1 U771 ( .A(G140), .B(n718), .ZN(G42) );
  XOR2_X1 U772 ( .A(n719), .B(G101), .Z(n720) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n732) );
  NOR2_X1 U775 ( .A1(n649), .A2(G953), .ZN(n724) );
  XOR2_X1 U776 ( .A(KEYINPUT125), .B(n724), .Z(n730) );
  XOR2_X1 U777 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n726) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(G69) );
  XNOR2_X1 U783 ( .A(n734), .B(n737), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n737), .B(G227), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U789 ( .A(n742), .B(G119), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U791 ( .A(G137), .B(n744), .ZN(G39) );
endmodule

