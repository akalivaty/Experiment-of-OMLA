//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n203), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g0010(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n203), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NOR2_X1   g0014(.A1(G58), .A2(G68), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n216), .A2(G50), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n211), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n210), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  INV_X1    g0031(.A(G50), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(G68), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G116), .Z(new_n240));
  INV_X1    g0040(.A(G107), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G97), .ZN(new_n242));
  INV_X1    g0042(.A(G97), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G107), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n217), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n248), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G50), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(new_n232), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n218), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n218), .B1(new_n215), .B2(new_n232), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n252), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G222), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n271), .B1(new_n272), .B2(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n282), .A3(G274), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n276), .A2(new_n280), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(G226), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n268), .B1(new_n288), .B2(G169), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n289), .A2(KEYINPUT67), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(KEYINPUT67), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n259), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n287), .A2(G200), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT74), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n268), .A2(new_n300), .B1(new_n288), .B2(G190), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n297), .A2(new_n299), .A3(new_n304), .A4(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n308), .A2(new_n310), .A3(G226), .A4(G1698), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(G223), .A4(new_n270), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G87), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n276), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(G232), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n283), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n291), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n276), .B2(new_n314), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(G169), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n308), .A2(new_n310), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT7), .B1(new_n323), .B2(new_n218), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  AOI211_X1 g0125(.A(new_n325), .B(G20), .C1(new_n308), .C2(new_n310), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n234), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n215), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n263), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n325), .B1(new_n269), .B2(G20), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n323), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n234), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n338), .B2(new_n332), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n339), .A3(new_n252), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n260), .B1(new_n248), .B2(G20), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n253), .B1(new_n260), .B2(new_n250), .ZN(new_n342));
  AOI211_X1 g0142(.A(KEYINPUT18), .B(new_n322), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(new_n322), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT75), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n342), .ZN(new_n349));
  INV_X1    g0149(.A(new_n252), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n327), .A2(new_n333), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n335), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(new_n334), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT18), .B1(new_n353), .B2(new_n322), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n345), .A2(new_n346), .A3(new_n344), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n315), .A2(new_n358), .A3(new_n319), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G200), .B2(new_n321), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n340), .A2(new_n342), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n340), .A2(new_n360), .A3(KEYINPUT17), .A4(new_n342), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n348), .A2(new_n357), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n269), .A2(G226), .A3(new_n270), .ZN(new_n370));
  INV_X1    g0170(.A(G232), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n370), .B1(new_n307), .B2(new_n243), .C1(new_n273), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n276), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n284), .B1(G238), .B2(new_n285), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n369), .A3(new_n374), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G200), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n250), .A2(new_n234), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT12), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n234), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n272), .B2(new_n261), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n253), .A2(G68), .A3(new_n254), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT11), .B1(new_n383), .B2(new_n252), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n376), .A2(G190), .A3(new_n377), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n379), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n378), .A2(G169), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT14), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n378), .A2(new_n394), .A3(G169), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n395), .C1(new_n291), .C2(new_n378), .ZN(new_n396));
  INV_X1    g0196(.A(new_n388), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n253), .A2(G77), .A3(new_n254), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n249), .A2(G77), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n260), .A2(new_n264), .B1(new_n218), .B2(new_n272), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT70), .ZN(new_n406));
  INV_X1    g0206(.A(new_n261), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n401), .B(new_n403), .C1(new_n350), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n408), .A2(new_n350), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(KEYINPUT72), .A3(new_n401), .A4(new_n403), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n285), .A2(G244), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n283), .ZN(new_n416));
  INV_X1    g0216(.A(new_n273), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(G238), .B1(G107), .B2(new_n323), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n269), .A2(G232), .A3(new_n270), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT68), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT68), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n269), .A2(new_n421), .A3(G232), .A4(new_n270), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n282), .B1(new_n424), .B2(KEYINPUT69), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT69), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n418), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n416), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n411), .B(new_n413), .C1(new_n414), .C2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n428), .A2(G190), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n409), .B1(new_n428), .B2(G169), .ZN(new_n432));
  AOI211_X1 g0232(.A(G179), .B(new_n416), .C1(new_n425), .C2(new_n427), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n306), .A2(new_n368), .A3(new_n398), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n438));
  NAND2_X1  g0238(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n242), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n440), .A2(KEYINPUT77), .B1(new_n245), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(KEYINPUT77), .A3(G97), .A4(new_n241), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT78), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(G97), .A3(new_n241), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT77), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT78), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n245), .A2(new_n441), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n443), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n445), .A2(G20), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n241), .B1(new_n336), .B2(new_n337), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(G77), .B2(new_n263), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n252), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n250), .A2(new_n243), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n248), .A2(G33), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n350), .A2(new_n249), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(new_n243), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n279), .A2(G1), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G257), .A3(new_n282), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  AND2_X1   g0268(.A1(G1), .A2(G13), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n281), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n467), .A2(KEYINPUT80), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT80), .B1(new_n467), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n308), .A2(new_n310), .A3(G244), .A4(new_n270), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n477), .A2(G1698), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(new_n308), .A3(new_n310), .A4(G244), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n269), .A2(KEYINPUT79), .A3(G244), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n276), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n475), .A2(new_n291), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n475), .A2(KEYINPUT81), .A3(new_n291), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n475), .A2(new_n488), .ZN(new_n494));
  INV_X1    g0294(.A(G169), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n462), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT85), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n494), .A2(G190), .ZN(new_n499));
  AOI21_X1  g0299(.A(G200), .B1(new_n475), .B2(new_n488), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n456), .B(new_n461), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n308), .A2(new_n310), .A3(G244), .A4(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n308), .A2(new_n310), .A3(G238), .A4(new_n270), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n503), .C1(new_n307), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n276), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n248), .A2(G45), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G250), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT82), .B1(new_n276), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n282), .A2(new_n510), .A3(G250), .A4(new_n507), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n509), .A2(new_n511), .B1(new_n470), .B2(new_n463), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n506), .A2(new_n512), .A3(G190), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n269), .A2(new_n218), .A3(G68), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n261), .B2(new_n243), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT83), .B(G87), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n520), .A2(new_n521), .B1(new_n218), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n252), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT70), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n405), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n250), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n253), .A2(G87), .A3(new_n458), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n506), .A2(new_n512), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n506), .A2(new_n512), .A3(KEYINPUT84), .A4(G190), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n515), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n495), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n524), .B(new_n527), .C1(new_n526), .C2(new_n459), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n506), .A2(new_n512), .A3(new_n291), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n497), .A2(new_n498), .A3(new_n501), .A4(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n491), .A2(new_n492), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n350), .B1(new_n452), .B2(new_n454), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n496), .B1(new_n541), .B2(new_n460), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n501), .B(new_n538), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT85), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT87), .B1(new_n250), .B2(new_n504), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT87), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n249), .A2(new_n546), .A3(G116), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n459), .A2(new_n504), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n251), .A2(new_n217), .B1(G20), .B2(new_n504), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n479), .B(new_n218), .C1(G33), .C2(new_n243), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n549), .A2(KEYINPUT20), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT20), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n466), .A2(KEYINPUT86), .A3(G270), .A4(new_n282), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n556), .A2(new_n472), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n308), .A2(new_n310), .A3(G264), .A4(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n308), .A2(new_n310), .A3(G257), .A4(new_n270), .ZN(new_n559));
  INV_X1    g0359(.A(G303), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n269), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n276), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n466), .A2(G270), .A3(new_n282), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT86), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n557), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n555), .A2(KEYINPUT21), .A3(G169), .A4(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n557), .A2(new_n562), .A3(G190), .A4(new_n565), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n557), .A2(new_n562), .A3(new_n565), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n554), .B(new_n568), .C1(new_n569), .C2(new_n414), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n291), .B1(new_n561), .B2(new_n276), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n571), .A2(new_n565), .A3(new_n557), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n555), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  OAI21_X1  g0374(.A(G169), .B1(new_n548), .B2(new_n553), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  AND4_X1   g0376(.A1(new_n567), .A2(new_n570), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n276), .B1(new_n463), .B2(new_n471), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G264), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n308), .A2(new_n310), .A3(G257), .A4(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G294), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n308), .A2(new_n310), .A3(G250), .A4(new_n270), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT88), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT88), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n269), .A2(new_n585), .A3(G250), .A4(new_n270), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT89), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n276), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n586), .ZN(new_n590));
  INV_X1    g0390(.A(new_n582), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n590), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n472), .B(new_n579), .C1(new_n589), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n495), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n269), .A2(new_n218), .A3(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT22), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT22), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n269), .A2(new_n597), .A3(new_n218), .A4(G87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n307), .A2(new_n504), .A3(G20), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n218), .B2(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n241), .A2(KEYINPUT23), .A3(G20), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n599), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n600), .B1(new_n599), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n252), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT25), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n249), .B2(G107), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n249), .A2(new_n609), .A3(G107), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n459), .A2(new_n241), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n590), .A2(new_n591), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT89), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n587), .A2(new_n588), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n276), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(new_n291), .A3(new_n472), .A4(new_n579), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n594), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n593), .A2(G200), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(G190), .A3(new_n472), .A4(new_n579), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n608), .A4(new_n614), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n577), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n437), .A2(new_n539), .A3(new_n544), .A4(new_n625), .ZN(G372));
  INV_X1    g0426(.A(KEYINPUT90), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n530), .A2(new_n627), .A3(G200), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n628), .A2(new_n529), .A3(new_n513), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n497), .A2(new_n501), .A3(new_n624), .A4(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n567), .A2(new_n576), .A3(new_n573), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n621), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n537), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n534), .A2(new_n536), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n629), .A2(new_n630), .B1(new_n636), .B2(new_n535), .ZN(new_n637));
  INV_X1    g0437(.A(new_n542), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n493), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n638), .A2(new_n538), .A3(new_n493), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n639), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n437), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n343), .A2(new_n347), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n396), .A2(new_n397), .B1(new_n390), .B2(new_n434), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n365), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n303), .A2(new_n305), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n295), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n649), .ZN(G369));
  AND2_X1   g0450(.A1(new_n624), .A2(new_n621), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n248), .A2(new_n218), .A3(G13), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT91), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(G343), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(G343), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n615), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n651), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n621), .B2(new_n660), .ZN(new_n664));
  INV_X1    g0464(.A(G330), .ZN(new_n665));
  OR3_X1    g0465(.A1(new_n633), .A2(new_n554), .A3(new_n660), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n577), .B1(new_n554), .B2(new_n660), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n633), .A2(new_n661), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n651), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n660), .B(KEYINPUT92), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n621), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0477(.A(new_n212), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n520), .A2(new_n504), .A3(new_n521), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(G1), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n216), .A2(G50), .A3(new_n220), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n680), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT94), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n643), .A2(new_n688), .A3(new_n672), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n641), .A2(new_n639), .ZN(new_n690));
  INV_X1    g0490(.A(new_n637), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT26), .B1(new_n691), .B2(new_n497), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n660), .B1(new_n693), .B2(new_n635), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n506), .A2(new_n512), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n572), .A2(new_n488), .A3(new_n475), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n619), .A2(new_n579), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(G179), .B1(new_n506), .B2(new_n512), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n566), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT95), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n566), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n704), .A2(new_n494), .A3(new_n593), .A4(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n698), .A2(new_n475), .A3(new_n488), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n282), .B1(new_n616), .B2(KEYINPUT89), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(new_n618), .B1(G264), .B2(new_n578), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n708), .A2(new_n710), .A3(KEYINPUT30), .A4(new_n572), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n701), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n661), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n672), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(KEYINPUT96), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT96), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n712), .A2(new_n716), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n712), .B2(new_n661), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n544), .A2(new_n539), .A3(new_n625), .A4(new_n672), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n696), .B1(G330), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n687), .B1(new_n725), .B2(G1), .ZN(G364));
  INV_X1    g0526(.A(new_n668), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n666), .A2(new_n665), .A3(new_n667), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n218), .A2(G13), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n248), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n679), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n269), .A2(G355), .A3(new_n212), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n238), .A2(new_n279), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n678), .A2(new_n269), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n684), .B2(G45), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n735), .B1(G116), .B2(new_n212), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n217), .B1(G20), .B2(new_n495), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n733), .B1(new_n739), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(KEYINPUT97), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(KEYINPUT97), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n414), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n218), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G283), .A2(new_n751), .B1(new_n754), .B2(G329), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n358), .A2(new_n414), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n749), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n755), .B(new_n323), .C1(new_n560), .C2(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(KEYINPUT98), .A2(G20), .A3(G179), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT98), .B1(G20), .B2(G179), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(G190), .A3(new_n414), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n761), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n358), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n768), .A2(G322), .B1(G311), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n218), .B1(new_n766), .B2(new_n291), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n765), .A2(KEYINPUT99), .A3(new_n756), .ZN(new_n777));
  AOI21_X1  g0577(.A(KEYINPUT99), .B1(new_n765), .B2(new_n756), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT101), .B(G326), .Z(new_n780));
  OAI221_X1 g0580(.A(new_n771), .B1(new_n772), .B2(new_n776), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n769), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n782), .A2(new_n272), .B1(new_n328), .B2(new_n767), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G68), .B2(new_n762), .ZN(new_n784));
  INV_X1    g0584(.A(new_n779), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G50), .ZN(new_n786));
  INV_X1    g0586(.A(new_n776), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G97), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n754), .A2(G159), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n269), .B1(new_n750), .B2(new_n241), .C1(new_n520), .C2(new_n757), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n784), .A2(new_n786), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n781), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n746), .B(new_n747), .C1(new_n794), .C2(new_n743), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n666), .A2(new_n667), .A3(new_n742), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n734), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n643), .A2(new_n672), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n409), .A2(new_n661), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n429), .B2(new_n430), .ZN(new_n802));
  INV_X1    g0602(.A(new_n434), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n432), .A2(new_n433), .A3(new_n661), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n805), .B1(new_n802), .B2(new_n803), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n672), .B(new_n809), .C1(new_n635), .C2(new_n642), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n724), .A2(G330), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n732), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n812), .B2(new_n811), .ZN(new_n814));
  INV_X1    g0614(.A(new_n757), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G107), .A2(new_n815), .B1(new_n751), .B2(G87), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n269), .B1(new_n754), .B2(G311), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n782), .A2(new_n504), .B1(new_n772), .B2(new_n767), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G283), .C2(new_n762), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n820), .B(new_n788), .C1(new_n560), .C2(new_n779), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT102), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n768), .A2(G143), .B1(G150), .B2(new_n762), .ZN(new_n823));
  INV_X1    g0623(.A(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n782), .C1(new_n779), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n776), .A2(new_n328), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G68), .A2(new_n751), .B1(new_n754), .B2(G132), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n831), .B(new_n269), .C1(new_n232), .C2(new_n757), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n743), .B1(new_n822), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n743), .A2(new_n740), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n733), .B1(new_n272), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n741), .C2(new_n809), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n814), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT103), .Z(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  NAND2_X1  g0640(.A1(new_n445), .A2(new_n451), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT35), .ZN(new_n842));
  OAI211_X1 g0642(.A(G116), .B(new_n219), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  OR3_X1    g0645(.A1(new_n684), .A2(new_n272), .A3(new_n329), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n248), .B(G13), .C1(new_n846), .C2(new_n233), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n345), .A2(new_n346), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n345), .A2(new_n655), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n361), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n850), .A2(new_n851), .A3(new_n854), .A4(new_n361), .ZN(new_n855));
  INV_X1    g0655(.A(new_n851), .ZN(new_n856));
  AOI221_X4 g0656(.A(new_n849), .B1(new_n853), .B2(new_n855), .C1(new_n367), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n367), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n853), .A2(new_n855), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT39), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT105), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n859), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT104), .B1(new_n363), .B2(new_n364), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n363), .A2(KEYINPUT104), .A3(new_n364), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n645), .A3(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(new_n856), .B1(new_n853), .B2(new_n855), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n863), .B(new_n864), .C1(KEYINPUT38), .C2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n861), .A2(new_n862), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n862), .B1(new_n861), .B2(new_n870), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n396), .A2(new_n397), .A3(new_n660), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n810), .A2(new_n806), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n397), .B(new_n661), .C1(new_n396), .C2(new_n391), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n395), .B1(new_n291), .B2(new_n378), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n394), .B1(new_n378), .B2(G169), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n397), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n388), .A2(new_n660), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n390), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n858), .A2(new_n859), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n849), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n863), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n645), .ZN(new_n891));
  INV_X1    g0691(.A(new_n655), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n877), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n696), .A2(new_n437), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n649), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n807), .B1(new_n879), .B2(new_n885), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n713), .A2(new_n714), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n721), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n723), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n867), .A2(new_n354), .A3(new_n356), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n856), .B1(new_n903), .B2(new_n865), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n904), .B2(new_n859), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n857), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT40), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT40), .B1(new_n889), .B2(new_n863), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n901), .A3(new_n898), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n436), .B1(new_n723), .B2(new_n900), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n665), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n911), .B2(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n897), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n248), .B2(new_n729), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n897), .A2(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n848), .B1(new_n915), .B2(new_n916), .ZN(G367));
  NAND2_X1  g0717(.A1(new_n762), .A2(G294), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT46), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n757), .B2(new_n504), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n918), .B1(KEYINPUT111), .B2(new_n920), .C1(new_n560), .C2(new_n767), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n785), .B2(G311), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n920), .A2(KEYINPUT111), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT112), .B(G317), .Z(new_n924));
  AOI21_X1  g0724(.A(new_n269), .B1(new_n754), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n926), .C1(new_n243), .C2(new_n750), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n923), .B(new_n927), .C1(G283), .C2(new_n769), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n922), .B(new_n928), .C1(new_n241), .C2(new_n776), .ZN(new_n929));
  AOI22_X1  g0729(.A1(G58), .A2(new_n815), .B1(new_n754), .B2(G137), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n767), .B2(new_n262), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G68), .B2(new_n787), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n785), .A2(G143), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n269), .B1(new_n750), .B2(new_n272), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT113), .ZN(new_n935));
  AOI22_X1  g0735(.A1(G50), .A2(new_n769), .B1(new_n762), .B2(G159), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n932), .A2(new_n933), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT47), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n743), .ZN(new_n940));
  INV_X1    g0740(.A(new_n737), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n744), .B1(new_n526), .B2(new_n212), .C1(new_n230), .C2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n942), .A2(KEYINPUT110), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(KEYINPUT110), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n943), .A2(new_n944), .A3(new_n733), .ZN(new_n945));
  INV_X1    g0745(.A(new_n742), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n529), .A2(new_n660), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n636), .A2(new_n947), .A3(new_n535), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n691), .B2(new_n947), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n940), .B(new_n945), .C1(new_n946), .C2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n462), .A2(new_n673), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n497), .A2(new_n501), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n638), .A2(new_n493), .A3(new_n673), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n651), .A3(new_n670), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n497), .B1(new_n953), .B2(new_n621), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n956), .A2(KEYINPUT42), .B1(new_n672), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT107), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(KEYINPUT107), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT108), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n967), .A2(KEYINPUT108), .A3(new_n968), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n965), .C2(new_n964), .ZN(new_n973));
  INV_X1    g0773(.A(new_n955), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n669), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n725), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n675), .A2(new_n955), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n675), .C2(new_n955), .ZN(new_n981));
  NOR2_X1   g0781(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n675), .A2(new_n955), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n669), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n980), .A2(new_n669), .A3(new_n981), .A4(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(new_n727), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n977), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n679), .B(KEYINPUT41), .Z(new_n996));
  OAI21_X1  g0796(.A(new_n730), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n951), .B1(new_n976), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT114), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(G387));
  OR2_X1    g0800(.A1(new_n664), .A2(new_n946), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n737), .B1(new_n227), .B2(new_n279), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n681), .A2(new_n212), .A3(new_n269), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n260), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1005));
  AOI21_X1  g0805(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT50), .B1(new_n260), .B2(G50), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1005), .A2(new_n682), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1004), .A2(new_n1008), .B1(new_n241), .B2(new_n678), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n744), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n732), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n785), .A2(G159), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n787), .A2(new_n406), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n269), .B1(new_n750), .B2(new_n243), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n757), .A2(new_n272), .B1(new_n753), .B2(new_n262), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n260), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1014), .B(new_n1015), .C1(new_n1016), .C2(new_n762), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n768), .A2(G50), .B1(G68), .B2(new_n769), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1012), .A2(new_n1013), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n768), .A2(new_n924), .B1(G311), .B2(new_n762), .ZN(new_n1020));
  INV_X1    g0820(.A(G322), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n560), .B2(new_n782), .C1(new_n779), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G283), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n776), .A2(new_n1025), .B1(new_n772), .B2(new_n757), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n269), .B1(new_n751), .B2(G116), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n780), .C2(new_n753), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT49), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1019), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1011), .B1(new_n1032), .B2(new_n743), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n994), .A2(new_n731), .B1(new_n1001), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n725), .A2(new_n994), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n679), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n725), .A2(new_n994), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  INV_X1    g0838(.A(KEYINPUT115), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n988), .B2(new_n989), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n989), .A2(new_n1039), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n730), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n974), .A2(new_n742), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n246), .A2(new_n737), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n744), .C1(new_n243), .C2(new_n212), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n732), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT116), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n779), .A2(new_n262), .B1(new_n824), .B2(new_n767), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  INV_X1    g0850(.A(G143), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n757), .A2(new_n234), .B1(new_n753), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n323), .B(new_n1052), .C1(G87), .C2(new_n751), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n762), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n232), .C1(new_n260), .C2(new_n782), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n776), .A2(new_n272), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n785), .A2(G317), .B1(G311), .B2(new_n768), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n269), .B1(new_n751), .B2(G107), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G283), .A2(new_n815), .B1(new_n754), .B2(G322), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n1054), .C2(new_n560), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G294), .B2(new_n769), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n504), .B2(new_n776), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1050), .A2(new_n1057), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1048), .B1(new_n1065), .B2(new_n743), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1044), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT117), .B1(new_n1043), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n990), .A2(KEYINPUT115), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n731), .A3(new_n1041), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT117), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1072), .A3(new_n1067), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1035), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n680), .B1(new_n991), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1035), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1078), .ZN(G390));
  AOI21_X1  g0879(.A(new_n864), .B1(new_n889), .B2(new_n863), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n857), .A2(new_n905), .A3(KEYINPUT39), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT105), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n887), .A2(new_n875), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n861), .A2(new_n862), .A3(new_n870), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n660), .B(new_n804), .C1(new_n693), .C2(new_n635), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n806), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n886), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n875), .B1(new_n857), .B2(new_n905), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n724), .A2(G330), .A3(new_n809), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1091), .A2(new_n1089), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1085), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n665), .B1(new_n900), .B2(new_n723), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n898), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n731), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n733), .B1(new_n260), .B2(new_n835), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n323), .B1(new_n754), .B2(G125), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n232), .B2(new_n750), .C1(new_n1054), .C2(new_n825), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G159), .B2(new_n787), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n785), .A2(G128), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n757), .A2(new_n262), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n768), .A2(G132), .B1(new_n769), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1056), .B1(G116), .B2(new_n768), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT121), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G87), .A2(new_n815), .B1(new_n754), .B2(G294), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n323), .C1(new_n234), .C2(new_n750), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G107), .B2(new_n762), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n243), .B2(new_n782), .C1(new_n1025), .C2(new_n779), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(KEYINPUT122), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(KEYINPUT122), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n743), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1099), .B1(new_n1117), .B2(new_n1119), .C1(new_n874), .C2(new_n741), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1094), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1089), .B1(new_n1121), .B2(new_n807), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1092), .A2(new_n1088), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1091), .A2(new_n1089), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1095), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT118), .B1(new_n1125), .B2(new_n878), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1091), .A2(new_n1089), .B1(new_n898), .B2(new_n1094), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT118), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n878), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1095), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n876), .B1(new_n878), .B2(new_n886), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n871), .A2(new_n872), .A3(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n876), .B(new_n906), .C1(new_n886), .C2(new_n1087), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1085), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n895), .B(new_n649), .C1(new_n436), .C2(new_n1121), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1131), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1125), .A2(KEYINPUT118), .A3(new_n878), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1128), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1138), .B1(new_n1145), .B2(new_n1123), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT119), .B1(new_n1097), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT120), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1136), .A2(KEYINPUT120), .A3(new_n1137), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1131), .A2(new_n1139), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n679), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1098), .B(new_n1120), .C1(new_n1148), .C2(new_n1154), .ZN(G378));
  OAI21_X1  g0955(.A(new_n1139), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n910), .A2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n268), .A2(new_n655), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n306), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n306), .A2(new_n1158), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR3_X1    g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1157), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(G330), .A3(new_n910), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n894), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n877), .A2(new_n1166), .A3(new_n893), .A4(new_n1168), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1097), .A2(new_n1146), .A3(KEYINPUT119), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1138), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(KEYINPUT57), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n679), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1165), .A2(new_n740), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n743), .A2(G50), .A3(new_n740), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n269), .A2(G41), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G50), .B(new_n1182), .C1(new_n307), .C2(new_n278), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n782), .A2(new_n526), .B1(new_n241), .B2(new_n767), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G77), .A2(new_n815), .B1(new_n751), .B2(G58), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n1182), .C1(new_n1025), .C2(new_n753), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G97), .C2(new_n762), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n234), .B2(new_n776), .C1(new_n504), .C2(new_n779), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n307), .B(new_n278), .C1(new_n750), .C2(new_n824), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G124), .B2(new_n754), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n768), .A2(G128), .B1(G137), .B2(new_n769), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n762), .A2(G132), .B1(new_n815), .B2(new_n1107), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n262), .C2(new_n776), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G125), .B2(new_n785), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT59), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1192), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1196), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1190), .B1(new_n1189), .B2(new_n1188), .C1(new_n1198), .C2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n733), .B(new_n1181), .C1(new_n1201), .C2(new_n743), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1172), .A2(new_n731), .B1(new_n1180), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1179), .A2(new_n1203), .ZN(G375));
  AOI21_X1  g1004(.A(new_n733), .B1(new_n234), .B2(new_n835), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT123), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G159), .A2(new_n815), .B1(new_n754), .B2(G128), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n269), .C1(new_n328), .C2(new_n750), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G150), .B2(new_n769), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n785), .A2(G132), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n787), .A2(G50), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n768), .A2(G137), .B1(new_n762), .B2(new_n1107), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n779), .A2(new_n772), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n323), .B1(new_n750), .B2(new_n272), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n757), .A2(new_n243), .B1(new_n753), .B2(new_n560), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n769), .C2(G107), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n768), .A2(G283), .B1(G116), .B2(new_n762), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1013), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1213), .B1(new_n1214), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1206), .B1(new_n1220), .B2(new_n743), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n886), .B2(new_n741), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1131), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n730), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1146), .A2(new_n996), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1138), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(G381));
  OR2_X1    g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G384), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G390), .B1(new_n1231), .B2(KEYINPUT124), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(KEYINPUT124), .B2(new_n1231), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(G387), .A2(G381), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1098), .A2(new_n1120), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1154), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G375), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1234), .A2(new_n1238), .A3(new_n1239), .ZN(G407));
  NAND3_X1  g1040(.A1(new_n657), .A2(new_n658), .A3(G213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1238), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  AOI22_X1  g1044(.A1(new_n1069), .A2(new_n1073), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1229), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1246), .B1(new_n1229), .B2(new_n1247), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1245), .B(KEYINPUT114), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1229), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1229), .A2(new_n1247), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT126), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(G390), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1255), .A2(new_n998), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n998), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1203), .C1(new_n1173), .C2(new_n1178), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1172), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1176), .A2(new_n996), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1203), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1238), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1226), .B1(new_n1265), .B2(new_n1146), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1131), .A2(new_n1265), .A3(new_n1139), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n680), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1224), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n839), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n839), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1264), .A2(new_n1241), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1264), .A2(KEYINPUT125), .A3(new_n1241), .A4(new_n1273), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT62), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1279));
  NAND2_X1  g1079(.A1(new_n1264), .A2(new_n1241), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1272), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G2897), .B(new_n1242), .C1(new_n1281), .C2(new_n1270), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1242), .A2(G2897), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1271), .A2(new_n1272), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1279), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1258), .B1(new_n1278), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1276), .A2(new_n1290), .A3(new_n1277), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1274), .A2(new_n1290), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1280), .A2(new_n1285), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1258), .A2(KEYINPUT61), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(new_n1258), .A2(new_n1273), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1272), .B(new_n1271), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1238), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1259), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1299), .B(new_n1301), .ZN(G402));
endmodule


