

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U547 ( .A(n645), .B(n644), .ZN(n667) );
  NOR2_X1 U548 ( .A1(n601), .A2(n600), .ZN(n603) );
  INV_X1 U549 ( .A(KEYINPUT95), .ZN(n620) );
  AND2_X1 U550 ( .A1(n710), .A2(n711), .ZN(n634) );
  INV_X1 U551 ( .A(KEYINPUT29), .ZN(n644) );
  INV_X1 U552 ( .A(KEYINPUT31), .ZN(n654) );
  NAND2_X1 U553 ( .A1(n711), .A2(n710), .ZN(n647) );
  INV_X1 U554 ( .A(n759), .ZN(n746) );
  AND2_X1 U555 ( .A1(n747), .A2(n746), .ZN(n748) );
  INV_X1 U556 ( .A(G651), .ZN(n525) );
  XOR2_X1 U557 ( .A(KEYINPUT73), .B(n614), .Z(n902) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n516), .ZN(n892) );
  NOR2_X1 U559 ( .A1(G651), .A2(n526), .ZN(n795) );
  NAND2_X1 U560 ( .A1(n603), .A2(n602), .ZN(n946) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n511) );
  XOR2_X2 U562 ( .A(KEYINPUT17), .B(n511), .Z(n890) );
  NAND2_X1 U563 ( .A1(n890), .A2(G138), .ZN(n514) );
  INV_X1 U564 ( .A(G2104), .ZN(n516) );
  NAND2_X1 U565 ( .A1(G102), .A2(n892), .ZN(n512) );
  XOR2_X1 U566 ( .A(KEYINPUT83), .B(n512), .Z(n513) );
  NAND2_X1 U567 ( .A1(n514), .A2(n513), .ZN(n520) );
  INV_X1 U568 ( .A(G2105), .ZN(n515) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n515), .ZN(n886) );
  NAND2_X1 U570 ( .A1(G126), .A2(n886), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n516), .A2(n515), .ZN(n887) );
  NAND2_X1 U572 ( .A1(G114), .A2(n887), .ZN(n517) );
  NAND2_X1 U573 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U574 ( .A1(n520), .A2(n519), .ZN(G164) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n526) );
  NAND2_X1 U576 ( .A1(n795), .A2(G52), .ZN(n524) );
  NOR2_X1 U577 ( .A1(G543), .A2(n525), .ZN(n521) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n521), .Z(n522) );
  XNOR2_X2 U579 ( .A(KEYINPUT66), .B(n522), .ZN(n796) );
  NAND2_X1 U580 ( .A1(G64), .A2(n796), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n531) );
  NOR2_X1 U582 ( .A1(n526), .A2(n525), .ZN(n799) );
  NAND2_X1 U583 ( .A1(G77), .A2(n799), .ZN(n528) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n800) );
  NAND2_X1 U585 ( .A1(G90), .A2(n800), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(n529), .Z(n530) );
  NOR2_X1 U588 ( .A1(n531), .A2(n530), .ZN(G171) );
  NAND2_X1 U589 ( .A1(n799), .A2(G75), .ZN(n534) );
  NAND2_X1 U590 ( .A1(G50), .A2(n795), .ZN(n532) );
  XOR2_X1 U591 ( .A(KEYINPUT81), .B(n532), .Z(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n800), .A2(G88), .ZN(n536) );
  NAND2_X1 U594 ( .A1(G62), .A2(n796), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n538), .A2(n537), .ZN(G166) );
  XOR2_X1 U597 ( .A(KEYINPUT84), .B(G166), .Z(G303) );
  INV_X1 U598 ( .A(KEYINPUT7), .ZN(n550) );
  NAND2_X1 U599 ( .A1(G63), .A2(n796), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n539), .B(KEYINPUT74), .ZN(n541) );
  NAND2_X1 U601 ( .A1(G51), .A2(n795), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT6), .B(n542), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n800), .A2(G89), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT4), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G76), .A2(n799), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U608 ( .A(n546), .B(KEYINPUT5), .Z(n547) );
  NOR2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT75), .B(n551), .Z(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G87), .A2(n526), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G74), .A2(G651), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U616 ( .A1(n796), .A2(n554), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n795), .A2(G49), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G288) );
  NAND2_X1 U619 ( .A1(n799), .A2(G73), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT2), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G86), .A2(n800), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G61), .A2(n796), .ZN(n560) );
  XNOR2_X1 U624 ( .A(KEYINPUT79), .B(n560), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT80), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G48), .A2(n795), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(G305) );
  AND2_X1 U629 ( .A1(G60), .A2(n796), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G72), .A2(n799), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G85), .A2(n800), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n795), .A2(G47), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(G290) );
  INV_X1 U636 ( .A(KEYINPUT85), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n892), .A2(G101), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT23), .B(n572), .Z(n574) );
  NAND2_X1 U639 ( .A1(n886), .A2(G125), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT65), .ZN(n768) );
  NAND2_X1 U642 ( .A1(G137), .A2(n890), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G113), .A2(n887), .ZN(n576) );
  AND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n769) );
  AND2_X1 U645 ( .A1(n769), .A2(G40), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n768), .A2(n578), .ZN(n581) );
  INV_X1 U647 ( .A(n581), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U649 ( .A1(KEYINPUT85), .A2(n581), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n710) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NOR2_X1 U652 ( .A1(n634), .A2(G1961), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT93), .ZN(n586) );
  XNOR2_X1 U654 ( .A(G2078), .B(KEYINPUT25), .ZN(n933) );
  NAND2_X1 U655 ( .A1(n634), .A2(n933), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n651) );
  NAND2_X1 U657 ( .A1(n651), .A2(G171), .ZN(n668) );
  NAND2_X1 U658 ( .A1(G8), .A2(n647), .ZN(n727) );
  NOR2_X1 U659 ( .A1(G1971), .A2(n727), .ZN(n588) );
  NOR2_X1 U660 ( .A1(G2090), .A2(n647), .ZN(n587) );
  NOR2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n589), .A2(G303), .ZN(n656) );
  INV_X1 U663 ( .A(n656), .ZN(n590) );
  OR2_X1 U664 ( .A1(n590), .A2(G286), .ZN(n658) );
  AND2_X1 U665 ( .A1(n668), .A2(n658), .ZN(n646) );
  XNOR2_X1 U666 ( .A(G1996), .B(KEYINPUT94), .ZN(n928) );
  NAND2_X1 U667 ( .A1(n928), .A2(n634), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n591), .B(KEYINPUT26), .ZN(n623) );
  XOR2_X1 U669 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n593) );
  NAND2_X1 U670 ( .A1(G56), .A2(n796), .ZN(n592) );
  XNOR2_X1 U671 ( .A(n593), .B(n592), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n799), .A2(G68), .ZN(n594) );
  XNOR2_X1 U673 ( .A(n594), .B(KEYINPUT70), .ZN(n598) );
  XOR2_X1 U674 ( .A(KEYINPUT69), .B(KEYINPUT12), .Z(n596) );
  NAND2_X1 U675 ( .A1(G81), .A2(n800), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U678 ( .A(KEYINPUT13), .B(n599), .Z(n600) );
  NAND2_X1 U679 ( .A1(n795), .A2(G43), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n647), .A2(G1341), .ZN(n622) );
  INV_X1 U681 ( .A(n622), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n946), .A2(n604), .ZN(n605) );
  AND2_X1 U683 ( .A1(n623), .A2(n605), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n796), .A2(G66), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT72), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G79), .A2(n799), .ZN(n608) );
  NAND2_X1 U687 ( .A1(G92), .A2(n800), .ZN(n607) );
  AND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G54), .A2(n795), .ZN(n609) );
  AND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT15), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n902), .ZN(n619) );
  NOR2_X1 U694 ( .A1(G2067), .A2(n647), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n634), .A2(G1348), .ZN(n616) );
  NOR2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(n620), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n946), .A2(n624), .ZN(n625) );
  OR2_X1 U701 ( .A1(n902), .A2(n625), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n639) );
  NAND2_X1 U703 ( .A1(n795), .A2(G53), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G65), .A2(n796), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G78), .A2(n799), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G91), .A2(n800), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n947) );
  NAND2_X1 U710 ( .A1(n634), .A2(G2072), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT27), .ZN(n637) );
  AND2_X1 U712 ( .A1(G1956), .A2(n647), .ZN(n636) );
  NOR2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n947), .A2(n640), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n947), .A2(n640), .ZN(n641) );
  XOR2_X1 U717 ( .A(n641), .B(KEYINPUT28), .Z(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n667), .ZN(n660) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n727), .ZN(n672) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n647), .ZN(n665) );
  NOR2_X1 U722 ( .A1(n672), .A2(n665), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G8), .A2(n648), .ZN(n649) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n649), .ZN(n650) );
  NOR2_X1 U725 ( .A1(n650), .A2(G168), .ZN(n653) );
  NOR2_X1 U726 ( .A1(G171), .A2(n651), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(n669) );
  NAND2_X1 U729 ( .A1(n669), .A2(n656), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n661), .B(KEYINPUT96), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n662), .A2(G8), .ZN(n664) );
  XOR2_X1 U734 ( .A(KEYINPUT97), .B(KEYINPUT32), .Z(n663) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(n719) );
  NAND2_X1 U736 ( .A1(G8), .A2(n665), .ZN(n666) );
  XNOR2_X1 U737 ( .A(KEYINPUT92), .B(n666), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n670) );
  AND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n718) );
  NAND2_X1 U742 ( .A1(G288), .A2(G1976), .ZN(n675) );
  XOR2_X1 U743 ( .A(KEYINPUT99), .B(n675), .Z(n953) );
  INV_X1 U744 ( .A(n953), .ZN(n676) );
  OR2_X1 U745 ( .A1(n676), .A2(n727), .ZN(n683) );
  INV_X1 U746 ( .A(n683), .ZN(n677) );
  AND2_X1 U747 ( .A1(n718), .A2(n677), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n719), .A2(n678), .ZN(n685) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n679) );
  XOR2_X1 U750 ( .A(KEYINPUT98), .B(n679), .Z(n950) );
  INV_X1 U751 ( .A(n950), .ZN(n681) );
  NOR2_X1 U752 ( .A1(G303), .A2(G1971), .ZN(n680) );
  NOR2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n682) );
  OR2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n687) );
  INV_X1 U756 ( .A(KEYINPUT64), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n687), .B(n686), .ZN(n689) );
  INV_X1 U758 ( .A(KEYINPUT33), .ZN(n688) );
  NAND2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n717) );
  NOR2_X1 U760 ( .A1(n950), .A2(n727), .ZN(n690) );
  NAND2_X1 U761 ( .A1(KEYINPUT33), .A2(n690), .ZN(n691) );
  XOR2_X1 U762 ( .A(G1981), .B(G305), .Z(n955) );
  NAND2_X1 U763 ( .A1(n691), .A2(n955), .ZN(n715) );
  NAND2_X1 U764 ( .A1(G129), .A2(n886), .ZN(n693) );
  NAND2_X1 U765 ( .A1(G117), .A2(n887), .ZN(n692) );
  NAND2_X1 U766 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n892), .A2(G105), .ZN(n694) );
  XOR2_X1 U768 ( .A(KEYINPUT38), .B(n694), .Z(n695) );
  NOR2_X1 U769 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n890), .A2(G141), .ZN(n697) );
  NAND2_X1 U771 ( .A1(n698), .A2(n697), .ZN(n871) );
  NAND2_X1 U772 ( .A1(G1996), .A2(n871), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n699), .B(KEYINPUT90), .ZN(n709) );
  NAND2_X1 U774 ( .A1(G107), .A2(n887), .ZN(n700) );
  XOR2_X1 U775 ( .A(KEYINPUT88), .B(n700), .Z(n705) );
  NAND2_X1 U776 ( .A1(G95), .A2(n892), .ZN(n702) );
  NAND2_X1 U777 ( .A1(G131), .A2(n890), .ZN(n701) );
  NAND2_X1 U778 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U779 ( .A(KEYINPUT89), .B(n703), .Z(n704) );
  NOR2_X1 U780 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U781 ( .A1(n886), .A2(G119), .ZN(n706) );
  NAND2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n872) );
  NAND2_X1 U783 ( .A1(G1991), .A2(n872), .ZN(n708) );
  NAND2_X1 U784 ( .A1(n709), .A2(n708), .ZN(n1009) );
  INV_X1 U785 ( .A(n710), .ZN(n712) );
  NOR2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U787 ( .A(n713), .B(KEYINPUT86), .ZN(n763) );
  NAND2_X1 U788 ( .A1(n1009), .A2(n763), .ZN(n714) );
  XNOR2_X1 U789 ( .A(n714), .B(KEYINPUT91), .ZN(n754) );
  NOR2_X1 U790 ( .A1(n715), .A2(n754), .ZN(n716) );
  NAND2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n734) );
  INV_X1 U792 ( .A(n754), .ZN(n732) );
  NAND2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n725) );
  NOR2_X1 U794 ( .A1(G2090), .A2(G303), .ZN(n720) );
  NAND2_X1 U795 ( .A1(G8), .A2(n720), .ZN(n723) );
  NOR2_X1 U796 ( .A1(G1981), .A2(G305), .ZN(n721) );
  XOR2_X1 U797 ( .A(n721), .B(KEYINPUT24), .Z(n722) );
  OR2_X1 U798 ( .A1(n727), .A2(n722), .ZN(n726) );
  AND2_X1 U799 ( .A1(n723), .A2(n726), .ZN(n724) );
  NAND2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n730) );
  INV_X1 U801 ( .A(n726), .ZN(n728) );
  OR2_X1 U802 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n747) );
  INV_X1 U806 ( .A(n763), .ZN(n745) );
  XNOR2_X1 U807 ( .A(G2067), .B(KEYINPUT37), .ZN(n761) );
  NAND2_X1 U808 ( .A1(G128), .A2(n886), .ZN(n736) );
  NAND2_X1 U809 ( .A1(G116), .A2(n887), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U811 ( .A(n737), .B(KEYINPUT35), .ZN(n742) );
  NAND2_X1 U812 ( .A1(G104), .A2(n892), .ZN(n739) );
  NAND2_X1 U813 ( .A1(G140), .A2(n890), .ZN(n738) );
  NAND2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U815 ( .A(KEYINPUT34), .B(n740), .Z(n741) );
  NAND2_X1 U816 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U817 ( .A(n743), .B(KEYINPUT36), .Z(n868) );
  OR2_X1 U818 ( .A1(n761), .A2(n868), .ZN(n744) );
  XOR2_X1 U819 ( .A(KEYINPUT87), .B(n744), .Z(n1017) );
  NOR2_X1 U820 ( .A1(n745), .A2(n1017), .ZN(n759) );
  XNOR2_X1 U821 ( .A(n748), .B(KEYINPUT100), .ZN(n750) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n962) );
  NAND2_X1 U823 ( .A1(n962), .A2(n763), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n766) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n871), .ZN(n1005) );
  NOR2_X1 U826 ( .A1(G1991), .A2(n872), .ZN(n1023) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n1023), .A2(n751), .ZN(n752) );
  XOR2_X1 U829 ( .A(KEYINPUT101), .B(n752), .Z(n753) );
  NOR2_X1 U830 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U831 ( .A(n755), .B(KEYINPUT102), .ZN(n756) );
  NOR2_X1 U832 ( .A1(n1005), .A2(n756), .ZN(n757) );
  XOR2_X1 U833 ( .A(KEYINPUT39), .B(n757), .Z(n758) );
  NOR2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U835 ( .A(n760), .B(KEYINPUT103), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n868), .A2(n761), .ZN(n1022) );
  NAND2_X1 U837 ( .A1(n762), .A2(n1022), .ZN(n764) );
  NAND2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n767), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U841 ( .A1(n769), .A2(n768), .ZN(G160) );
  NAND2_X1 U842 ( .A1(G123), .A2(n886), .ZN(n770) );
  XOR2_X1 U843 ( .A(KEYINPUT18), .B(n770), .Z(n775) );
  NAND2_X1 U844 ( .A1(G99), .A2(n892), .ZN(n772) );
  NAND2_X1 U845 ( .A1(G111), .A2(n887), .ZN(n771) );
  NAND2_X1 U846 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U847 ( .A(KEYINPUT77), .B(n773), .Z(n774) );
  NOR2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U849 ( .A1(n890), .A2(G135), .ZN(n776) );
  NAND2_X1 U850 ( .A1(n777), .A2(n776), .ZN(n1021) );
  XNOR2_X1 U851 ( .A(G2096), .B(n1021), .ZN(n778) );
  OR2_X1 U852 ( .A1(G2100), .A2(n778), .ZN(G156) );
  INV_X1 U853 ( .A(G57), .ZN(G237) );
  INV_X1 U854 ( .A(G132), .ZN(G219) );
  INV_X1 U855 ( .A(G82), .ZN(G220) );
  NAND2_X1 U856 ( .A1(G94), .A2(G452), .ZN(n779) );
  XNOR2_X1 U857 ( .A(n779), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n780) );
  XNOR2_X1 U859 ( .A(n780), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U860 ( .A(G223), .ZN(n830) );
  NAND2_X1 U861 ( .A1(n830), .A2(G567), .ZN(n781) );
  XOR2_X1 U862 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  XNOR2_X1 U863 ( .A(G860), .B(KEYINPUT71), .ZN(n786) );
  OR2_X1 U864 ( .A1(n946), .A2(n786), .ZN(G153) );
  INV_X1 U865 ( .A(G171), .ZN(G301) );
  NAND2_X1 U866 ( .A1(G868), .A2(G301), .ZN(n783) );
  INV_X1 U867 ( .A(n902), .ZN(n963) );
  INV_X1 U868 ( .A(G868), .ZN(n815) );
  NAND2_X1 U869 ( .A1(n963), .A2(n815), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(G284) );
  INV_X1 U871 ( .A(n947), .ZN(G299) );
  NOR2_X1 U872 ( .A1(G286), .A2(n815), .ZN(n785) );
  NOR2_X1 U873 ( .A1(G868), .A2(G299), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n786), .A2(G559), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n787), .A2(n902), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n788), .B(KEYINPUT76), .ZN(n789) );
  XNOR2_X1 U878 ( .A(KEYINPUT16), .B(n789), .ZN(G148) );
  NOR2_X1 U879 ( .A1(G868), .A2(n946), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G868), .A2(n902), .ZN(n790) );
  NOR2_X1 U881 ( .A1(G559), .A2(n790), .ZN(n791) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(G282) );
  XNOR2_X1 U883 ( .A(n946), .B(KEYINPUT78), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n902), .A2(G559), .ZN(n793) );
  XNOR2_X1 U885 ( .A(n794), .B(n793), .ZN(n812) );
  NOR2_X1 U886 ( .A1(G860), .A2(n812), .ZN(n805) );
  NAND2_X1 U887 ( .A1(n795), .A2(G55), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G67), .A2(n796), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G80), .A2(n799), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G93), .A2(n800), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n814) );
  XOR2_X1 U894 ( .A(n805), .B(n814), .Z(G145) );
  XNOR2_X1 U895 ( .A(n947), .B(G290), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n806), .B(G305), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n807) );
  XNOR2_X1 U898 ( .A(G288), .B(n807), .ZN(n808) );
  XOR2_X1 U899 ( .A(n809), .B(n808), .Z(n811) );
  XOR2_X1 U900 ( .A(G166), .B(n814), .Z(n810) );
  XNOR2_X1 U901 ( .A(n811), .B(n810), .ZN(n901) );
  XNOR2_X1 U902 ( .A(n812), .B(n901), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n822) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n822), .Z(n823) );
  NOR2_X1 U914 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G96), .A2(n824), .ZN(n834) );
  NAND2_X1 U916 ( .A1(n834), .A2(G2106), .ZN(n828) );
  NAND2_X1 U917 ( .A1(G108), .A2(G120), .ZN(n825) );
  NOR2_X1 U918 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U919 ( .A1(G69), .A2(n826), .ZN(n835) );
  NAND2_X1 U920 ( .A1(n835), .A2(G567), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n857) );
  NAND2_X1 U922 ( .A1(G661), .A2(G483), .ZN(n829) );
  NOR2_X1 U923 ( .A1(n857), .A2(n829), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U927 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U930 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  XNOR2_X1 U932 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  XOR2_X1 U936 ( .A(KEYINPUT110), .B(G2678), .Z(n837) );
  XNOR2_X1 U937 ( .A(KEYINPUT43), .B(G2096), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n838), .B(KEYINPUT42), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2072), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U942 ( .A(G2100), .B(G2090), .Z(n842) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2084), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U946 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1971), .B(G1961), .Z(n848) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U951 ( .A(G1976), .B(G1956), .Z(n850) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U953 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U954 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(G2474), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U957 ( .A(G1981), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G229) );
  INV_X1 U959 ( .A(n857), .ZN(G319) );
  NAND2_X1 U960 ( .A1(G124), .A2(n886), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n892), .A2(G100), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G136), .A2(n890), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G112), .A2(n887), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n1021), .B(n867), .ZN(n870) );
  XOR2_X1 U972 ( .A(G164), .B(n868), .Z(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n875) );
  XNOR2_X1 U974 ( .A(G162), .B(n871), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U976 ( .A(n875), .B(n874), .Z(n885) );
  NAND2_X1 U977 ( .A1(G103), .A2(n892), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G139), .A2(n890), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n887), .A2(G115), .ZN(n878) );
  XOR2_X1 U981 ( .A(KEYINPUT113), .B(n878), .Z(n880) );
  NAND2_X1 U982 ( .A1(n886), .A2(G127), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n1012) );
  XNOR2_X1 U986 ( .A(G160), .B(n1012), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n899) );
  NAND2_X1 U988 ( .A1(G130), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G118), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n897) );
  NAND2_X1 U991 ( .A1(n890), .A2(G142), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n891), .B(KEYINPUT112), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G106), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(n895), .B(KEYINPUT45), .Z(n896) );
  NOR2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U998 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U999 ( .A(n901), .B(G286), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G171), .B(n902), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n905), .B(n946), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n921) );
  XNOR2_X1 U1007 ( .A(G2451), .B(G2446), .ZN(n918) );
  XOR2_X1 U1008 ( .A(G2430), .B(KEYINPUT105), .Z(n910) );
  XNOR2_X1 U1009 ( .A(G2454), .B(G2435), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1011 ( .A(G2438), .B(KEYINPUT104), .Z(n912) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1014 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1015 ( .A(G2443), .B(G2427), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(G14), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n924), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(n924), .ZN(G401) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n1029) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G35), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(G1991), .B(G25), .ZN(n926) );
  XNOR2_X1 U1029 ( .A(G33), .B(G2072), .ZN(n925) );
  NOR2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1031 ( .A(G2067), .B(G26), .Z(n927) );
  NAND2_X1 U1032 ( .A1(n927), .A2(G28), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(G32), .B(n928), .ZN(n929) );
  NOR2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1036 ( .A(G27), .B(n933), .Z(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(KEYINPUT53), .B(n936), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n941) );
  XOR2_X1 U1040 ( .A(G2084), .B(G34), .Z(n939) );
  XNOR2_X1 U1041 ( .A(KEYINPUT54), .B(n939), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(n1029), .B(n942), .ZN(n944) );
  INV_X1 U1044 ( .A(G29), .ZN(n943) );
  NAND2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n945), .ZN(n1003) );
  XNOR2_X1 U1047 ( .A(G16), .B(KEYINPUT56), .ZN(n973) );
  XOR2_X1 U1048 ( .A(n946), .B(G1341), .Z(n949) );
  XNOR2_X1 U1049 ( .A(n947), .B(G1956), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1051 ( .A(n950), .B(KEYINPUT122), .Z(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n957), .B(KEYINPUT120), .ZN(n958) );
  XOR2_X1 U1057 ( .A(KEYINPUT57), .B(n958), .Z(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(G1961), .B(G301), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT121), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(n964), .B(n963), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1064 ( .A(G1971), .B(G303), .Z(n967) );
  XNOR2_X1 U1065 ( .A(KEYINPUT123), .B(n967), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n1001) );
  INV_X1 U1069 ( .A(G16), .ZN(n999) );
  XNOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n974), .B(G4), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G1341), .B(G19), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G20), .ZN(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT125), .B(G1981), .Z(n979) );
  XNOR2_X1 U1077 ( .A(G6), .B(n979), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(KEYINPUT60), .B(n982), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(G1976), .B(G23), .ZN(n983) );
  NOR2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1083 ( .A(KEYINPUT126), .B(n985), .Z(n987) );
  XNOR2_X1 U1084 ( .A(G1986), .B(G24), .ZN(n986) );
  NOR2_X1 U1085 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1086 ( .A(n988), .B(KEYINPUT58), .ZN(n989) );
  XNOR2_X1 U1087 ( .A(n989), .B(KEYINPUT127), .ZN(n992) );
  XNOR2_X1 U1088 ( .A(KEYINPUT124), .B(G1961), .ZN(n990) );
  XNOR2_X1 U1089 ( .A(G5), .B(n990), .ZN(n991) );
  NOR2_X1 U1090 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1092 ( .A(G21), .B(G1966), .ZN(n995) );
  NOR2_X1 U1093 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1094 ( .A(KEYINPUT61), .B(n997), .ZN(n998) );
  NAND2_X1 U1095 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1096 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1033) );
  XNOR2_X1 U1098 ( .A(G160), .B(G2084), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1100 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1006), .Z(n1007) );
  XNOR2_X1 U1102 ( .A(n1007), .B(KEYINPUT117), .ZN(n1008) );
  NOR2_X1 U1103 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1104 ( .A1(n1011), .A2(n1010), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1015) );
  XOR2_X1 U1106 ( .A(n1012), .B(KEYINPUT118), .Z(n1013) );
  XNOR2_X1 U1107 ( .A(G2072), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1108 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1109 ( .A(n1016), .B(KEYINPUT50), .ZN(n1018) );
  NAND2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT119), .B(n1027), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT52), .B(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(G29), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

