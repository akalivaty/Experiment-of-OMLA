

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596;

  INV_X1 U324 ( .A(KEYINPUT55), .ZN(n460) );
  INV_X1 U325 ( .A(n525), .ZN(n497) );
  XNOR2_X1 U326 ( .A(G36GAT), .B(G190GAT), .ZN(n408) );
  XNOR2_X1 U327 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U328 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U329 ( .A1(n497), .A2(n496), .ZN(n498) );
  XOR2_X1 U330 ( .A(n458), .B(n457), .Z(n556) );
  XOR2_X1 U331 ( .A(KEYINPUT40), .B(n507), .Z(n292) );
  XOR2_X1 U332 ( .A(n361), .B(n360), .Z(n293) );
  XNOR2_X1 U333 ( .A(n414), .B(KEYINPUT114), .ZN(n415) );
  XNOR2_X1 U334 ( .A(n416), .B(n415), .ZN(n422) );
  XNOR2_X1 U335 ( .A(n430), .B(n429), .ZN(n431) );
  INV_X1 U336 ( .A(n495), .ZN(n496) );
  XNOR2_X1 U337 ( .A(n362), .B(n293), .ZN(n363) );
  XNOR2_X1 U338 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U339 ( .A(n364), .B(n363), .ZN(n367) );
  XNOR2_X1 U340 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XOR2_X1 U341 ( .A(n437), .B(n436), .Z(n504) );
  XNOR2_X1 U342 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n465) );
  XNOR2_X1 U343 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(G176GAT), .B(KEYINPUT20), .Z(n295) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(KEYINPUT87), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n311) );
  XOR2_X1 U347 ( .A(KEYINPUT18), .B(KEYINPUT85), .Z(n297) );
  XNOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(KEYINPUT17), .B(n298), .Z(n434) );
  XOR2_X1 U351 ( .A(G15GAT), .B(G127GAT), .Z(n376) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n299), .B(KEYINPUT0), .ZN(n450) );
  XOR2_X1 U354 ( .A(n376), .B(n450), .Z(n301) );
  NAND2_X1 U355 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n434), .B(n302), .ZN(n309) );
  XOR2_X1 U358 ( .A(G183GAT), .B(KEYINPUT88), .Z(n304) );
  XNOR2_X1 U359 ( .A(G190GAT), .B(G99GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U361 ( .A(n305), .B(KEYINPUT84), .Z(n307) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n365) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(n365), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X2 U366 ( .A(n311), .B(n310), .Z(n540) );
  INV_X1 U367 ( .A(n540), .ZN(n506) );
  XNOR2_X1 U368 ( .A(G211GAT), .B(G218GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n312), .B(KEYINPUT21), .ZN(n313) );
  XOR2_X1 U370 ( .A(n313), .B(KEYINPUT89), .Z(n315) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G204GAT), .ZN(n314) );
  XOR2_X1 U372 ( .A(n315), .B(n314), .Z(n435) );
  XOR2_X1 U373 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n317) );
  XNOR2_X1 U374 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U376 ( .A(KEYINPUT3), .B(n318), .Z(n449) );
  XOR2_X1 U377 ( .A(n435), .B(n449), .Z(n331) );
  XOR2_X1 U378 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n320) );
  XNOR2_X1 U379 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U381 ( .A(KEYINPUT92), .B(n321), .Z(n323) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n326) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G148GAT), .Z(n325) );
  XNOR2_X1 U385 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n359) );
  XOR2_X1 U387 ( .A(n326), .B(n359), .Z(n329) );
  XOR2_X1 U388 ( .A(G141GAT), .B(G22GAT), .Z(n334) );
  XNOR2_X1 U389 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n327), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U391 ( .A(n334), .B(n409), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n474) );
  XOR2_X1 U394 ( .A(G169GAT), .B(G8GAT), .Z(n429) );
  XOR2_X1 U395 ( .A(KEYINPUT69), .B(G1GAT), .Z(n378) );
  XOR2_X1 U396 ( .A(n429), .B(n378), .Z(n333) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n335) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U400 ( .A(G15GAT), .B(G113GAT), .Z(n337) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(G36GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U403 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n339) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U406 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n345) );
  INV_X1 U408 ( .A(KEYINPUT68), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U410 ( .A(G29GAT), .B(G43GAT), .Z(n347) );
  XNOR2_X1 U411 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n403) );
  XNOR2_X1 U413 ( .A(n403), .B(KEYINPUT30), .ZN(n348) );
  XOR2_X1 U414 ( .A(n349), .B(n348), .Z(n541) );
  INV_X1 U415 ( .A(n541), .ZN(n581) );
  XOR2_X1 U416 ( .A(G99GAT), .B(G85GAT), .Z(n402) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(G92GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n350), .B(G64GAT), .ZN(n428) );
  XNOR2_X1 U419 ( .A(n402), .B(n428), .ZN(n354) );
  INV_X1 U420 ( .A(n354), .ZN(n352) );
  AND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  INV_X1 U422 ( .A(n353), .ZN(n351) );
  NAND2_X1 U423 ( .A1(n352), .A2(n351), .ZN(n356) );
  NAND2_X1 U424 ( .A1(n354), .A2(n353), .ZN(n355) );
  NAND2_X1 U425 ( .A1(n356), .A2(n355), .ZN(n358) );
  INV_X1 U426 ( .A(KEYINPUT31), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n359), .B(KEYINPUT71), .ZN(n362) );
  XOR2_X1 U429 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n361) );
  XNOR2_X1 U430 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n360) );
  XOR2_X1 U431 ( .A(G57GAT), .B(KEYINPUT13), .Z(n377) );
  XNOR2_X1 U432 ( .A(n365), .B(n377), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n586) );
  XNOR2_X1 U434 ( .A(n586), .B(KEYINPUT41), .ZN(n512) );
  NAND2_X1 U435 ( .A1(n581), .A2(n512), .ZN(n370) );
  XOR2_X1 U436 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n368) );
  XNOR2_X1 U437 ( .A(KEYINPUT112), .B(n368), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n413) );
  XOR2_X1 U439 ( .A(KEYINPUT80), .B(G64GAT), .Z(n372) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(G155GAT), .ZN(n371) );
  XNOR2_X1 U441 ( .A(n372), .B(n371), .ZN(n390) );
  XOR2_X1 U442 ( .A(G183GAT), .B(KEYINPUT79), .Z(n427) );
  XOR2_X1 U443 ( .A(n427), .B(KEYINPUT12), .Z(n374) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n388) );
  XOR2_X1 U447 ( .A(n377), .B(G78GAT), .Z(n380) );
  XNOR2_X1 U448 ( .A(n378), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U450 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n382) );
  XNOR2_X1 U451 ( .A(KEYINPUT14), .B(KEYINPUT81), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U453 ( .A(n384), .B(n383), .Z(n386) );
  XNOR2_X1 U454 ( .A(G22GAT), .B(G71GAT), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U457 ( .A(n390), .B(n389), .Z(n589) );
  INV_X1 U458 ( .A(n589), .ZN(n548) );
  XOR2_X1 U459 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n392) );
  XNOR2_X1 U460 ( .A(KEYINPUT75), .B(KEYINPUT78), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U462 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n394) );
  XNOR2_X1 U463 ( .A(G134GAT), .B(G92GAT), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U465 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U466 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n398) );
  NAND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U469 ( .A(G106GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n401), .B(n400), .ZN(n407) );
  XOR2_X1 U471 ( .A(KEYINPUT74), .B(n402), .Z(n405) );
  XNOR2_X1 U472 ( .A(n403), .B(G218GAT), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U474 ( .A(n407), .B(n406), .Z(n411) );
  XNOR2_X1 U475 ( .A(n408), .B(KEYINPUT77), .ZN(n424) );
  XNOR2_X1 U476 ( .A(n409), .B(n424), .ZN(n410) );
  XOR2_X1 U477 ( .A(n411), .B(n410), .Z(n552) );
  AND2_X1 U478 ( .A1(n548), .A2(n552), .ZN(n412) );
  AND2_X1 U479 ( .A1(n413), .A2(n412), .ZN(n416) );
  INV_X1 U480 ( .A(KEYINPUT47), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n552), .B(KEYINPUT102), .ZN(n417) );
  XNOR2_X1 U482 ( .A(KEYINPUT36), .B(n417), .ZN(n594) );
  NOR2_X1 U483 ( .A1(n594), .A2(n548), .ZN(n418) );
  XNOR2_X1 U484 ( .A(KEYINPUT45), .B(n418), .ZN(n419) );
  NAND2_X1 U485 ( .A1(n419), .A2(n586), .ZN(n420) );
  NOR2_X1 U486 ( .A1(n420), .A2(n581), .ZN(n421) );
  NOR2_X1 U487 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(KEYINPUT48), .B(n423), .ZN(n537) );
  XOR2_X1 U489 ( .A(KEYINPUT97), .B(n424), .Z(n426) );
  NAND2_X1 U490 ( .A1(G226GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U492 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n437) );
  INV_X1 U494 ( .A(n435), .ZN(n436) );
  NOR2_X1 U495 ( .A1(n537), .A2(n504), .ZN(n438) );
  XNOR2_X1 U496 ( .A(KEYINPUT54), .B(n438), .ZN(n459) );
  XOR2_X1 U497 ( .A(G120GAT), .B(G127GAT), .Z(n440) );
  XNOR2_X1 U498 ( .A(G29GAT), .B(G141GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U500 ( .A(G162GAT), .B(G85GAT), .Z(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n456) );
  XOR2_X1 U502 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n444) );
  XNOR2_X1 U503 ( .A(KEYINPUT6), .B(KEYINPUT95), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U505 ( .A(KEYINPUT94), .B(G57GAT), .Z(n446) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(G148GAT), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n454) );
  XOR2_X1 U509 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n452) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n458) );
  NAND2_X1 U514 ( .A1(G225GAT), .A2(G233GAT), .ZN(n457) );
  INV_X1 U515 ( .A(n556), .ZN(n500) );
  NAND2_X1 U516 ( .A1(n459), .A2(n500), .ZN(n579) );
  NOR2_X1 U517 ( .A1(n474), .A2(n579), .ZN(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n506), .A2(n464), .ZN(n576) );
  INV_X1 U520 ( .A(n552), .ZN(n566) );
  NAND2_X1 U521 ( .A1(n576), .A2(n566), .ZN(n466) );
  XNOR2_X1 U522 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n484) );
  NAND2_X1 U523 ( .A1(n581), .A2(n586), .ZN(n495) );
  INV_X1 U524 ( .A(n504), .ZN(n528) );
  XOR2_X1 U525 ( .A(KEYINPUT27), .B(n528), .Z(n475) );
  NAND2_X1 U526 ( .A1(n506), .A2(n474), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT98), .ZN(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT26), .B(n468), .ZN(n578) );
  NOR2_X1 U529 ( .A1(n475), .A2(n578), .ZN(n557) );
  NOR2_X1 U530 ( .A1(n506), .A2(n504), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n469), .A2(n474), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT25), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT99), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n557), .A2(n472), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n473), .A2(n556), .ZN(n479) );
  XOR2_X1 U536 ( .A(n474), .B(KEYINPUT28), .Z(n509) );
  INV_X1 U537 ( .A(n509), .ZN(n531) );
  NOR2_X1 U538 ( .A1(n500), .A2(n531), .ZN(n477) );
  INV_X1 U539 ( .A(n475), .ZN(n476) );
  NAND2_X1 U540 ( .A1(n477), .A2(n476), .ZN(n538) );
  NOR2_X1 U541 ( .A1(n540), .A2(n538), .ZN(n478) );
  NOR2_X1 U542 ( .A1(n479), .A2(n478), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n566), .A2(n548), .ZN(n481) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT83), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(n482) );
  OR2_X1 U546 ( .A1(n491), .A2(n482), .ZN(n513) );
  NOR2_X1 U547 ( .A1(n495), .A2(n513), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n488), .A2(n556), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n484), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n488), .A2(n528), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U553 ( .A1(n488), .A2(n540), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n531), .A2(n488), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n489), .B(KEYINPUT100), .ZN(n490) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  NOR2_X1 U558 ( .A1(n491), .A2(n589), .ZN(n492) );
  XNOR2_X1 U559 ( .A(n492), .B(KEYINPUT103), .ZN(n493) );
  NOR2_X1 U560 ( .A1(n594), .A2(n493), .ZN(n494) );
  XNOR2_X1 U561 ( .A(KEYINPUT37), .B(n494), .ZN(n525) );
  XNOR2_X1 U562 ( .A(KEYINPUT38), .B(n499), .ZN(n508) );
  NOR2_X1 U563 ( .A1(n500), .A2(n508), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n501) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(n501), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n504), .A2(n508), .ZN(n505) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n505), .Z(G1329GAT) );
  NOR2_X1 U569 ( .A1(n506), .A2(n508), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n292), .ZN(G1330GAT) );
  NOR2_X1 U571 ( .A1(n509), .A2(n508), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(G1331GAT) );
  INV_X1 U574 ( .A(n512), .ZN(n543) );
  NAND2_X1 U575 ( .A1(n541), .A2(n512), .ZN(n524) );
  NOR2_X1 U576 ( .A1(n524), .A2(n513), .ZN(n514) );
  XNOR2_X1 U577 ( .A(KEYINPUT106), .B(n514), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n520), .A2(n556), .ZN(n517) );
  XOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT107), .Z(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n528), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n540), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n531), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n523), .ZN(G1335GAT) );
  XOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT109), .Z(n527) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n532), .A2(n556), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n528), .A2(n532), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n540), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n536) );
  XOR2_X1 U599 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n534) );
  NAND2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n538), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n551) );
  NOR2_X1 U605 ( .A1(n541), .A2(n551), .ZN(n542) );
  XOR2_X1 U606 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  NOR2_X1 U607 ( .A1(n543), .A2(n551), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n548), .A2(n551), .ZN(n549) );
  XOR2_X1 U614 ( .A(n550), .B(n549), .Z(G1342GAT) );
  NOR2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U618 ( .A(G134GAT), .B(n555), .Z(G1343GAT) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U620 ( .A1(n537), .A2(n558), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n567), .A2(n581), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n561) );
  NAND2_X1 U625 ( .A1(n567), .A2(n512), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  XOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U629 ( .A1(n567), .A2(n589), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n581), .A2(n576), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(n573), .Z(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n512), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  NAND2_X1 U642 ( .A1(n576), .A2(n589), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT125), .B(n580), .ZN(n593) );
  INV_X1 U646 ( .A(n593), .ZN(n590) );
  NAND2_X1 U647 ( .A1(n590), .A2(n581), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  OR2_X1 U653 ( .A1(n593), .A2(n586), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U655 ( .A(G211GAT), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1354GAT) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(KEYINPUT62), .B(n595), .Z(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

