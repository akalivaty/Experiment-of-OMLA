//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n192), .A2(new_n195), .A3(new_n198), .A4(new_n193), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT81), .B(G107), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G104), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n201), .A2(new_n203), .B1(KEYINPUT3), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(G101), .B1(new_n202), .B2(G107), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n201), .B2(G104), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(G101), .ZN(new_n209));
  OR2_X1    g023(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G128), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  OAI21_X1  g032(.A(G128), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n209), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n203), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n205), .A2(KEYINPUT3), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n207), .ZN(new_n230));
  INV_X1    g044(.A(new_n205), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n227), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n202), .ZN(new_n233));
  INV_X1    g047(.A(G101), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n221), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n214), .B2(new_n219), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT82), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT10), .B1(new_n224), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT0), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n213), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n240), .A2(new_n241), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n216), .A2(new_n218), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n202), .A2(G107), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n228), .A2(new_n229), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n234), .B1(new_n206), .B2(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n230), .A2(KEYINPUT4), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n246), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n215), .A2(G146), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n210), .B2(new_n211), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n220), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n209), .A2(new_n257), .A3(KEYINPUT10), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n200), .B1(new_n239), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT86), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT86), .B(new_n200), .C1(new_n239), .C2(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT85), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n200), .B(KEYINPUT83), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n239), .A2(new_n259), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G140), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT80), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n265), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n223), .B1(new_n209), .B2(new_n222), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT82), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n266), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n258), .A3(new_n253), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT85), .A3(new_n272), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n264), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT84), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n200), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI22_X1  g099(.A1(new_n276), .A2(new_n277), .B1(new_n257), .B2(new_n209), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n200), .ZN(new_n287));
  INV_X1    g101(.A(new_n257), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n224), .A2(new_n238), .B1(new_n288), .B2(new_n235), .ZN(new_n289));
  INV_X1    g103(.A(new_n200), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n289), .A2(new_n290), .A3(new_n284), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n280), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n273), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n282), .A2(new_n293), .A3(G469), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n280), .B(new_n272), .C1(new_n287), .C2(new_n291), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n267), .B1(new_n262), .B2(new_n263), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n272), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n295), .A3(new_n296), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT95), .ZN(new_n305));
  INV_X1    g119(.A(G217), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n187), .A2(new_n306), .A3(G953), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT67), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G116), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(G122), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n308), .A2(G122), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n201), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n215), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n241), .A2(G143), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n191), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(G134), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT14), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n308), .B2(G122), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n322), .B1(new_n312), .B2(new_n324), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n314), .B(new_n321), .C1(new_n329), .C2(new_n204), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n312), .A2(new_n313), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n232), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n314), .ZN(new_n333));
  OAI21_X1  g147(.A(G134), .B1(new_n315), .B2(KEYINPUT13), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(KEYINPUT13), .B2(new_n318), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n191), .B2(new_n318), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n330), .A2(KEYINPUT94), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n328), .A2(new_n327), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n204), .B1(new_n338), .B2(new_n325), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n321), .A2(new_n314), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n339), .A2(KEYINPUT94), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n307), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT94), .B1(new_n339), .B2(new_n340), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n333), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n339), .A2(KEYINPUT94), .A3(new_n340), .ZN(new_n346));
  INV_X1    g160(.A(new_n307), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n296), .B1(new_n342), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G478), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(KEYINPUT15), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n341), .A2(new_n343), .A3(new_n344), .A4(new_n307), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n351), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n296), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(G234), .A2(G237), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(G952), .A3(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n358), .A2(G902), .A3(G953), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT21), .B(G898), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n352), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT16), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT16), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n366), .A3(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT74), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(new_n371), .A3(new_n366), .A4(G125), .ZN(new_n375));
  AND4_X1   g189(.A1(G146), .A2(new_n370), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n217), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n378), .B2(KEYINPUT75), .ZN(new_n379));
  INV_X1    g193(.A(G237), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n359), .A3(G214), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(new_n215), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G131), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n381), .A2(new_n215), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n215), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n198), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT75), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(new_n389), .A3(new_n217), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(KEYINPUT17), .A3(G131), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n379), .A2(new_n388), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n202), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n381), .B(G143), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n397), .ZN(new_n399));
  XNOR2_X1  g213(.A(G125), .B(G140), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n217), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n394), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n394), .B1(new_n392), .B2(new_n402), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT92), .B(new_n296), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G475), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n392), .A2(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(new_n394), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(G902), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT92), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n383), .A2(new_n387), .ZN(new_n414));
  INV_X1    g228(.A(new_n376), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n400), .B(KEYINPUT19), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n414), .B(new_n415), .C1(G146), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n402), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n403), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n413), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n422), .ZN(new_n424));
  AOI211_X1 g238(.A(KEYINPUT20), .B(new_n424), .C1(new_n420), .C2(new_n403), .ZN(new_n425));
  OAI22_X1  g239(.A1(new_n407), .A2(new_n412), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n305), .B1(new_n365), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G475), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n411), .B2(KEYINPUT92), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n296), .B1(new_n404), .B2(new_n405), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n421), .A2(new_n422), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT20), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(new_n413), .A3(new_n422), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n429), .A2(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n356), .B1(new_n355), .B2(new_n296), .ZN(new_n437));
  AOI211_X1 g251(.A(G902), .B(new_n351), .C1(new_n353), .C2(new_n354), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT95), .A4(new_n364), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n427), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n309), .A2(new_n311), .A3(G119), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n308), .A2(G119), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT2), .A2(G113), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT66), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT66), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT2), .A3(G113), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT2), .ZN(new_n454));
  INV_X1    g268(.A(G113), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n450), .A2(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n447), .A3(new_n445), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n458), .A2(new_n460), .B1(new_n248), .B2(new_n249), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n248), .A2(G101), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n230), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n445), .A2(KEYINPUT5), .A3(new_n447), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n455), .B1(new_n446), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT67), .B(G116), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n446), .B1(new_n467), .B2(G119), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n464), .A2(new_n466), .B1(new_n468), .B2(new_n459), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n461), .A2(new_n463), .B1(new_n209), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G122), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n444), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n461), .A2(new_n463), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n209), .A2(new_n469), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n476), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n472), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n257), .A2(new_n368), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n246), .A2(G125), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n359), .A2(G224), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT88), .B(new_n472), .C1(new_n475), .C2(new_n478), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n476), .A2(new_n477), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n471), .B1(new_n488), .B2(KEYINPUT87), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n444), .C1(KEYINPUT87), .C2(new_n488), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n481), .A2(new_n486), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n484), .A2(new_n492), .A3(new_n485), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n470), .B2(new_n471), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n485), .B1(KEYINPUT89), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(KEYINPUT89), .B2(new_n492), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n482), .A2(new_n483), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n471), .B(KEYINPUT8), .Z(new_n500));
  OR2_X1    g314(.A1(new_n209), .A2(new_n469), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n477), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n497), .A2(new_n498), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n499), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n494), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n491), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n491), .A2(new_n505), .A3(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n443), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n304), .A2(new_n441), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n306), .B1(G234), .B2(new_n296), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT22), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(G137), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n379), .A2(new_n390), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n241), .A2(G119), .ZN(new_n522));
  INV_X1    g336(.A(G119), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G128), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT24), .B(G110), .Z(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT72), .ZN(new_n528));
  INV_X1    g342(.A(G110), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n530), .A2(KEYINPUT23), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(KEYINPUT23), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n531), .A2(new_n524), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n528), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n521), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n400), .A2(new_n217), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n415), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n525), .A2(new_n526), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT76), .B(G110), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n520), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(new_n519), .C1(new_n521), .C2(new_n534), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n544), .A3(new_n296), .ZN(new_n545));
  NOR2_X1   g359(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n546), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n544), .A3(new_n296), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n516), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n542), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT78), .B1(new_n542), .B2(new_n544), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n515), .A2(G902), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n553), .B(KEYINPUT79), .Z(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n191), .A2(G137), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n194), .A2(G134), .ZN(new_n559));
  OAI21_X1  g373(.A(G131), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n199), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n257), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n200), .A2(new_n246), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT30), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n458), .A2(new_n460), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n199), .A2(new_n197), .B1(new_n242), .B2(new_n245), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n199), .A2(new_n560), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n220), .A2(new_n256), .B1(new_n567), .B2(KEYINPUT64), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n567), .A2(KEYINPUT64), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n564), .B(new_n565), .C1(new_n570), .C2(KEYINPUT30), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n380), .A2(new_n359), .A3(G210), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT27), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT26), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n576), .A2(new_n577), .A3(G101), .ZN(new_n578));
  AOI21_X1  g392(.A(G101), .B1(new_n576), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n565), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n562), .A2(new_n581), .A3(new_n563), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT31), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n567), .A2(KEYINPUT64), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n569), .A2(new_n257), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n563), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n565), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT28), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n562), .A2(new_n581), .A3(KEYINPUT28), .A4(new_n563), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n580), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT31), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n571), .A2(new_n595), .A3(new_n580), .A4(new_n582), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n584), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(G472), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT32), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(KEYINPUT32), .A3(new_n598), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT29), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n562), .A2(new_n563), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n565), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT70), .A3(new_n582), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT70), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n610), .A3(new_n565), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n606), .B(new_n590), .C1(new_n612), .C2(new_n589), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n296), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n571), .A2(new_n582), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n593), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT68), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n588), .A2(new_n580), .A3(new_n590), .A4(new_n591), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n605), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n615), .A2(KEYINPUT68), .A3(new_n593), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n614), .B1(new_n622), .B2(KEYINPUT69), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT69), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n618), .A2(new_n620), .A3(new_n624), .A4(new_n621), .ZN(new_n625));
  AOI211_X1 g439(.A(KEYINPUT71), .B(new_n604), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT71), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(KEYINPUT69), .ZN(new_n628));
  INV_X1    g442(.A(new_n614), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n630), .B2(G472), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n603), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n304), .A2(new_n441), .A3(KEYINPUT96), .A4(new_n511), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n514), .A2(new_n557), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  NAND2_X1  g449(.A1(new_n349), .A2(new_n350), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n355), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n350), .A2(G902), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n345), .B2(new_n346), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n307), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT33), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n307), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n638), .B(new_n639), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n436), .B1(new_n636), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n363), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n491), .A2(new_n505), .A3(new_n507), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n507), .B1(new_n491), .B2(new_n505), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n442), .B1(new_n510), .B2(KEYINPUT97), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n509), .A2(KEYINPUT97), .A3(new_n510), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT98), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n648), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n302), .A2(new_n295), .A3(new_n296), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n294), .A2(new_n298), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n188), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n557), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n597), .A2(new_n296), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n599), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  NAND3_X1  g485(.A1(new_n434), .A2(KEYINPUT101), .A3(new_n435), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(new_n423), .B2(new_n425), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n672), .B(new_n674), .C1(new_n437), .C2(new_n438), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n363), .B1(new_n429), .B2(new_n432), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT102), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n672), .A2(new_n674), .ZN(new_n679));
  INV_X1    g493(.A(new_n439), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n676), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n683), .A2(new_n655), .A3(new_n658), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n668), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NAND2_X1  g501(.A1(new_n547), .A2(new_n549), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n535), .A2(new_n541), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n689), .B(new_n690), .Z(new_n691));
  AOI22_X1  g505(.A1(new_n688), .A2(new_n515), .B1(new_n691), .B2(new_n554), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n667), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n514), .A2(new_n633), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  AND2_X1   g510(.A1(new_n655), .A2(new_n658), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n429), .A2(new_n432), .ZN(new_n698));
  INV_X1    g512(.A(new_n360), .ZN(new_n699));
  INV_X1    g513(.A(new_n361), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT103), .B(G900), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n663), .A2(new_n675), .A3(new_n692), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n697), .A2(new_n632), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XNOR2_X1  g521(.A(new_n703), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n304), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT40), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n509), .A2(new_n510), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT38), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n612), .A2(new_n593), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n296), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n593), .B1(new_n582), .B2(new_n571), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n601), .A2(new_n602), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n692), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n436), .A2(new_n439), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n442), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n712), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n710), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G143), .ZN(G45));
  INV_X1    g537(.A(new_n692), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n304), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n646), .A2(new_n703), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n697), .A2(new_n632), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  AND2_X1   g543(.A1(new_n632), .A2(new_n557), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n302), .A2(new_n296), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(new_n188), .A3(new_n303), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n188), .A3(new_n303), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n730), .A2(new_n660), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n632), .A2(new_n557), .A3(new_n737), .A4(new_n735), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n683), .A2(new_n655), .A3(new_n658), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n308), .ZN(G18));
  AOI21_X1  g559(.A(new_n692), .B1(new_n427), .B2(new_n440), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n632), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n655), .A2(new_n658), .A3(new_n733), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n655), .A2(new_n658), .A3(new_n750), .A4(new_n733), .ZN(new_n751));
  AOI211_X1 g565(.A(KEYINPUT107), .B(new_n747), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n751), .ZN(new_n754));
  INV_X1    g568(.A(new_n747), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n523), .ZN(G21));
  OAI21_X1  g572(.A(new_n590), .B1(new_n612), .B2(new_n589), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n593), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n584), .A3(new_n596), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n598), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT108), .B(G472), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n665), .A2(new_n763), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n557), .A2(new_n762), .A3(new_n364), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n735), .A2(new_n737), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n655), .A2(new_n658), .A3(new_n719), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  AND2_X1   g583(.A1(new_n762), .A2(new_n764), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n724), .ZN(new_n771));
  INV_X1    g585(.A(new_n726), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n749), .B2(new_n751), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n368), .ZN(G27));
  NAND3_X1  g589(.A1(new_n509), .A2(new_n442), .A3(new_n510), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n663), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n632), .A2(new_n557), .A3(new_n772), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  NOR2_X1   g595(.A1(new_n675), .A2(new_n704), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n632), .A2(new_n557), .A3(new_n782), .A4(new_n777), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT109), .B(G134), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G36));
  NAND2_X1  g599(.A1(new_n724), .A2(new_n667), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT111), .Z(new_n787));
  NAND2_X1  g601(.A1(new_n645), .A2(new_n636), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n436), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT43), .Z(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n776), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n790), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n282), .A2(new_n293), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n295), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n282), .A2(new_n293), .A3(KEYINPUT45), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n297), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT110), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n661), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n188), .A3(new_n708), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n796), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n194), .ZN(G39));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n188), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(new_n632), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n814), .A3(new_n188), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n726), .A2(new_n557), .A3(new_n776), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NOR2_X1   g632(.A1(new_n736), .A2(new_n776), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n790), .A2(new_n360), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n730), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n664), .A2(new_n717), .A3(new_n699), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT120), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n647), .ZN(new_n826));
  INV_X1    g640(.A(G952), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(G953), .ZN(new_n828));
  INV_X1    g642(.A(new_n754), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n790), .A2(new_n360), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n770), .A2(new_n557), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n822), .B(new_n828), .C1(new_n829), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n820), .A2(new_n771), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT119), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n825), .A2(new_n426), .A3(new_n788), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n712), .A2(new_n443), .A3(new_n733), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n839), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT50), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(KEYINPUT118), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n732), .A2(new_n303), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n189), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT116), .Z(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n812), .B2(new_n815), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n830), .A2(new_n831), .A3(new_n794), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT114), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n843), .B(new_n851), .C1(KEYINPUT118), .C2(new_n842), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n842), .A2(new_n835), .A3(new_n837), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n812), .A2(new_n815), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n854), .B2(new_n846), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT51), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n833), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n730), .A2(new_n684), .A3(new_n738), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n739), .A2(new_n858), .A3(new_n768), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n754), .A2(new_n755), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT107), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n754), .A2(new_n753), .A3(new_n755), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n188), .B(new_n703), .C1(new_n661), .C2(new_n662), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n718), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n655), .A3(new_n658), .A4(new_n719), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n773), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n754), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n697), .B(new_n632), .C1(new_n727), .C2(new_n705), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n778), .B(KEYINPUT42), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n646), .B1(new_n436), .B2(new_n680), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n668), .A3(new_n511), .A4(new_n364), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n634), .A2(new_n694), .A3(new_n783), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n725), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n794), .ZN(new_n880));
  INV_X1    g694(.A(new_n704), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n632), .A2(new_n439), .A3(new_n679), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n772), .A2(new_n770), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n874), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n871), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n774), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n888), .A3(new_n868), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n863), .A2(new_n873), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n742), .A2(new_n659), .B1(new_n767), .B2(new_n766), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n744), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n752), .B2(new_n756), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n634), .A2(new_n694), .A3(new_n783), .A4(new_n877), .ZN(new_n896));
  INV_X1    g710(.A(new_n884), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n780), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n873), .A4(new_n889), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  XOR2_X1   g716(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n903));
  AND3_X1   g717(.A1(new_n892), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n857), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(G952), .B2(G953), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n844), .B(KEYINPUT49), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n557), .A2(new_n188), .A3(new_n442), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n909), .A2(new_n717), .A3(new_n789), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n712), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n359), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n296), .B1(new_n892), .B2(new_n900), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n915), .B2(G210), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n481), .A2(new_n487), .A3(new_n490), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n486), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n916), .B2(new_n920), .ZN(G51));
  AND2_X1   g736(.A1(new_n915), .A2(new_n801), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n297), .B(KEYINPUT57), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n903), .B1(new_n892), .B2(new_n900), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n904), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n302), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n302), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(G54));
  NAND3_X1  g745(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  INV_X1    g746(.A(new_n421), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n913), .ZN(G60));
  NOR2_X1   g750(.A1(new_n643), .A2(new_n644), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n355), .B2(new_n637), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n905), .A2(new_n902), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT59), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n904), .A2(new_n925), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n914), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n942), .A2(new_n945), .ZN(G63));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT122), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n892), .B2(new_n900), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n913), .B1(new_n952), .B2(new_n691), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n551), .A2(new_n552), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n957), .B2(new_n952), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  OAI221_X1 g773(.A(new_n953), .B1(new_n954), .B2(new_n947), .C1(new_n957), .C2(new_n952), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  NAND4_X1  g775(.A1(new_n863), .A2(new_n634), .A3(new_n694), .A4(new_n877), .ZN(new_n962));
  NAND2_X1  g776(.A1(G224), .A2(G953), .ZN(new_n963));
  OAI22_X1  g777(.A1(new_n962), .A2(G953), .B1(new_n362), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT124), .Z(new_n965));
  INV_X1    g779(.A(G898), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n917), .B1(new_n966), .B2(G953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  MUX2_X1   g782(.A(new_n570), .B(new_n607), .S(KEYINPUT30), .Z(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(new_n417), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n887), .A2(new_n722), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n817), .A3(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n709), .A2(new_n875), .A3(new_n776), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n730), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n796), .B2(new_n808), .ZN(new_n978));
  OR3_X1    g792(.A1(new_n975), .A2(G953), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n971), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n730), .A2(new_n697), .A3(new_n719), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n783), .B1(new_n808), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n809), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n984), .A2(new_n780), .A3(new_n817), .A4(new_n887), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n359), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n270), .A2(G900), .A3(G953), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n970), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n981), .A2(new_n988), .A3(KEYINPUT125), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  OR2_X1    g809(.A1(new_n962), .A2(new_n978), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n975), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n715), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(new_n1000), .A3(new_n715), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n615), .A2(new_n580), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n995), .B1(new_n985), .B2(new_n962), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1004), .A2(KEYINPUT127), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1006), .B(new_n995), .C1(new_n985), .C2(new_n962), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1003), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n995), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n618), .A2(new_n621), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n583), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n913), .B1(new_n901), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1002), .A2(new_n1009), .A3(new_n1013), .ZN(G57));
endmodule


