

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n769), .A2(n752), .ZN(n516) );
  INV_X1 U550 ( .A(n734), .ZN(n719) );
  XNOR2_X1 U551 ( .A(n725), .B(KEYINPUT30), .ZN(n726) );
  INV_X1 U552 ( .A(n938), .ZN(n752) );
  AND2_X1 U553 ( .A1(n753), .A2(n516), .ZN(n754) );
  XNOR2_X1 U554 ( .A(G651), .B(KEYINPUT66), .ZN(n519) );
  NOR2_X1 U555 ( .A1(G651), .A2(n650), .ZN(n644) );
  NOR2_X2 U556 ( .A1(G2105), .A2(n537), .ZN(n881) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n538), .Z(n882) );
  XOR2_X1 U558 ( .A(KEYINPUT1), .B(n525), .Z(n649) );
  NOR2_X1 U559 ( .A1(G543), .A2(G651), .ZN(n634) );
  NAND2_X1 U560 ( .A1(G89), .A2(n634), .ZN(n517) );
  XOR2_X1 U561 ( .A(KEYINPUT75), .B(n517), .Z(n518) );
  XNOR2_X1 U562 ( .A(n518), .B(KEYINPUT4), .ZN(n522) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n650) );
  INV_X1 U564 ( .A(n519), .ZN(n524) );
  OR2_X1 U565 ( .A1(n650), .A2(n524), .ZN(n520) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT67), .ZN(n637) );
  NAND2_X1 U567 ( .A1(G76), .A2(n637), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(KEYINPUT5), .ZN(n531) );
  NOR2_X1 U570 ( .A1(G543), .A2(n524), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n649), .A2(G63), .ZN(n526) );
  XNOR2_X1 U572 ( .A(n526), .B(KEYINPUT76), .ZN(n528) );
  NAND2_X1 U573 ( .A1(G51), .A2(n644), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U575 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U576 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U577 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U578 ( .A(G2104), .ZN(n537) );
  NAND2_X1 U579 ( .A1(G101), .A2(n881), .ZN(n533) );
  XNOR2_X1 U580 ( .A(n533), .B(KEYINPUT23), .ZN(n534) );
  XNOR2_X1 U581 ( .A(n534), .B(KEYINPUT65), .ZN(n536) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U583 ( .A1(G113), .A2(n886), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n536), .A2(n535), .ZN(n542) );
  AND2_X1 U585 ( .A1(n537), .A2(G2105), .ZN(n885) );
  NAND2_X1 U586 ( .A1(G125), .A2(n885), .ZN(n540) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G137), .A2(n882), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U590 ( .A1(n542), .A2(n541), .ZN(G160) );
  XNOR2_X1 U591 ( .A(G168), .B(KEYINPUT8), .ZN(n543) );
  XNOR2_X1 U592 ( .A(n543), .B(KEYINPUT77), .ZN(G286) );
  XNOR2_X1 U593 ( .A(G2446), .B(KEYINPUT108), .ZN(n553) );
  XOR2_X1 U594 ( .A(G2430), .B(G2427), .Z(n545) );
  XNOR2_X1 U595 ( .A(G2435), .B(G2438), .ZN(n544) );
  XNOR2_X1 U596 ( .A(n545), .B(n544), .ZN(n549) );
  XOR2_X1 U597 ( .A(G2454), .B(KEYINPUT109), .Z(n547) );
  INV_X1 U598 ( .A(G1341), .ZN(n934) );
  XOR2_X1 U599 ( .A(G1348), .B(n934), .Z(n546) );
  XNOR2_X1 U600 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U601 ( .A(n549), .B(n548), .Z(n551) );
  XNOR2_X1 U602 ( .A(G2443), .B(G2451), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n553), .B(n552), .ZN(n554) );
  AND2_X1 U605 ( .A1(n554), .A2(G14), .ZN(G401) );
  NAND2_X1 U606 ( .A1(G52), .A2(n644), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G64), .A2(n649), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U609 ( .A1(G90), .A2(n634), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G77), .A2(n637), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U613 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U618 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(G223), .B(KEYINPUT72), .Z(n827) );
  NAND2_X1 U620 ( .A1(n827), .A2(G567), .ZN(n563) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U622 ( .A1(n634), .A2(G81), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G68), .A2(n637), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n567), .Z(n571) );
  NAND2_X1 U627 ( .A1(G56), .A2(n649), .ZN(n568) );
  XNOR2_X1 U628 ( .A(n568), .B(KEYINPUT73), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT14), .ZN(n570) );
  NOR2_X1 U630 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n644), .A2(G43), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n933) );
  INV_X1 U633 ( .A(G860), .ZN(n615) );
  OR2_X1 U634 ( .A1(n933), .A2(n615), .ZN(G153) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G54), .A2(n644), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G66), .A2(n649), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G92), .A2(n634), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G79), .A2(n637), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X2 U643 ( .A(n580), .B(KEYINPUT15), .Z(n930) );
  INV_X1 U644 ( .A(n930), .ZN(n707) );
  INV_X1 U645 ( .A(G868), .ZN(n661) );
  NAND2_X1 U646 ( .A1(n707), .A2(n661), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT74), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G53), .A2(n644), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G78), .A2(n637), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G91), .A2(n634), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G65), .A2(n649), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n927) );
  XOR2_X1 U657 ( .A(n927), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U658 ( .A1(G299), .A2(G868), .ZN(n591) );
  NOR2_X1 U659 ( .A1(G286), .A2(n661), .ZN(n590) );
  NOR2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U661 ( .A1(n615), .A2(G559), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n592), .A2(n930), .ZN(n593) );
  XNOR2_X1 U663 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U664 ( .A1(n930), .A2(G868), .ZN(n594) );
  NOR2_X1 U665 ( .A1(G559), .A2(n594), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT78), .ZN(n597) );
  NOR2_X1 U667 ( .A1(n933), .A2(G868), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U669 ( .A1(G123), .A2(n885), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G99), .A2(n881), .ZN(n599) );
  XOR2_X1 U672 ( .A(KEYINPUT79), .B(n599), .Z(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G135), .A2(n882), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G111), .A2(n886), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n988) );
  XOR2_X1 U678 ( .A(G2096), .B(n988), .Z(n606) );
  NOR2_X1 U679 ( .A1(G2100), .A2(n606), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT80), .B(n607), .Z(G156) );
  NAND2_X1 U681 ( .A1(G93), .A2(n634), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G80), .A2(n637), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G55), .A2(n644), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G67), .A2(n649), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n660) );
  NAND2_X1 U688 ( .A1(G559), .A2(n930), .ZN(n614) );
  XOR2_X1 U689 ( .A(n933), .B(n614), .Z(n658) );
  NAND2_X1 U690 ( .A1(n615), .A2(n658), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT81), .ZN(n617) );
  XOR2_X1 U692 ( .A(n660), .B(n617), .Z(G145) );
  NAND2_X1 U693 ( .A1(G50), .A2(n644), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT84), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G75), .A2(n637), .ZN(n619) );
  XOR2_X1 U696 ( .A(KEYINPUT85), .B(n619), .Z(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G88), .A2(n634), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G62), .A2(n649), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(G166) );
  INV_X1 U702 ( .A(G166), .ZN(G303) );
  NAND2_X1 U703 ( .A1(n649), .A2(G60), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n637), .A2(G72), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n634), .A2(G85), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G47), .A2(n644), .ZN(n628) );
  XOR2_X1 U708 ( .A(KEYINPUT68), .B(n628), .Z(n629) );
  NOR2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U711 ( .A(KEYINPUT69), .B(n633), .Z(G290) );
  NAND2_X1 U712 ( .A1(n644), .A2(G48), .ZN(n642) );
  NAND2_X1 U713 ( .A1(G86), .A2(n634), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G61), .A2(n649), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n637), .A2(G73), .ZN(n638) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT83), .B(n643), .Z(G305) );
  NAND2_X1 U721 ( .A1(G49), .A2(n644), .ZN(n646) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U724 ( .A(KEYINPUT82), .B(n647), .ZN(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(G288) );
  XOR2_X1 U728 ( .A(KEYINPUT19), .B(n660), .Z(n657) );
  XNOR2_X1 U729 ( .A(G299), .B(G290), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G305), .ZN(n654) );
  XOR2_X1 U731 ( .A(G303), .B(n654), .Z(n655) );
  XNOR2_X1 U732 ( .A(n655), .B(G288), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n895) );
  XNOR2_X1 U734 ( .A(n895), .B(n658), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U744 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U745 ( .A1(G219), .A2(G220), .ZN(n668) );
  XNOR2_X1 U746 ( .A(KEYINPUT22), .B(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n669), .A2(G96), .ZN(n670) );
  NOR2_X1 U748 ( .A1(G218), .A2(n670), .ZN(n671) );
  XOR2_X1 U749 ( .A(KEYINPUT86), .B(n671), .Z(n832) );
  NAND2_X1 U750 ( .A1(n832), .A2(G2106), .ZN(n675) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U752 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G108), .A2(n673), .ZN(n831) );
  NAND2_X1 U754 ( .A1(G567), .A2(n831), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n675), .A2(n674), .ZN(n833) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U757 ( .A1(n833), .A2(n676), .ZN(n830) );
  NAND2_X1 U758 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(n882), .A2(G138), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G126), .A2(n885), .ZN(n677) );
  XOR2_X1 U761 ( .A(KEYINPUT87), .B(n677), .Z(n678) );
  NAND2_X1 U762 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G102), .A2(n881), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G114), .A2(n886), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U766 ( .A1(n683), .A2(n682), .ZN(G164) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U768 ( .A(n774), .ZN(n684) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NAND2_X1 U770 ( .A1(n684), .A2(n775), .ZN(n685) );
  XNOR2_X2 U771 ( .A(n685), .B(KEYINPUT64), .ZN(n734) );
  NAND2_X1 U772 ( .A1(G2072), .A2(n719), .ZN(n686) );
  XNOR2_X1 U773 ( .A(n686), .B(KEYINPUT27), .ZN(n688) );
  INV_X1 U774 ( .A(G1956), .ZN(n926) );
  NOR2_X1 U775 ( .A1(n719), .A2(n926), .ZN(n687) );
  NOR2_X1 U776 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U777 ( .A1(n692), .A2(n927), .ZN(n691) );
  XNOR2_X1 U778 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n689), .B(KEYINPUT98), .ZN(n690) );
  XNOR2_X1 U780 ( .A(n691), .B(n690), .ZN(n715) );
  NAND2_X1 U781 ( .A1(n692), .A2(n927), .ZN(n713) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n707), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n693), .A2(n934), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n694), .A2(n734), .ZN(n695) );
  XNOR2_X1 U785 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n695), .A2(n698), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n719), .A2(G1996), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n703) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n698), .ZN(n700) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n707), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n719), .A2(n701), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U794 ( .A1(n933), .A2(n704), .ZN(n710) );
  NAND2_X1 U795 ( .A1(G2067), .A2(n719), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n734), .A2(G1348), .ZN(n705) );
  NAND2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n708) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U800 ( .A(KEYINPUT101), .B(n711), .Z(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U803 ( .A(KEYINPUT102), .B(KEYINPUT29), .Z(n716) );
  XNOR2_X1 U804 ( .A(n717), .B(n716), .ZN(n723) );
  NOR2_X1 U805 ( .A1(G1961), .A2(n719), .ZN(n718) );
  XNOR2_X1 U806 ( .A(n718), .B(KEYINPUT97), .ZN(n721) );
  XNOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .ZN(n909) );
  NAND2_X1 U808 ( .A1(n909), .A2(n719), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n727) );
  NAND2_X1 U810 ( .A1(n727), .A2(G171), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n732) );
  NAND2_X1 U812 ( .A1(n734), .A2(G8), .ZN(n769) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n769), .ZN(n745) );
  NOR2_X1 U814 ( .A1(n734), .A2(G2084), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n745), .A2(n742), .ZN(n724) );
  NAND2_X1 U816 ( .A1(G8), .A2(n724), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n726), .A2(G168), .ZN(n729) );
  NOR2_X1 U818 ( .A1(G171), .A2(n727), .ZN(n728) );
  NOR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n730), .Z(n731) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U822 ( .A1(n743), .A2(G286), .ZN(n739) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n769), .ZN(n733) );
  XOR2_X1 U824 ( .A(KEYINPUT103), .B(n733), .Z(n736) );
  NOR2_X1 U825 ( .A1(n734), .A2(G2090), .ZN(n735) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U827 ( .A1(G303), .A2(n737), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U830 ( .A(n741), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U831 ( .A1(G8), .A2(n742), .ZN(n747) );
  INV_X1 U832 ( .A(n743), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n762) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n755), .A2(n750), .ZN(n937) );
  NAND2_X1 U839 ( .A1(n762), .A2(n937), .ZN(n753) );
  NAND2_X1 U840 ( .A1(G288), .A2(G1976), .ZN(n751) );
  XNOR2_X1 U841 ( .A(n751), .B(KEYINPUT104), .ZN(n938) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n754), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n756), .A2(n769), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n944) );
  NAND2_X1 U847 ( .A1(n759), .A2(n944), .ZN(n773) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U849 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n769), .A2(n763), .ZN(n764) );
  XNOR2_X1 U852 ( .A(n764), .B(KEYINPUT105), .ZN(n771) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XNOR2_X1 U854 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n765) );
  XNOR2_X1 U855 ( .A(n765), .B(KEYINPUT95), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n767), .B(n766), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n787) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n822) );
  XNOR2_X1 U861 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  XNOR2_X1 U862 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G128), .A2(n885), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G116), .A2(n886), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n779), .B(n778), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n882), .A2(G140), .ZN(n780) );
  XNOR2_X1 U868 ( .A(n780), .B(KEYINPUT88), .ZN(n782) );
  NAND2_X1 U869 ( .A1(G104), .A2(n881), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n783), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n786), .ZN(n878) );
  NOR2_X1 U874 ( .A1(n811), .A2(n878), .ZN(n987) );
  NAND2_X1 U875 ( .A1(n822), .A2(n987), .ZN(n818) );
  AND2_X1 U876 ( .A1(n787), .A2(n818), .ZN(n810) );
  XOR2_X1 U877 ( .A(KEYINPUT91), .B(G1991), .Z(n915) );
  NAND2_X1 U878 ( .A1(G119), .A2(n885), .ZN(n789) );
  NAND2_X1 U879 ( .A1(G95), .A2(n881), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n886), .A2(G107), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT90), .B(n790), .Z(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n882), .A2(G131), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n863) );
  NAND2_X1 U886 ( .A1(n915), .A2(n863), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G105), .A2(n881), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT38), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G141), .A2(n882), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G117), .A2(n886), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n885), .A2(G129), .ZN(n798) );
  XOR2_X1 U893 ( .A(KEYINPUT92), .B(n798), .Z(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n874) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n874), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U898 ( .A(KEYINPUT93), .B(n805), .ZN(n984) );
  INV_X1 U899 ( .A(n822), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n984), .A2(n806), .ZN(n814) );
  XNOR2_X1 U901 ( .A(KEYINPUT94), .B(n814), .ZN(n808) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n936) );
  AND2_X1 U903 ( .A1(n936), .A2(n822), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n825) );
  NAND2_X1 U906 ( .A1(n811), .A2(n878), .ZN(n1007) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n874), .ZN(n994) );
  NOR2_X1 U908 ( .A1(n915), .A2(n863), .ZN(n989) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n989), .A2(n812), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n994), .A2(n815), .ZN(n816) );
  XNOR2_X1 U913 ( .A(KEYINPUT106), .B(n816), .ZN(n817) );
  XNOR2_X1 U914 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n1007), .A2(n820), .ZN(n821) );
  XOR2_X1 U917 ( .A(KEYINPUT107), .B(n821), .Z(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT40), .B(n826), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(KEYINPUT110), .B(n833), .Z(G319) );
  XOR2_X1 U933 ( .A(KEYINPUT42), .B(G2090), .Z(n835) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2072), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U936 ( .A(n836), .B(G2100), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2084), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n840) );
  XNOR2_X1 U940 ( .A(KEYINPUT111), .B(G2678), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(G227) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1971), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1976), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n845), .B(KEYINPUT112), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n926), .B(G1961), .ZN(n849) );
  XNOR2_X1 U950 ( .A(G1981), .B(G1966), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U952 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U953 ( .A(KEYINPUT113), .B(G2474), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n885), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT114), .ZN(n855) );
  XNOR2_X1 U957 ( .A(KEYINPUT44), .B(n855), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G112), .A2(n886), .ZN(n856) );
  XOR2_X1 U959 ( .A(KEYINPUT115), .B(n856), .Z(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G100), .A2(n881), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G136), .A2(n882), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U964 ( .A1(n862), .A2(n861), .ZN(G162) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n863), .B(n988), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U968 ( .A(G160), .B(n866), .Z(n877) );
  NAND2_X1 U969 ( .A1(G130), .A2(n885), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G118), .A2(n886), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G106), .A2(n881), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G142), .A2(n882), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U975 ( .A(n871), .B(KEYINPUT45), .Z(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n878), .B(G162), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n893) );
  NAND2_X1 U981 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U984 ( .A1(G127), .A2(n885), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G115), .A2(n886), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n998) );
  XOR2_X1 U989 ( .A(n998), .B(G164), .Z(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U991 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n933), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n930), .B(G171), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G37), .A2(n899), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n900) );
  XOR2_X1 U998 ( .A(KEYINPUT49), .B(n900), .Z(n901) );
  NAND2_X1 U999 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n902), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n903), .B(KEYINPUT116), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1006 ( .A(G2067), .B(G26), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(G33), .B(G2072), .ZN(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n914) );
  XOR2_X1 U1009 ( .A(G1996), .B(G32), .Z(n908) );
  NAND2_X1 U1010 ( .A1(n908), .A2(G28), .ZN(n912) );
  XOR2_X1 U1011 ( .A(G27), .B(n909), .Z(n910) );
  XNOR2_X1 U1012 ( .A(KEYINPUT122), .B(n910), .ZN(n911) );
  NOR2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(G25), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1017 ( .A(KEYINPUT53), .B(n918), .Z(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT54), .B(G34), .Z(n919) );
  XNOR2_X1 U1019 ( .A(G2084), .B(n919), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(G35), .B(G2090), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1023 ( .A(KEYINPUT55), .B(n924), .Z(n925) );
  NOR2_X1 U1024 ( .A1(G29), .A2(n925), .ZN(n981) );
  INV_X1 U1025 ( .A(G16), .ZN(n977) );
  XOR2_X1 U1026 ( .A(n977), .B(KEYINPUT56), .Z(n953) );
  XOR2_X1 U1027 ( .A(n927), .B(n926), .Z(n929) );
  XOR2_X1 U1028 ( .A(G301), .B(G1961), .Z(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1030 ( .A(G1348), .B(n930), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n951) );
  XOR2_X1 U1032 ( .A(n934), .B(n933), .Z(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n943) );
  AND2_X1 U1034 ( .A1(G303), .A2(G1971), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(KEYINPUT124), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G168), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(n946), .B(KEYINPUT57), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT123), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n979) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G21), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G5), .B(G1961), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n966) );
  XOR2_X1 U1049 ( .A(G1341), .B(G19), .Z(n957) );
  XOR2_X1 U1050 ( .A(G1956), .B(G20), .Z(n956) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n963) );
  XOR2_X1 U1052 ( .A(G1981), .B(G6), .Z(n961) );
  XOR2_X1 U1053 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n958) );
  XNOR2_X1 U1054 ( .A(G4), .B(n958), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n959), .B(G1348), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT60), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n973) );
  XNOR2_X1 U1060 ( .A(G1976), .B(G23), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G1971), .B(G22), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n970) );
  XOR2_X1 U1063 ( .A(G1986), .B(G24), .Z(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT58), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT61), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT126), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n982), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n983), .B(KEYINPUT127), .ZN(n1014) );
  XNOR2_X1 U1074 ( .A(G160), .B(G2084), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n991) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(KEYINPUT117), .B(n992), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1082 ( .A(KEYINPUT51), .B(n995), .Z(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1005) );
  XNOR2_X1 U1084 ( .A(G164), .B(G2078), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G2072), .B(n998), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(n999), .B(KEYINPUT118), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(n1002), .B(KEYINPUT50), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT119), .B(n1003), .Z(n1004) );
  NOR2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(n1008), .B(KEYINPUT52), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(n1009), .B(KEYINPUT120), .ZN(n1010) );
  NOR2_X1 U1094 ( .A1(KEYINPUT55), .A2(n1010), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT121), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1096 ( .A1(n1012), .A2(G29), .ZN(n1013) );
  NAND2_X1 U1097 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1015), .ZN(G150) );
  INV_X1 U1099 ( .A(G150), .ZN(G311) );
endmodule

