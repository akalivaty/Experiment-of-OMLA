//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT71), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n201), .B2(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT70), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT24), .B(G110), .Z(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n197), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n196), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G125), .B(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n194), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n213), .B1(new_n210), .B2(new_n212), .ZN(new_n220));
  INV_X1    g034(.A(G110), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(new_n199), .C1(new_n202), .C2(new_n204), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n219), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n215), .B1(new_n217), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n226), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n215), .B(new_n229), .C1(new_n217), .C2(new_n224), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT73), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G217), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(G234), .B2(new_n232), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n236), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n232), .A4(new_n233), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT73), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n231), .A2(new_n233), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n239), .A2(G902), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n240), .A2(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n248), .A2(G134), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(G134), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n253));
  OAI211_X1 g067(.A(G134), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n248), .A2(G134), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(KEYINPUT66), .A3(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT64), .A2(G143), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(G146), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n266), .A2(G146), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT64), .A2(G143), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT64), .A2(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n194), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n194), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT1), .B1(new_n266), .B2(G146), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n276), .A2(new_n278), .B1(G128), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n256), .B(new_n264), .C1(new_n273), .C2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n251), .A2(new_n255), .A3(new_n254), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n255), .B1(new_n251), .B2(new_n254), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n269), .A2(new_n271), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT64), .B(G143), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n277), .B1(new_n287), .B2(new_n194), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT0), .B(G128), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n281), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n269), .A2(new_n271), .A3(new_n285), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n289), .B1(new_n276), .B2(new_n278), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n253), .ZN(new_n298));
  NAND2_X1  g112(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n261), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n257), .B2(G137), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n258), .ZN(new_n302));
  OAI21_X1  g116(.A(G131), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n256), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n286), .B(KEYINPUT67), .C1(new_n288), .C2(new_n289), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n297), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT30), .A3(new_n281), .ZN(new_n307));
  XNOR2_X1  g121(.A(G116), .B(G119), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT2), .B(G113), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n310), .A3(new_n281), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G237), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n227), .A3(G210), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT27), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT26), .B(G101), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n313), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n291), .A2(new_n311), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n306), .A2(KEYINPUT28), .A3(new_n310), .A4(new_n281), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n319), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n314), .B2(new_n320), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT68), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n306), .A2(new_n281), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n311), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT69), .A3(new_n313), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n336), .A3(new_n311), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(KEYINPUT28), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n338), .A2(KEYINPUT29), .A3(new_n319), .A4(new_n324), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n330), .A2(new_n232), .A3(new_n332), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G472), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n312), .A2(new_n319), .A3(new_n313), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT31), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n320), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n312), .A2(new_n346), .A3(new_n319), .A4(new_n313), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n247), .B1(new_n341), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G478), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT15), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  INV_X1    g172(.A(G122), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G116), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n360), .B2(KEYINPUT14), .ZN(new_n361));
  XNOR2_X1  g175(.A(G116), .B(G122), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT88), .B1(new_n287), .B2(new_n198), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n274), .A2(new_n275), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G128), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n198), .A2(G143), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n257), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n257), .B1(new_n368), .B2(new_n369), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n368), .A2(KEYINPUT89), .A3(new_n257), .A4(new_n369), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n362), .B(G107), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n368), .A2(new_n380), .B1(new_n198), .B2(G143), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n364), .A2(new_n367), .A3(KEYINPUT13), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n257), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n373), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n385), .A2(new_n238), .A3(G953), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n373), .B(new_n386), .C1(new_n379), .C2(new_n383), .ZN(new_n389));
  AOI21_X1  g203(.A(G902), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT90), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT90), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n357), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n368), .A2(new_n380), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n382), .A3(new_n369), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G134), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n377), .B1(new_n370), .B2(new_n374), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n376), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n386), .B1(new_n401), .B2(new_n373), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n393), .B(new_n232), .C1(new_n396), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n357), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(G234), .A2(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(G952), .A3(new_n227), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT21), .B(G898), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT92), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(G902), .A3(G953), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n395), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  INV_X1    g229(.A(G104), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n196), .B(KEYINPUT72), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n315), .A2(new_n227), .A3(G143), .A4(G214), .ZN(new_n419));
  INV_X1    g233(.A(G214), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n420), .A2(G237), .A3(G953), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n287), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G131), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n255), .B(new_n419), .C1(new_n287), .C2(new_n421), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n218), .B(KEYINPUT19), .Z(new_n426));
  OAI211_X1 g240(.A(new_n418), .B(new_n425), .C1(G146), .C2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n218), .B(new_n194), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n255), .ZN(new_n430));
  OAI221_X1 g244(.A(new_n428), .B1(new_n422), .B2(new_n430), .C1(new_n423), .C2(new_n429), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n417), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(KEYINPUT17), .A3(G131), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(KEYINPUT85), .A3(new_n195), .A4(new_n196), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n423), .A2(new_n435), .A3(new_n424), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n191), .A2(G146), .A3(new_n192), .ZN(new_n438));
  AOI21_X1  g252(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT85), .B1(new_n440), .B2(new_n433), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n417), .B(new_n431), .C1(new_n437), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n422), .A2(KEYINPUT17), .A3(G131), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n197), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n436), .A3(new_n434), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n448), .A2(KEYINPUT86), .A3(new_n417), .A4(new_n431), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n432), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G475), .A2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT20), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OR3_X1    g269(.A1(new_n450), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT87), .B(KEYINPUT20), .C1(new_n450), .C2(new_n452), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n417), .B1(new_n448), .B2(new_n431), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n444), .B2(new_n449), .ZN(new_n460));
  OAI21_X1  g274(.A(G475), .B1(new_n460), .B2(G902), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n414), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT3), .B1(new_n416), .B2(G107), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n358), .A3(G104), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n416), .A2(G107), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(G101), .ZN(new_n470));
  INV_X1    g284(.A(G101), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n467), .A3(new_n471), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT4), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT75), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(G101), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT75), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT4), .A4(new_n472), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT4), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n469), .A2(new_n479), .A3(G101), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT76), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT76), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n469), .A2(new_n482), .A3(new_n479), .A4(G101), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n310), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n309), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n308), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT5), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n201), .A3(G116), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G113), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n487), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n358), .A2(KEYINPUT77), .A3(G104), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT77), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n416), .B2(G107), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n358), .A2(G104), .ZN(new_n496));
  OAI211_X1 g310(.A(G101), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n472), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n485), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT80), .ZN(new_n502));
  XNOR2_X1  g316(.A(G110), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT79), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n499), .B1(new_n478), .B2(new_n484), .ZN(new_n506));
  INV_X1    g320(.A(new_n504), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT80), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n501), .A2(new_n509), .A3(new_n504), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT81), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n290), .A2(G125), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n276), .A2(new_n278), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n279), .A2(G128), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n189), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n227), .A2(G224), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT82), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n520), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT81), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n501), .A2(new_n524), .A3(new_n509), .A4(new_n504), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n511), .A2(new_n513), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n504), .A2(KEYINPUT8), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n504), .A2(KEYINPUT8), .ZN(new_n528));
  INV_X1    g342(.A(new_n498), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n492), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT83), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n488), .B1(new_n531), .B2(new_n491), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n490), .A2(KEYINPUT83), .A3(G113), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n498), .B1(new_n534), .B2(new_n487), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT7), .B(new_n521), .C1(new_n520), .C2(KEYINPUT84), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n514), .A2(new_n519), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n506), .A2(new_n507), .ZN(new_n542));
  AOI21_X1  g356(.A(G902), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G210), .B1(G237), .B2(G902), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n526), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n526), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n464), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT74), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G110), .B(G140), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n227), .A2(G227), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n269), .A2(new_n271), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT1), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n287), .B2(new_n194), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n557), .B2(new_n198), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n498), .B1(new_n558), .B2(new_n518), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n517), .A2(new_n498), .A3(new_n518), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n304), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT12), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT12), .B(new_n304), .C1(new_n559), .C2(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n558), .A2(new_n518), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n529), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n517), .B2(new_n518), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n567), .A2(new_n568), .B1(new_n529), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n304), .B(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n481), .A2(new_n483), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n478), .A2(new_n297), .A3(new_n305), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n554), .B1(new_n565), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n478), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n572), .A2(new_n297), .A3(new_n305), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n569), .A2(new_n529), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n559), .B2(KEYINPUT10), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n304), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n574), .A3(new_n554), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(G469), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(G469), .A2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n284), .B1(new_n570), .B2(new_n573), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n553), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n565), .A2(new_n574), .A3(new_n554), .ZN(new_n590));
  AOI211_X1 g404(.A(G469), .B(G902), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n550), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n547), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n355), .A2(new_n463), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n348), .B2(new_n232), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n349), .B2(new_n348), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n574), .A2(new_n554), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n588), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n575), .ZN(new_n601));
  OAI21_X1  g415(.A(G469), .B1(new_n601), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n590), .ZN(new_n603));
  INV_X1    g417(.A(G469), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n232), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n549), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n606), .A3(new_n246), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT93), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n598), .A2(new_n606), .A3(new_n609), .A4(new_n246), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT94), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n396), .B2(new_n402), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n388), .A2(new_n614), .A3(new_n389), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(G478), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n356), .A2(new_n232), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n390), .B2(new_n356), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n462), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n464), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n526), .A2(new_n543), .ZN(new_n623));
  INV_X1    g437(.A(new_n544), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n526), .A2(new_n543), .A3(new_n544), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n413), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n612), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT34), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AND3_X1   g445(.A1(new_n455), .A2(KEYINPUT95), .A3(new_n457), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT95), .B1(new_n455), .B2(new_n457), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n456), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n461), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n395), .B2(new_n407), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n413), .B(KEYINPUT96), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n634), .A2(new_n640), .A3(new_n636), .A4(new_n637), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n627), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n612), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n358), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n229), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(new_n225), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n245), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n241), .A2(KEYINPUT73), .A3(new_n242), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n237), .A2(new_n239), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(new_n598), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n593), .A3(new_n463), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n627), .A2(new_n606), .ZN(new_n665));
  AOI22_X1  g479(.A1(G472), .A2(new_n340), .B1(new_n351), .B2(new_n353), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n665), .A2(new_n666), .A3(new_n658), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n412), .A2(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n409), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n634), .A2(new_n636), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n670), .A3(KEYINPUT102), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n341), .A2(new_n354), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n593), .A2(new_n673), .A3(new_n659), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n634), .A2(new_n636), .A3(new_n669), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT103), .B(G128), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G30));
  XNOR2_X1  g493(.A(new_n669), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n606), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n240), .A2(new_n243), .B1(new_n245), .B2(new_n650), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n682), .A2(new_n464), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n545), .A2(new_n546), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n314), .A2(new_n319), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n335), .A2(new_n337), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n232), .B(new_n688), .C1(new_n689), .C2(new_n319), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G472), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n354), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n395), .A2(new_n407), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n462), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n685), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n365), .ZN(G45));
  INV_X1    g510(.A(new_n669), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n619), .C1(new_n458), .C2(new_n461), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n674), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n194), .ZN(G48));
  INV_X1    g515(.A(new_n590), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n554), .B1(new_n582), .B2(new_n574), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n232), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n548), .A3(new_n605), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n708), .A3(new_n548), .A4(new_n605), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n628), .ZN(new_n711));
  INV_X1    g525(.A(new_n621), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n355), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND2_X1  g529(.A1(new_n339), .A2(new_n232), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT68), .B1(new_n331), .B2(new_n327), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n596), .B1(new_n718), .B2(new_n332), .ZN(new_n719));
  INV_X1    g533(.A(new_n353), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n352), .B1(new_n348), .B2(new_n349), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n246), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n707), .A2(new_n709), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n639), .A2(new_n725), .A3(new_n627), .A4(new_n641), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  AOI21_X1  g541(.A(new_n658), .B1(new_n354), .B2(new_n341), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n710), .A2(new_n728), .A3(new_n627), .A4(new_n463), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AND2_X1   g544(.A1(new_n458), .A2(new_n461), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n406), .B1(new_n405), .B2(new_n391), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n394), .A2(new_n357), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n731), .A2(new_n547), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n348), .A2(new_n232), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G472), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n319), .B1(new_n338), .B2(new_n324), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n343), .A2(new_n347), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n349), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(new_n740), .A3(new_n246), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n737), .A2(new_n740), .A3(new_n743), .A4(new_n246), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n710), .A2(new_n735), .A3(new_n745), .A4(new_n637), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  INV_X1    g561(.A(new_n349), .ZN(new_n748));
  INV_X1    g562(.A(new_n739), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n338), .A2(new_n324), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n320), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n683), .A3(new_n597), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n707), .A2(new_n753), .A3(new_n627), .A4(new_n709), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n699), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n189), .ZN(G27));
  NAND3_X1  g570(.A1(new_n625), .A2(new_n464), .A3(new_n626), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n548), .B1(new_n586), .B2(new_n591), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n355), .A2(new_n698), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n355), .A2(new_n698), .A3(KEYINPUT106), .A4(new_n759), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n355), .A2(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n355), .A2(KEYINPUT107), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n698), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n255), .ZN(G33));
  NOR4_X1   g585(.A1(new_n675), .A2(new_n723), .A3(new_n758), .A4(new_n757), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT108), .B(G134), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G36));
  OR2_X1    g588(.A1(new_n462), .A2(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n731), .A2(new_n620), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n777), .B1(new_n462), .B2(KEYINPUT109), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n731), .A3(new_n620), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n598), .B(new_n683), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT44), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n545), .A2(new_n546), .A3(new_n622), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n780), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n598), .A2(new_n683), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n601), .A2(KEYINPUT45), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n600), .B2(new_n575), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(G469), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n585), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n591), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n548), .A3(new_n680), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n782), .A2(new_n783), .A3(new_n788), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  NOR4_X1   g613(.A1(new_n699), .A2(new_n673), .A3(new_n246), .A4(new_n757), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n796), .A2(KEYINPUT47), .A3(new_n548), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT47), .B1(new_n796), .B2(new_n548), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT110), .B(G140), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G42));
  AOI21_X1  g619(.A(new_n409), .B1(new_n742), .B2(new_n744), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n784), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n687), .A2(new_n710), .A3(new_n622), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n801), .A2(new_n802), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n705), .A2(new_n549), .A3(new_n605), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n807), .A2(new_n757), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n710), .A2(new_n783), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n409), .B1(new_n819), .B2(KEYINPUT116), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n354), .A2(new_n246), .A3(new_n691), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n731), .A3(new_n619), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n753), .A3(new_n784), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(KEYINPUT117), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n812), .B(new_n818), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n814), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n815), .B(KEYINPUT115), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n817), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n826), .A3(new_n825), .ZN(new_n833));
  INV_X1    g647(.A(new_n812), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n813), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n820), .A2(new_n821), .A3(new_n712), .A4(new_n824), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(G952), .A3(new_n227), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n820), .A2(new_n784), .A3(new_n821), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n766), .A2(new_n767), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n838), .A2(KEYINPUT48), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT48), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n807), .A2(new_n547), .A3(new_n724), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT118), .Z(new_n844));
  AND3_X1   g658(.A1(new_n842), .A2(new_n844), .A3(KEYINPUT119), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT119), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n829), .B(new_n835), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n627), .A2(new_n639), .A3(new_n641), .A4(new_n725), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n746), .A2(new_n729), .A3(new_n713), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n729), .A2(new_n713), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n726), .A4(new_n746), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n772), .B1(new_n765), .B2(new_n769), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n621), .B1(new_n462), .B2(new_n734), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n627), .A2(new_n637), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n608), .A2(new_n856), .A3(new_n610), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n635), .A2(new_n697), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n783), .A2(new_n734), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n456), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n455), .A2(new_n457), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT95), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n455), .A2(KEYINPUT95), .A3(new_n457), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT113), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n395), .A2(new_n860), .A3(new_n407), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n757), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n634), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n872), .A3(new_n606), .A4(new_n728), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n593), .B(new_n463), .C1(new_n660), .C2(new_n355), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n698), .A2(new_n759), .A3(new_n753), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n859), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n851), .A2(new_n854), .A3(new_n855), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n699), .B1(new_n674), .B2(new_n754), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n671), .B2(new_n676), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n758), .A2(new_n654), .A3(new_n697), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n735), .A2(new_n880), .A3(new_n692), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n877), .B(new_n886), .C1(new_n887), .C2(KEYINPUT53), .ZN(new_n888));
  INV_X1    g702(.A(new_n878), .ZN(new_n889));
  AND4_X1   g703(.A1(KEYINPUT52), .A2(new_n677), .A3(new_n889), .A4(new_n881), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(new_n879), .B2(new_n881), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n851), .A2(new_n854), .A3(new_n876), .A4(new_n855), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n848), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n876), .A2(new_n855), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n849), .A2(new_n850), .A3(new_n893), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n898), .A2(new_n848), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n847), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(G952), .A2(G953), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT120), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n776), .A2(new_n247), .A3(new_n549), .A4(new_n622), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT111), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n705), .A2(new_n605), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT49), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n692), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n687), .A3(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n903), .A2(new_n905), .B1(new_n908), .B2(new_n913), .ZN(G75));
  AOI21_X1  g728(.A(new_n232), .B1(new_n898), .B2(new_n901), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n511), .A2(new_n513), .A3(new_n525), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n523), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT55), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(KEYINPUT56), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n916), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n916), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n227), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  INV_X1    g740(.A(new_n792), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n585), .B(KEYINPUT57), .Z(new_n931));
  AOI21_X1  g745(.A(new_n848), .B1(new_n898), .B2(new_n901), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n902), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n603), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n925), .B1(new_n930), .B2(new_n934), .ZN(G54));
  NAND3_X1  g749(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n450), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n450), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n925), .ZN(G60));
  XNOR2_X1  g753(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n617), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n897), .B2(new_n902), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n613), .A2(new_n615), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  INV_X1    g760(.A(new_n944), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n941), .C1(new_n902), .C2(new_n932), .ZN(new_n948));
  INV_X1    g762(.A(new_n925), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n898), .B2(new_n901), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n650), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n955), .B(new_n949), .C1(new_n244), .C2(new_n954), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G66));
  AOI21_X1  g772(.A(new_n227), .B1(new_n411), .B2(G224), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n851), .A2(new_n854), .A3(new_n859), .A4(new_n874), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n959), .B1(new_n964), .B2(new_n227), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n917), .B1(G898), .B2(new_n227), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n965), .B(new_n966), .Z(G69));
  NAND4_X1  g781(.A1(new_n796), .A2(new_n548), .A3(new_n680), .A4(new_n735), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n839), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n970), .A2(new_n798), .A3(new_n803), .A4(new_n879), .ZN(new_n971));
  INV_X1    g785(.A(new_n855), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n227), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n293), .A2(new_n307), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n426), .ZN(new_n976));
  NAND2_X1  g790(.A1(G900), .A2(G953), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n681), .A2(new_n757), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n856), .A2(new_n979), .A3(new_n355), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n797), .B(new_n783), .C1(new_n781), .C2(KEYINPUT44), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n786), .A2(new_n787), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n803), .B(new_n980), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n879), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n984), .A2(KEYINPUT62), .A3(new_n695), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  INV_X1    g800(.A(new_n695), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n879), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(G953), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n978), .B1(new_n990), .B2(new_n976), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n227), .B1(G227), .B2(G900), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n992), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n978), .B(new_n994), .C1(new_n990), .C2(new_n976), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(G72));
  NAND3_X1  g810(.A1(new_n973), .A2(new_n963), .A3(new_n962), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n314), .A2(new_n319), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n888), .A2(new_n896), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n321), .A2(new_n342), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n999), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1002), .B(new_n949), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n989), .A2(new_n963), .A3(new_n962), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n688), .B1(new_n1007), .B2(new_n999), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT127), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1006), .A2(new_n1009), .ZN(G57));
endmodule


