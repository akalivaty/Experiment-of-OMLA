

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  NOR2_X1 U322 ( .A1(n553), .A2(n476), .ZN(n586) );
  XNOR2_X1 U323 ( .A(n464), .B(KEYINPUT48), .ZN(n555) );
  XNOR2_X1 U324 ( .A(n310), .B(n309), .ZN(n454) );
  XOR2_X1 U325 ( .A(KEYINPUT73), .B(n335), .Z(n381) );
  XNOR2_X1 U326 ( .A(n367), .B(n290), .ZN(n370) );
  XNOR2_X1 U327 ( .A(KEYINPUT37), .B(KEYINPUT101), .ZN(n445) );
  XNOR2_X1 U328 ( .A(n381), .B(n380), .ZN(n386) );
  XOR2_X1 U329 ( .A(n339), .B(n338), .Z(n566) );
  XOR2_X1 U330 ( .A(n324), .B(n336), .Z(n578) );
  XOR2_X1 U331 ( .A(n366), .B(n365), .Z(n290) );
  XOR2_X1 U332 ( .A(n381), .B(n336), .Z(n291) );
  XNOR2_X1 U333 ( .A(G190GAT), .B(G218GAT), .ZN(n332) );
  XNOR2_X1 U334 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n460) );
  XNOR2_X1 U335 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U336 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U337 ( .A(n437), .B(n364), .ZN(n309) );
  XNOR2_X1 U338 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U339 ( .A(KEYINPUT36), .B(n547), .Z(n471) );
  XOR2_X1 U340 ( .A(KEYINPUT74), .B(n566), .Z(n547) );
  XNOR2_X1 U341 ( .A(n447), .B(KEYINPUT107), .ZN(n534) );
  XNOR2_X1 U342 ( .A(n388), .B(n376), .ZN(n538) );
  XNOR2_X1 U343 ( .A(n483), .B(n482), .ZN(n511) );
  XNOR2_X1 U344 ( .A(n472), .B(G218GAT), .ZN(n473) );
  XNOR2_X1 U345 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n479) );
  XNOR2_X1 U346 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U347 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U348 ( .A(n474), .B(n473), .ZN(G1355GAT) );
  XNOR2_X1 U349 ( .A(n480), .B(n479), .ZN(G1351GAT) );
  XNOR2_X1 U350 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G106GAT), .Z(n293) );
  XNOR2_X1 U352 ( .A(G85GAT), .B(KEYINPUT69), .ZN(n292) );
  XNOR2_X1 U353 ( .A(n293), .B(n292), .ZN(n330) );
  XNOR2_X1 U354 ( .A(n330), .B(KEYINPUT32), .ZN(n297) );
  INV_X1 U355 ( .A(n297), .ZN(n295) );
  AND2_X1 U356 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  INV_X1 U357 ( .A(n296), .ZN(n294) );
  NAND2_X1 U358 ( .A1(n295), .A2(n294), .ZN(n299) );
  NAND2_X1 U359 ( .A1(n297), .A2(n296), .ZN(n298) );
  NAND2_X1 U360 ( .A1(n299), .A2(n298), .ZN(n303) );
  XOR2_X1 U361 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n301) );
  XNOR2_X1 U362 ( .A(G92GAT), .B(KEYINPUT31), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U365 ( .A(KEYINPUT71), .B(G204GAT), .Z(n305) );
  XNOR2_X1 U366 ( .A(G64GAT), .B(G176GAT), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n382) );
  XNOR2_X1 U368 ( .A(G148GAT), .B(G78GAT), .ZN(n306) );
  XNOR2_X1 U369 ( .A(n306), .B(KEYINPUT68), .ZN(n355) );
  XOR2_X1 U370 ( .A(n382), .B(n355), .Z(n307) );
  XNOR2_X1 U371 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U372 ( .A(G57GAT), .B(KEYINPUT13), .Z(n437) );
  XNOR2_X1 U373 ( .A(G120GAT), .B(G71GAT), .ZN(n364) );
  XOR2_X1 U374 ( .A(KEYINPUT41), .B(n454), .Z(n572) );
  INV_X1 U375 ( .A(n572), .ZN(n559) );
  XOR2_X1 U376 ( .A(G8GAT), .B(G169GAT), .Z(n379) );
  XOR2_X1 U377 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n312) );
  XNOR2_X1 U378 ( .A(G15GAT), .B(G197GAT), .ZN(n311) );
  XNOR2_X1 U379 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n379), .B(n313), .ZN(n317) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n345) );
  XOR2_X1 U382 ( .A(KEYINPUT29), .B(n345), .Z(n315) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U384 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U385 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U386 ( .A(n318), .B(G50GAT), .Z(n320) );
  XOR2_X1 U387 ( .A(G113GAT), .B(G1GAT), .Z(n401) );
  XNOR2_X1 U388 ( .A(n401), .B(G36GAT), .ZN(n319) );
  XNOR2_X1 U389 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U390 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n322) );
  XNOR2_X1 U391 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n321) );
  XNOR2_X1 U392 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(n323), .ZN(n336) );
  NOR2_X1 U394 ( .A1(n559), .A2(n578), .ZN(n515) );
  XNOR2_X1 U395 ( .A(G162GAT), .B(G50GAT), .ZN(n325) );
  XNOR2_X1 U396 ( .A(n325), .B(KEYINPUT72), .ZN(n356) );
  XOR2_X1 U397 ( .A(n356), .B(G134GAT), .Z(n327) );
  NAND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U399 ( .A(n327), .B(n326), .ZN(n339) );
  XOR2_X1 U400 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n329) );
  XNOR2_X1 U401 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n328) );
  XNOR2_X1 U402 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U403 ( .A(n331), .B(n330), .Z(n337) );
  INV_X1 U404 ( .A(n332), .ZN(n334) );
  XNOR2_X1 U405 ( .A(G92GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U406 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U407 ( .A(n337), .B(n291), .ZN(n338) );
  XOR2_X1 U408 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n341) );
  XNOR2_X1 U409 ( .A(KEYINPUT84), .B(G197GAT), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U411 ( .A(G211GAT), .B(n342), .Z(n387) );
  XOR2_X1 U412 ( .A(G155GAT), .B(KEYINPUT2), .Z(n344) );
  XNOR2_X1 U413 ( .A(KEYINPUT86), .B(KEYINPUT3), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n409) );
  XOR2_X1 U415 ( .A(n409), .B(n345), .Z(n347) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U417 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n387), .B(n348), .ZN(n360) );
  XOR2_X1 U419 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n350) );
  XNOR2_X1 U420 ( .A(G218GAT), .B(G106GAT), .ZN(n349) );
  XNOR2_X1 U421 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U422 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n352) );
  XNOR2_X1 U423 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U425 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U426 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n360), .B(n359), .ZN(n475) );
  XOR2_X1 U429 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n362) );
  XNOR2_X1 U430 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U432 ( .A(G183GAT), .B(n363), .Z(n388) );
  XNOR2_X1 U433 ( .A(n364), .B(G99GAT), .ZN(n367) );
  XOR2_X1 U434 ( .A(G15GAT), .B(G169GAT), .Z(n366) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(G134GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n368), .B(KEYINPUT0), .ZN(n410) );
  XNOR2_X1 U438 ( .A(n410), .B(G190GAT), .ZN(n369) );
  XOR2_X1 U439 ( .A(G176GAT), .B(KEYINPUT20), .Z(n372) );
  XNOR2_X1 U440 ( .A(G43GAT), .B(KEYINPUT80), .ZN(n371) );
  XNOR2_X1 U441 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U442 ( .A(G113GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  NAND2_X1 U444 ( .A1(n475), .A2(n538), .ZN(n377) );
  XNOR2_X1 U445 ( .A(KEYINPUT26), .B(n377), .ZN(n553) );
  XOR2_X1 U446 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n378) );
  XOR2_X1 U447 ( .A(n382), .B(KEYINPUT91), .Z(n384) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U450 ( .A(n386), .B(n385), .Z(n390) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n390), .B(n389), .Z(n531) );
  XOR2_X1 U453 ( .A(n531), .B(KEYINPUT27), .Z(n417) );
  NOR2_X1 U454 ( .A1(n553), .A2(n417), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n391), .B(KEYINPUT93), .ZN(n395) );
  INV_X1 U456 ( .A(n531), .ZN(n519) );
  NOR2_X1 U457 ( .A1(n519), .A2(n538), .ZN(n392) );
  NOR2_X1 U458 ( .A1(n475), .A2(n392), .ZN(n393) );
  XNOR2_X1 U459 ( .A(KEYINPUT25), .B(n393), .ZN(n394) );
  NAND2_X1 U460 ( .A1(n395), .A2(n394), .ZN(n415) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n397) );
  XNOR2_X1 U462 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n405) );
  XOR2_X1 U464 ( .A(G141GAT), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U465 ( .A(G162GAT), .B(G85GAT), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U467 ( .A(n400), .B(G120GAT), .Z(n403) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(n401), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n414) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n407) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U474 ( .A(n408), .B(KEYINPUT1), .Z(n412) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U477 ( .A(n414), .B(n413), .Z(n516) );
  NAND2_X1 U478 ( .A1(n415), .A2(n516), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n416), .B(KEYINPUT94), .ZN(n420) );
  OR2_X1 U480 ( .A1(n516), .A2(n417), .ZN(n552) );
  XOR2_X1 U481 ( .A(n475), .B(KEYINPUT28), .Z(n522) );
  INV_X1 U482 ( .A(n522), .ZN(n512) );
  NOR2_X1 U483 ( .A1(n552), .A2(n512), .ZN(n536) );
  XNOR2_X1 U484 ( .A(n536), .B(KEYINPUT92), .ZN(n418) );
  NAND2_X1 U485 ( .A1(n418), .A2(n538), .ZN(n419) );
  NAND2_X1 U486 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U487 ( .A(KEYINPUT95), .B(n421), .ZN(n494) );
  INV_X1 U488 ( .A(n494), .ZN(n442) );
  XOR2_X1 U489 ( .A(KEYINPUT12), .B(G8GAT), .Z(n423) );
  XNOR2_X1 U490 ( .A(G1GAT), .B(G64GAT), .ZN(n422) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U492 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n425) );
  XNOR2_X1 U493 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U496 ( .A(G71GAT), .B(G183GAT), .Z(n429) );
  XNOR2_X1 U497 ( .A(G127GAT), .B(G15GAT), .ZN(n428) );
  XNOR2_X1 U498 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U499 ( .A(G22GAT), .B(G211GAT), .Z(n431) );
  XNOR2_X1 U500 ( .A(G155GAT), .B(G78GAT), .ZN(n430) );
  XNOR2_X1 U501 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U502 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U503 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n435) );
  NAND2_X1 U504 ( .A1(G231GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U506 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U507 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U508 ( .A(n441), .B(n440), .Z(n563) );
  INV_X1 U509 ( .A(n563), .ZN(n585) );
  NAND2_X1 U510 ( .A1(n442), .A2(n563), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n443), .B(KEYINPUT100), .ZN(n444) );
  NOR2_X1 U512 ( .A1(n471), .A2(n444), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n446), .B(n445), .ZN(n481) );
  NAND2_X1 U514 ( .A1(n515), .A2(n481), .ZN(n447) );
  NAND2_X1 U515 ( .A1(n534), .A2(n512), .ZN(n451) );
  XNOR2_X1 U516 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n449) );
  XOR2_X1 U517 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n448) );
  XNOR2_X1 U518 ( .A(n451), .B(n450), .ZN(G1339GAT) );
  XOR2_X1 U519 ( .A(n519), .B(KEYINPUT118), .Z(n465) );
  NOR2_X1 U520 ( .A1(n471), .A2(n563), .ZN(n453) );
  XNOR2_X1 U521 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n452) );
  XNOR2_X1 U522 ( .A(n453), .B(n452), .ZN(n456) );
  NOR2_X1 U523 ( .A1(n454), .A2(n578), .ZN(n455) );
  NAND2_X1 U524 ( .A1(n456), .A2(n455), .ZN(n463) );
  INV_X1 U525 ( .A(n578), .ZN(n556) );
  NOR2_X1 U526 ( .A1(n556), .A2(n559), .ZN(n457) );
  XNOR2_X1 U527 ( .A(n457), .B(KEYINPUT46), .ZN(n458) );
  NOR2_X1 U528 ( .A1(n585), .A2(n458), .ZN(n459) );
  NAND2_X1 U529 ( .A1(n459), .A2(n566), .ZN(n461) );
  NAND2_X1 U530 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U531 ( .A1(n465), .A2(n555), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n466), .B(KEYINPUT54), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n467), .B(KEYINPUT119), .ZN(n468) );
  NAND2_X1 U534 ( .A1(n468), .A2(n516), .ZN(n469) );
  XNOR2_X1 U535 ( .A(n469), .B(KEYINPUT64), .ZN(n476) );
  INV_X1 U536 ( .A(n586), .ZN(n470) );
  NOR2_X1 U537 ( .A1(n471), .A2(n470), .ZN(n474) );
  XNOR2_X1 U538 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n472) );
  NOR2_X1 U539 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NOR2_X2 U541 ( .A1(n538), .A2(n478), .ZN(n573) );
  NAND2_X1 U542 ( .A1(n573), .A2(n547), .ZN(n480) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n483) );
  NOR2_X1 U544 ( .A1(n556), .A2(n454), .ZN(n495) );
  NAND2_X1 U545 ( .A1(n495), .A2(n481), .ZN(n482) );
  INV_X1 U546 ( .A(n538), .ZN(n533) );
  NAND2_X1 U547 ( .A1(n511), .A2(n533), .ZN(n487) );
  XOR2_X1 U548 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n485) );
  INV_X1 U549 ( .A(G43GAT), .ZN(n484) );
  NAND2_X1 U550 ( .A1(n573), .A2(n585), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n488) );
  XNOR2_X1 U552 ( .A(n488), .B(G183GAT), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1350GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n498) );
  INV_X1 U555 ( .A(n516), .ZN(n528) );
  XOR2_X1 U556 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n492) );
  OR2_X1 U557 ( .A1(n563), .A2(n547), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(n493) );
  NOR2_X1 U559 ( .A1(n494), .A2(n493), .ZN(n514) );
  NAND2_X1 U560 ( .A1(n514), .A2(n495), .ZN(n496) );
  XOR2_X1 U561 ( .A(KEYINPUT96), .B(n496), .Z(n504) );
  NAND2_X1 U562 ( .A1(n528), .A2(n504), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n531), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(KEYINPUT98), .ZN(n501) );
  XNOR2_X1 U567 ( .A(G8GAT), .B(n501), .ZN(G1325GAT) );
  XOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U569 ( .A1(n533), .A2(n504), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  XOR2_X1 U571 ( .A(G22GAT), .B(KEYINPUT99), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n512), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(G1327GAT) );
  NAND2_X1 U574 ( .A1(n528), .A2(n511), .ZN(n508) );
  XOR2_X1 U575 ( .A(G29GAT), .B(KEYINPUT39), .Z(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  XOR2_X1 U577 ( .A(G36GAT), .B(KEYINPUT103), .Z(n510) );
  NAND2_X1 U578 ( .A1(n511), .A2(n531), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n510), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U580 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n513), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n523) );
  NOR2_X1 U583 ( .A1(n516), .A2(n523), .ZN(n517) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n517), .Z(n518) );
  XNOR2_X1 U585 ( .A(KEYINPUT42), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U586 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U587 ( .A(G64GAT), .B(n520), .Z(G1333GAT) );
  NOR2_X1 U588 ( .A1(n538), .A2(n523), .ZN(n521) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n521), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n527) );
  XOR2_X1 U591 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n525) );
  XNOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  NAND2_X1 U595 ( .A1(n534), .A2(n528), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT108), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n531), .A2(n534), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n540) );
  NAND2_X1 U603 ( .A1(n536), .A2(n555), .ZN(n537) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n548), .A2(n578), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n543) );
  NAND2_X1 U609 ( .A1(n548), .A2(n572), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n585), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n565) );
  NOR2_X1 U621 ( .A1(n556), .A2(n565), .ZN(n558) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n565), .ZN(n561) );
  XNOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U632 ( .A1(n578), .A2(n573), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n570) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT120), .B(n571), .Z(n575) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT124), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(n577), .Z(n580) );
  NAND2_X1 U643 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U646 ( .A1(n586), .A2(n454), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n584) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT125), .Z(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
endmodule

