//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT82), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G104), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n202), .A3(new_n204), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n198), .A2(G104), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(new_n205), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(KEYINPUT84), .A3(new_n202), .A4(new_n201), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n202), .B1(new_n199), .B2(new_n204), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT1), .A3(G146), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n220), .B(new_n222), .C1(G128), .C2(new_n217), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n214), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n202), .B1(new_n212), .B2(new_n201), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n221), .A2(G146), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT64), .B1(new_n217), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n233), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n235), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n204), .B1(new_n197), .B2(new_n199), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n206), .B1(new_n205), .B2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n228), .B(G101), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n230), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n220), .ZN(new_n250));
  AOI21_X1  g064(.A(G128), .B1(new_n232), .B2(new_n233), .ZN(new_n251));
  INV_X1    g065(.A(new_n222), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT67), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n254), .B(new_n222), .C1(new_n217), .C2(G128), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n225), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n215), .B1(new_n210), .B2(new_n213), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n226), .A2(new_n249), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G137), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(G137), .ZN(new_n264));
  INV_X1    g078(.A(G137), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT11), .A3(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n263), .A2(new_n266), .A3(new_n270), .A4(new_n264), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n267), .A2(KEYINPUT65), .A3(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT86), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT86), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n260), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n226), .A2(new_n249), .A3(new_n274), .A4(new_n259), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT85), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n230), .A2(new_n248), .B1(new_n257), .B2(new_n258), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n274), .A4(new_n226), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n196), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n195), .B1(new_n282), .B2(new_n285), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n214), .A2(new_n216), .A3(new_n223), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n253), .A2(new_n255), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n220), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n258), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n275), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT12), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT12), .B(new_n275), .C1(new_n289), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n190), .B(new_n191), .C1(new_n287), .C2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n190), .A2(new_n191), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n286), .A2(new_n196), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT86), .B(new_n274), .C1(new_n283), .C2(new_n226), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n278), .B1(new_n260), .B2(new_n275), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n282), .A2(new_n285), .B1(new_n295), .B2(new_n296), .ZN(new_n307));
  OAI22_X1  g121(.A1(new_n303), .A2(new_n306), .B1(new_n307), .B2(new_n196), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n286), .A2(new_n297), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n195), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n280), .A2(new_n288), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT87), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(G469), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n189), .B1(new_n302), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G237), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n193), .A3(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT27), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(KEYINPUT68), .A2(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT68), .A2(G116), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(G119), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(G119), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT2), .B(G113), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n326), .A2(G119), .ZN(new_n330));
  AND2_X1   g144(.A1(KEYINPUT68), .A2(G116), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT68), .A2(G116), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n333), .B2(G119), .ZN(new_n334));
  INV_X1    g148(.A(new_n328), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n235), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n217), .A2(new_n236), .A3(KEYINPUT64), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n241), .B1(new_n238), .B2(new_n240), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n265), .A2(G134), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n262), .A2(G137), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n271), .A2(new_n344), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n274), .A2(new_n341), .B1(new_n256), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n243), .A2(new_n273), .A3(new_n272), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(KEYINPUT70), .C1(new_n345), .C2(new_n256), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT66), .B1(new_n271), .B2(new_n344), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n256), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n243), .A2(new_n273), .A3(new_n272), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n337), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n337), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n349), .B(new_n359), .C1(new_n345), .C2(new_n256), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n352), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n322), .B1(new_n351), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT30), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n256), .A2(new_n345), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(new_n349), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n337), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(new_n360), .A3(new_n321), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n360), .ZN(new_n370));
  INV_X1    g184(.A(new_n354), .ZN(new_n371));
  INV_X1    g185(.A(new_n355), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n291), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n364), .A3(new_n349), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n346), .A2(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n370), .B(new_n322), .C1(new_n376), .C2(new_n337), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT31), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n362), .B(new_n369), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G472), .A2(G902), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(KEYINPUT32), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT32), .B1(new_n380), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n370), .B1(new_n376), .B2(new_n337), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n322), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n321), .B1(new_n351), .B2(new_n361), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n322), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n346), .A2(new_n347), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n350), .A3(new_n359), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n352), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n346), .A2(new_n337), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n360), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT28), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(KEYINPUT71), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n352), .B1(new_n395), .B2(new_n360), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n391), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G472), .B1(new_n388), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G472), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(new_n191), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n359), .B1(new_n373), .B2(new_n349), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT28), .B1(new_n409), .B2(new_n370), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n322), .B1(new_n394), .B2(new_n410), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n370), .B(new_n321), .C1(new_n376), .C2(new_n337), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n389), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n351), .A2(new_n399), .A3(new_n400), .ZN(new_n414));
  INV_X1    g228(.A(new_n401), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n390), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n408), .B(G472), .C1(new_n417), .C2(G902), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n384), .A2(new_n407), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT73), .B(G217), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(G234), .B2(new_n191), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT22), .B(G137), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(KEYINPUT23), .C1(new_n218), .C2(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT76), .ZN(new_n428));
  INV_X1    g242(.A(G119), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(G128), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT75), .B1(new_n218), .B2(G119), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n218), .A2(KEYINPUT76), .A3(G119), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT23), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n436), .A3(G110), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT77), .ZN(new_n438));
  INV_X1    g252(.A(G140), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G125), .ZN(new_n440));
  INV_X1    g254(.A(G125), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G140), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT16), .ZN(new_n443));
  OR3_X1    g257(.A1(new_n441), .A2(KEYINPUT16), .A3(G140), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(G146), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT78), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n231), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n444), .A3(new_n449), .A4(G146), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT77), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n432), .A2(new_n436), .A3(new_n452), .A4(G110), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n454), .A2(new_n218), .A3(G119), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT74), .B1(new_n429), .B2(G128), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n430), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT24), .B(G110), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n438), .A2(new_n451), .A3(new_n453), .A4(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n437), .A2(KEYINPUT77), .B1(new_n458), .B2(new_n460), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n465), .A2(KEYINPUT79), .A3(new_n451), .A4(new_n453), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G125), .B(G140), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n231), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n445), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G110), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n430), .B1(new_n427), .B2(KEYINPUT76), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT80), .B(new_n471), .C1(new_n472), .C2(new_n435), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n459), .B1(new_n457), .B2(new_n430), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n472), .B2(new_n435), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n470), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT81), .B1(new_n467), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n482), .B(new_n479), .C1(new_n464), .C2(new_n466), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n425), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n467), .A2(new_n480), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n424), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT25), .B1(new_n487), .B2(new_n191), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n489), .B(G902), .C1(new_n484), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n421), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n421), .A2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G478), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n420), .A2(new_n187), .A3(G953), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n326), .A2(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT96), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n333), .A2(G122), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n198), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(G128), .B(G143), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(G134), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(G134), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n501), .A2(KEYINPUT14), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(KEYINPUT14), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n500), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(G107), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n511), .A2(KEYINPUT13), .B1(new_n221), .B2(G128), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n511), .A2(KEYINPUT13), .ZN(new_n513));
  OAI21_X1  g327(.A(G134), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n503), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n500), .A2(new_n501), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G107), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n517), .B2(new_n502), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n498), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n500), .B1(KEYINPUT14), .B2(new_n501), .ZN(new_n520));
  INV_X1    g334(.A(new_n508), .ZN(new_n521));
  OAI21_X1  g335(.A(G107), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n522), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n502), .ZN(new_n524));
  INV_X1    g338(.A(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n526), .A3(new_n497), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT98), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n530), .B(G902), .C1(new_n519), .C2(new_n527), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n496), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n531), .A2(new_n496), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n317), .A2(new_n193), .A3(G214), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n221), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n535), .B(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n270), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n468), .B(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n231), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n445), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(KEYINPUT18), .B(G131), .C1(new_n536), .C2(KEYINPUT92), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n545));
  NAND2_X1  g359(.A1(KEYINPUT18), .A2(G131), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n538), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n468), .B(new_n231), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G113), .B(G122), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT94), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT93), .B(G104), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n536), .A2(KEYINPUT17), .A3(G131), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n540), .B2(KEYINPUT17), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n554), .B(new_n549), .C1(new_n558), .C2(new_n451), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT20), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n564), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT95), .B(G475), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n549), .B1(new_n558), .B2(new_n451), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n555), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(new_n559), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n568), .B1(new_n571), .B2(G902), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n193), .A2(G952), .ZN(new_n574));
  INV_X1    g388(.A(G234), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n317), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(G902), .B(G953), .C1(new_n575), .C2(new_n317), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n578), .B(KEYINPUT99), .Z(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n534), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G210), .B1(G237), .B2(G902), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT91), .Z(new_n585));
  AOI22_X1  g399(.A1(new_n329), .A2(new_n336), .B1(new_n227), .B2(new_n228), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n325), .B(KEYINPUT5), .C1(new_n326), .C2(G119), .ZN(new_n587));
  INV_X1    g401(.A(G113), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT5), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n330), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n587), .A2(new_n590), .B1(new_n334), .B2(new_n335), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n230), .A2(new_n586), .B1(new_n258), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G122), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n592), .A2(KEYINPUT6), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n341), .A2(G125), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n290), .A2(new_n441), .A3(new_n220), .ZN(new_n596));
  INV_X1    g410(.A(G224), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G953), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n595), .B2(new_n596), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n214), .A2(new_n216), .A3(new_n591), .ZN(new_n603));
  OAI21_X1  g417(.A(G101), .B1(new_n244), .B2(new_n246), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT4), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n210), .B2(new_n213), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n337), .A2(new_n247), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n603), .B(new_n593), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT89), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n592), .A2(new_n610), .A3(new_n593), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT6), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n614));
  INV_X1    g428(.A(new_n593), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n594), .B(new_n602), .C1(new_n612), .C2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n609), .A2(new_n611), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n600), .A2(new_n601), .B1(KEYINPUT7), .B2(new_n598), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT90), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n258), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n591), .ZN(new_n622));
  INV_X1    g436(.A(new_n336), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n587), .A2(new_n590), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n258), .B(new_n620), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n593), .B(KEYINPUT8), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n595), .A2(new_n596), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT7), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n599), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n619), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n191), .B1(new_n618), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n585), .B1(new_n617), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n612), .A2(new_n616), .ZN(new_n634));
  INV_X1    g448(.A(new_n594), .ZN(new_n635));
  INV_X1    g449(.A(new_n602), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n619), .A2(new_n627), .A3(new_n630), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n638), .B2(new_n612), .ZN(new_n639));
  INV_X1    g453(.A(new_n585), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(G214), .B1(G237), .B2(G902), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT88), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n583), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n316), .A2(new_n419), .A3(new_n494), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G101), .ZN(G3));
  NAND2_X1  g462(.A1(new_n491), .A2(new_n493), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n380), .A2(new_n191), .ZN(new_n650));
  NAND2_X1  g464(.A1(KEYINPUT100), .A2(G472), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n650), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n316), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT101), .ZN(new_n656));
  INV_X1    g470(.A(new_n643), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n640), .B1(new_n637), .B2(new_n639), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(KEYINPUT102), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n633), .A2(new_n660), .A3(new_n641), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n659), .A2(KEYINPUT103), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n662), .A2(new_n663), .A3(new_n581), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n519), .A2(new_n527), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT33), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT33), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(G478), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n495), .A2(new_n191), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n528), .B2(new_n495), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n570), .A2(new_n559), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n567), .B1(new_n672), .B2(new_n191), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n563), .B2(new_n565), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n656), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT104), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n673), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n566), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n532), .A2(new_n533), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n664), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n656), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NOR2_X1   g503(.A1(new_n481), .A2(new_n483), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n425), .A2(KEYINPUT36), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT106), .Z(new_n692));
  AND2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n492), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n653), .B1(new_n491), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n316), .A3(new_n646), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  INV_X1    g513(.A(new_n189), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n315), .A2(new_n301), .A3(new_n299), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n491), .A2(new_n695), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n579), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n576), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n566), .A2(new_n682), .A3(new_n534), .A4(new_n705), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n633), .A2(new_n660), .A3(new_n641), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n643), .B1(new_n633), .B2(new_n660), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n659), .A2(new_n661), .A3(KEYINPUT103), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(new_n419), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n707), .A2(new_n713), .A3(KEYINPUT107), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n419), .A3(new_n712), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n701), .A2(new_n702), .A3(new_n700), .A4(new_n706), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G128), .ZN(G30));
  XNOR2_X1  g534(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n642), .B(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n383), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n380), .A2(KEYINPUT32), .A3(new_n381), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n385), .A2(new_n322), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n191), .B1(new_n396), .B2(new_n321), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n491), .A3(new_n695), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n684), .A2(new_n674), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n643), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n723), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n705), .B(KEYINPUT39), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n316), .A2(KEYINPUT40), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT40), .B1(new_n316), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n737), .B(KEYINPUT109), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G143), .ZN(G45));
  AND2_X1   g553(.A1(new_n675), .A2(new_n705), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n701), .A2(new_n702), .A3(new_n700), .A4(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n716), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  NAND2_X1  g557(.A1(new_n494), .A2(new_n419), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n190), .A2(KEYINPUT110), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n286), .B1(new_n304), .B2(new_n305), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n746), .A2(new_n195), .B1(new_n297), .B2(new_n288), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n747), .B2(G902), .ZN(new_n748));
  INV_X1    g562(.A(new_n745), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n191), .B(new_n749), .C1(new_n287), .C2(new_n298), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n700), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n676), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND2_X1  g569(.A1(new_n686), .A2(new_n752), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NOR2_X1   g571(.A1(new_n662), .A2(new_n663), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n748), .A2(new_n700), .A3(new_n750), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n583), .B1(new_n491), .B2(new_n695), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(new_n419), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  NOR2_X1   g576(.A1(new_n751), .A2(new_n581), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n711), .A3(new_n712), .A4(new_n731), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n398), .A2(new_n401), .A3(new_n322), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n367), .A2(new_n360), .ZN(new_n767));
  OAI22_X1  g581(.A1(new_n767), .A2(new_n322), .B1(new_n378), .B2(KEYINPUT31), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n768), .A3(new_n369), .ZN(new_n769));
  AOI22_X1  g583(.A1(G472), .A2(new_n650), .B1(new_n769), .B2(new_n381), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n491), .A2(new_n770), .A3(new_n493), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  NAND3_X1  g588(.A1(new_n711), .A2(new_n759), .A3(new_n712), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n702), .A2(new_n740), .A3(new_n770), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  OAI211_X1 g594(.A(new_n299), .B(new_n301), .C1(new_n190), .C2(new_n308), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n642), .A2(new_n657), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n700), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n419), .A3(new_n494), .A4(new_n740), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n744), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT42), .A3(new_n740), .A4(new_n783), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  AND4_X1   g604(.A1(new_n419), .A2(new_n783), .A3(new_n494), .A4(new_n706), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n262), .ZN(G36));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n310), .B2(new_n314), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  OAI21_X1  g608(.A(G469), .B1(new_n308), .B2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT46), .B(new_n301), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT112), .A3(new_n299), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n793), .A2(new_n795), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n300), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(KEYINPUT46), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n796), .B2(new_n299), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n700), .B(new_n734), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT43), .B1(new_n671), .B2(new_n573), .ZN(new_n803));
  INV_X1    g617(.A(new_n671), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n674), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n653), .A2(new_n702), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT44), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT113), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT113), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(KEYINPUT44), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n782), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n802), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n265), .ZN(G39));
  OAI21_X1  g628(.A(new_n700), .B1(new_n800), .B2(new_n801), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT47), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(KEYINPUT47), .B(new_n700), .C1(new_n800), .C2(new_n801), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n649), .A2(new_n740), .A3(new_n782), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n419), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NAND2_X1  g637(.A1(new_n759), .A2(new_n782), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n649), .A3(new_n576), .A4(new_n729), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n675), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n574), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n771), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n806), .A2(new_n577), .A3(new_n803), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n776), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n832), .A2(new_n744), .A3(new_n824), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(KEYINPUT48), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n827), .B(new_n836), .C1(KEYINPUT48), .C2(new_n835), .ZN(new_n837));
  NOR2_X1   g651(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n722), .A2(new_n643), .A3(new_n751), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(KEYINPUT118), .A3(KEYINPUT50), .ZN(new_n841));
  NAND2_X1  g655(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n833), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n832), .A2(new_n824), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n702), .A2(new_n770), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n804), .A2(new_n573), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n844), .A2(new_n845), .B1(new_n825), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n841), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n748), .A2(new_n750), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n817), .B(new_n818), .C1(new_n700), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n782), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n829), .A2(new_n832), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n837), .B1(new_n854), .B2(KEYINPUT51), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n853), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n855), .B1(new_n861), .B2(KEYINPUT120), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(KEYINPUT120), .B2(new_n861), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n534), .A2(new_n674), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n573), .A2(new_n668), .A3(new_n670), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n645), .A3(new_n581), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n654), .A3(new_n316), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n647), .A2(new_n869), .A3(new_n697), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n760), .A2(new_n419), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n765), .A2(new_n772), .B1(new_n872), .B2(new_n776), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n684), .A2(new_n705), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n683), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n316), .A2(new_n702), .A3(new_n782), .A4(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n876), .A2(new_n419), .B1(new_n778), .B2(new_n783), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n752), .B(new_n664), .C1(new_n675), .C2(new_n685), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n871), .A2(new_n873), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n716), .A2(new_n741), .B1(new_n775), .B2(new_n777), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n711), .A2(new_n712), .A3(new_n731), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n781), .A2(new_n700), .A3(new_n705), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n730), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n719), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT107), .B1(new_n707), .B2(new_n713), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n716), .A2(new_n717), .A3(new_n715), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n882), .A2(new_n730), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n758), .A3(new_n731), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n742), .A2(new_n891), .A3(new_n779), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT52), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n791), .B1(new_n786), .B2(new_n788), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n879), .A2(new_n886), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n864), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n884), .A2(new_n885), .A3(new_n719), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n885), .B1(new_n884), .B2(new_n719), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT115), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n893), .A2(new_n901), .A3(new_n886), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n761), .B1(new_n829), .B2(new_n764), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n870), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n894), .A2(new_n904), .A3(new_n878), .A4(new_n877), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n896), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n904), .A2(new_n894), .A3(new_n878), .A4(new_n877), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n893), .A2(new_n886), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(KEYINPUT115), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n864), .A3(KEYINPUT53), .A4(new_n902), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(KEYINPUT54), .A3(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n909), .A2(new_n908), .A3(new_n896), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n896), .B2(new_n906), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n863), .A2(new_n917), .B1(G952), .B2(G953), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n850), .A2(KEYINPUT49), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT114), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n700), .A2(new_n644), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n804), .A2(new_n674), .A3(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n922), .B(new_n722), .C1(KEYINPUT49), .C2(new_n850), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n649), .A2(new_n729), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n918), .A2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n634), .A2(new_n635), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n636), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT55), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n585), .A2(G902), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n906), .A2(new_n896), .ZN(new_n931));
  INV_X1    g745(.A(new_n913), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n929), .B1(new_n933), .B2(KEYINPUT56), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  INV_X1    g749(.A(new_n929), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n935), .B(new_n936), .C1(new_n914), .C2(new_n930), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n193), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n934), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT121), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n934), .A2(new_n942), .A3(new_n937), .A4(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(G51));
  XNOR2_X1  g758(.A(new_n300), .B(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n931), .A2(new_n932), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n914), .A2(new_n915), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n747), .B(KEYINPUT122), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(G902), .A3(new_n798), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n938), .B1(new_n951), .B2(new_n952), .ZN(G54));
  NAND4_X1  g767(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n954));
  INV_X1    g768(.A(new_n560), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n938), .ZN(G60));
  NAND2_X1  g772(.A1(new_n666), .A2(new_n667), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n669), .B(KEYINPUT59), .Z(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n960), .C1(new_n947), .C2(new_n948), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n939), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n917), .B2(new_n960), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G63));
  INV_X1    g778(.A(new_n487), .ZN(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n914), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n693), .A2(new_n694), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT123), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT53), .B1(new_n910), .B2(new_n902), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n969), .B(new_n971), .C1(new_n972), .C2(new_n913), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n968), .A2(new_n973), .A3(new_n939), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT124), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n975), .A3(new_n939), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT61), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n967), .B1(new_n931), .B2(new_n932), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n938), .B1(new_n978), .B2(new_n971), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(new_n968), .C1(new_n975), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n977), .A2(new_n981), .ZN(G66));
  OAI21_X1  g796(.A(G953), .B1(new_n580), .B2(new_n597), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n904), .A2(new_n878), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n927), .B1(G898), .B2(new_n193), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(G227), .A2(G900), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n889), .A2(new_n880), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n894), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n802), .A2(new_n744), .A3(new_n881), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n703), .A2(G953), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT125), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n376), .B(new_n541), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(G953), .B(new_n989), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n995), .B2(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n989), .A2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n316), .A2(new_n734), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n852), .A2(new_n867), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(new_n787), .A3(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n990), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n738), .A2(new_n991), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(G953), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1003), .B(new_n1004), .C1(new_n1013), .C2(new_n1000), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1002), .A2(new_n1014), .ZN(G72));
  NAND4_X1  g829(.A1(new_n1012), .A2(new_n990), .A3(new_n985), .A4(new_n1008), .ZN(new_n1016));
  XNOR2_X1  g830(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(new_n405), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n726), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n386), .A2(new_n1018), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n726), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n907), .A2(new_n911), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n990), .A2(new_n985), .A3(new_n994), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n1018), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n938), .B1(new_n1025), .B2(new_n412), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(G57));
endmodule


