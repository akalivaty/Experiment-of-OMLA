//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT88), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n187), .A2(KEYINPUT3), .A3(G107), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n191), .A4(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n188), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n187), .A2(G107), .ZN(new_n195));
  OAI21_X1  g009(.A(G101), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n202), .A2(KEYINPUT1), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT89), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(new_n207), .A3(KEYINPUT1), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(G128), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n204), .B1(new_n202), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n197), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT10), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G101), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n193), .ZN(new_n216));
  INV_X1    g030(.A(new_n202), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n198), .B2(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n200), .A2(KEYINPUT64), .A3(G143), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n199), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n217), .A2(new_n218), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n214), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n204), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n205), .A2(G128), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n222), .A2(KEYINPUT69), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT69), .B1(new_n222), .B2(new_n230), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n193), .A4(new_n196), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n213), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT66), .A2(G134), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n238), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n242), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT67), .B1(new_n248), .B2(G137), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT66), .A2(G134), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT66), .A2(G134), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT67), .B(G137), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n247), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n247), .B(new_n257), .C1(new_n249), .C2(new_n253), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(KEYINPUT68), .A3(G131), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n236), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n222), .A2(new_n230), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n204), .B1(new_n266), .B2(new_n231), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n197), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n211), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT90), .A3(KEYINPUT12), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n272), .B(new_n274), .Z(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT90), .A2(KEYINPUT12), .ZN(new_n276));
  OR2_X1    g090(.A1(KEYINPUT90), .A2(KEYINPUT12), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n262), .A2(new_n269), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n263), .A2(new_n271), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n279), .A2(KEYINPUT91), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n236), .B(new_n262), .ZN(new_n281));
  INV_X1    g095(.A(new_n275), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT91), .A3(new_n279), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n280), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(G469), .A2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n275), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n263), .A2(new_n271), .A3(new_n282), .A4(new_n278), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G469), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT9), .B(G234), .Z(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(KEYINPUT87), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n303));
  INV_X1    g117(.A(G113), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(KEYINPUT71), .A2(KEYINPUT2), .A3(G113), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n305), .A2(new_n306), .B1(new_n303), .B2(new_n304), .ZN(new_n307));
  XNOR2_X1  g121(.A(G116), .B(G119), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n310), .A2(KEYINPUT5), .A3(G119), .ZN(new_n311));
  AOI211_X1 g125(.A(new_n304), .B(new_n311), .C1(KEYINPUT5), .C2(new_n308), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(new_n197), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n307), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n216), .A2(new_n318), .A3(new_n227), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(G110), .B(G122), .Z(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT92), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT92), .ZN(new_n326));
  INV_X1    g140(.A(new_n321), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n314), .A2(new_n319), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n325), .A2(new_n328), .B1(new_n321), .B2(new_n320), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n329), .B2(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n225), .A2(G125), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n267), .B2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G224), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G953), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n328), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n332), .B(KEYINPUT7), .C1(new_n333), .C2(G953), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n313), .B(new_n197), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n321), .B(KEYINPUT8), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n332), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT7), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(new_n334), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n338), .A2(new_n339), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n286), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G210), .B1(G237), .B2(G902), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT93), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n337), .A2(new_n286), .A3(new_n348), .A4(new_n346), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n301), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n273), .A3(G214), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(G143), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n257), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n356), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G131), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT17), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n356), .A2(KEYINPUT96), .A3(new_n257), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n359), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT98), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(KEYINPUT17), .A3(G131), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(KEYINPUT98), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n368), .A2(KEYINPUT16), .A3(G140), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(G146), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT97), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n365), .A2(new_n366), .A3(new_n367), .A4(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n187), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n370), .B(new_n200), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT95), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT18), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n356), .B1(new_n257), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n378), .B(new_n381), .C1(new_n361), .C2(new_n380), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n359), .A2(new_n361), .A3(new_n363), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n371), .A2(G146), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n370), .B(KEYINPUT19), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n384), .B(new_n385), .C1(G146), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n382), .ZN(new_n389));
  INV_X1    g203(.A(new_n377), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(G475), .A2(G902), .ZN(new_n393));
  XOR2_X1   g207(.A(new_n393), .B(KEYINPUT99), .Z(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(KEYINPUT20), .B2(new_n395), .ZN(new_n398));
  INV_X1    g212(.A(new_n383), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n377), .B1(new_n375), .B2(new_n382), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n286), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G475), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n310), .A2(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT100), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n310), .A2(G122), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT14), .ZN(new_n407));
  OAI21_X1  g221(.A(G107), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT102), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n406), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G107), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G128), .B(G143), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n248), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n248), .A2(new_n415), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n410), .B(new_n414), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT101), .B(KEYINPUT13), .Z(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(G128), .A3(new_n198), .ZN(new_n421));
  INV_X1    g235(.A(new_n415), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n421), .B(G134), .C1(new_n422), .C2(new_n420), .ZN(new_n423));
  INV_X1    g237(.A(new_n414), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n412), .A2(new_n413), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n416), .B(new_n423), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G217), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n296), .A2(new_n428), .A3(G953), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n419), .A2(new_n426), .A3(new_n429), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n286), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n434), .B(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n273), .A2(G952), .ZN(new_n438));
  NAND2_X1  g252(.A1(G234), .A2(G237), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(G902), .A3(G953), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n403), .A2(new_n437), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n299), .A2(new_n353), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT23), .B1(new_n203), .B2(G119), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT83), .B1(new_n203), .B2(G119), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G119), .B(G128), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT24), .B(G110), .Z(new_n453));
  OAI22_X1  g267(.A1(new_n451), .A2(G110), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n370), .A2(new_n200), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n385), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(G110), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n372), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n452), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT82), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(G137), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n461), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n286), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT25), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(G217), .B1(new_n470), .B2(G902), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT81), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT85), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n476), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n466), .A2(new_n286), .A3(new_n472), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G472), .A2(G902), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n243), .B1(G134), .B2(new_n237), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n258), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT70), .B1(new_n483), .B2(new_n267), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n234), .A2(new_n485), .A3(new_n258), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n259), .A2(new_n260), .A3(new_n225), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT73), .B1(new_n483), .B2(new_n267), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT73), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n234), .A2(new_n492), .A3(new_n258), .A4(new_n482), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n488), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n318), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(G101), .ZN(new_n499));
  INV_X1    g313(.A(G210), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n500), .A2(G237), .A3(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n499), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT76), .B(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n317), .B(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n494), .A2(new_n506), .A3(new_n489), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT74), .B(new_n318), .C1(new_n490), .C2(new_n495), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n498), .A2(new_n504), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT31), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n494), .A2(new_n506), .A3(new_n489), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n317), .B1(new_n487), .B2(new_n489), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT77), .B(KEYINPUT28), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n487), .A2(new_n489), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n318), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n516), .B2(new_n507), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n489), .B(new_n506), .C1(new_n483), .C2(new_n267), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(new_n514), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n513), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n504), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT78), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(KEYINPUT78), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n480), .B1(new_n510), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT32), .ZN(new_n529));
  INV_X1    g343(.A(new_n480), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n494), .A2(new_n489), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT30), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT74), .B1(new_n534), .B2(new_n318), .ZN(new_n535));
  INV_X1    g349(.A(new_n508), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n504), .A4(new_n507), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT31), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n509), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n521), .A2(KEYINPUT78), .A3(new_n522), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT78), .B1(new_n521), .B2(new_n522), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n530), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT32), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n529), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n506), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n531), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT79), .A3(new_n507), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT79), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n531), .A2(new_n552), .A3(new_n549), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(KEYINPUT28), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n519), .A2(new_n514), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n513), .B(new_n504), .C1(new_n517), .C2(new_n520), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n556), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n498), .A2(new_n507), .A3(new_n508), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n522), .ZN(new_n562));
  AOI211_X1 g376(.A(G902), .B(new_n558), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G472), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT80), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n558), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n561), .A2(new_n522), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n559), .A2(new_n556), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n286), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(G472), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AOI211_X1 g386(.A(KEYINPUT86), .B(new_n479), .C1(new_n548), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n545), .A2(new_n546), .ZN(new_n575));
  AOI211_X1 g389(.A(KEYINPUT32), .B(new_n530), .C1(new_n541), .C2(new_n544), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n560), .B2(new_n562), .ZN(new_n577));
  AOI211_X1 g391(.A(KEYINPUT80), .B(new_n564), .C1(new_n577), .C2(new_n566), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n570), .B1(new_n569), .B2(G472), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n575), .A2(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n479), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n448), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  AND2_X1   g398(.A1(new_n509), .A2(new_n539), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n509), .A2(new_n539), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n525), .B(new_n526), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n564), .B1(new_n587), .B2(new_n286), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n528), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n581), .A2(new_n297), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n348), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n347), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n301), .B1(new_n594), .B2(new_n352), .ZN(new_n595));
  INV_X1    g409(.A(new_n446), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n433), .A2(KEYINPUT33), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n431), .A2(new_n599), .A3(new_n432), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(G478), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n433), .A2(new_n435), .A3(new_n286), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n435), .A2(new_n286), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n403), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n592), .A2(new_n293), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  AND2_X1   g425(.A1(new_n437), .A2(new_n402), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n397), .A2(KEYINPUT103), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n395), .A2(new_n396), .ZN(new_n615));
  INV_X1    g429(.A(new_n394), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n383), .B2(new_n391), .ZN(new_n617));
  INV_X1    g431(.A(new_n396), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT103), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT104), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n614), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n615), .B1(new_n614), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n612), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n597), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n592), .A2(new_n293), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n475), .A2(new_n477), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n465), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT105), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(new_n461), .Z(new_n632));
  NOR3_X1   g446(.A1(new_n632), .A2(G902), .A3(new_n473), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n448), .A2(new_n528), .A3(new_n589), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT37), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(G110), .Z(G12));
  NAND3_X1  g452(.A1(new_n595), .A2(new_n297), .A3(new_n293), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n640));
  OR3_X1    g454(.A1(new_n444), .A2(new_n640), .A3(G900), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n640), .B1(new_n444), .B2(G900), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n440), .A3(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n612), .B(new_n643), .C1(new_n621), .C2(new_n622), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n580), .A2(new_n645), .A3(new_n635), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT107), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n634), .B1(new_n548), .B2(new_n572), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n645), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  NAND2_X1  g466(.A1(new_n351), .A2(new_n352), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT38), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n643), .B(KEYINPUT39), .Z(new_n655));
  NOR2_X1   g469(.A1(new_n298), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n301), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n575), .A2(new_n576), .ZN(new_n660));
  INV_X1    g474(.A(new_n561), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n522), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n551), .A2(new_n553), .ZN(new_n664));
  AOI21_X1  g478(.A(G902), .B1(new_n664), .B2(new_n522), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n564), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n437), .ZN(new_n669));
  INV_X1    g483(.A(new_n403), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n669), .B(new_n670), .C1(new_n656), .C2(new_n657), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n659), .A2(new_n634), .A3(new_n668), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  INV_X1    g487(.A(new_n639), .ZN(new_n674));
  INV_X1    g488(.A(new_n643), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n607), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n580), .A2(new_n635), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT108), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n648), .A2(new_n679), .A3(new_n674), .A4(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NAND3_X1  g496(.A1(new_n280), .A2(new_n284), .A3(new_n286), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(KEYINPUT109), .A3(G469), .ZN(new_n684));
  NAND2_X1  g498(.A1(KEYINPUT109), .A2(G469), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n280), .A2(new_n284), .A3(new_n286), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n297), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT110), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n684), .A2(new_n689), .A3(new_n297), .A4(new_n686), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n580), .A2(new_n691), .A3(new_n581), .A4(new_n608), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n580), .A2(new_n691), .A3(new_n581), .A4(new_n624), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT111), .B(G116), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G18));
  AND4_X1   g511(.A1(new_n447), .A2(new_n688), .A3(new_n595), .A4(new_n690), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n648), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  NOR2_X1   g514(.A1(new_n670), .A2(new_n669), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n596), .A2(new_n688), .A3(new_n595), .A4(new_n690), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n554), .A2(new_n555), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n522), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n530), .B1(new_n541), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n286), .B1(new_n510), .B2(new_n527), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n703), .B1(new_n708), .B2(new_n581), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n588), .A2(KEYINPUT112), .A3(new_n706), .A4(new_n479), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n701), .B(new_n702), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  NAND3_X1  g526(.A1(new_n691), .A2(new_n595), .A3(new_n676), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n635), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n368), .ZN(G27));
  INV_X1    g530(.A(new_n676), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n288), .B(KEYINPUT113), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n291), .A2(KEYINPUT114), .A3(G469), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT114), .B1(new_n291), .B2(G469), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n287), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n297), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n653), .A2(new_n301), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n580), .A2(new_n723), .A3(new_n581), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n479), .B1(new_n548), .B2(new_n572), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n723), .A4(new_n724), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n257), .ZN(G33));
  NOR2_X1   g545(.A1(new_n644), .A2(new_n722), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n727), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND3_X1  g548(.A1(new_n606), .A2(new_n398), .A3(new_n402), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT116), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT43), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n590), .A3(KEYINPUT44), .A4(new_n635), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n724), .B(KEYINPUT117), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT118), .ZN(new_n741));
  INV_X1    g555(.A(new_n718), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n291), .A2(KEYINPUT45), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n289), .A2(new_n290), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(G469), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n748), .A3(G469), .A4(new_n745), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n742), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n287), .B1(new_n750), .B2(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n297), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(new_n655), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n737), .A2(new_n590), .A3(new_n635), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n741), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  INV_X1    g573(.A(new_n724), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n753), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(KEYINPUT47), .B(new_n297), .C1(new_n751), .C2(new_n752), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n717), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n580), .A2(new_n581), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n768));
  INV_X1    g582(.A(new_n709), .ZN(new_n769));
  INV_X1    g583(.A(new_n710), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n737), .A2(new_n441), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n771), .A2(new_n739), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n684), .A2(new_n686), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n762), .B(new_n763), .C1(new_n297), .C2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n714), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n688), .A2(new_n690), .A3(new_n724), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT119), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT119), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n774), .A2(new_n776), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n479), .B(new_n440), .C1(new_n779), .C2(new_n780), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n667), .A3(new_n670), .A4(new_n605), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n654), .A2(new_n300), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n771), .A2(new_n691), .A3(new_n773), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT50), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n768), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n787), .B(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n782), .A3(KEYINPUT51), .A4(new_n784), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n783), .A2(new_n403), .A3(new_n606), .A4(new_n667), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(new_n792), .A3(new_n438), .A4(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n595), .A2(new_n771), .A3(new_n691), .A4(new_n773), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n781), .A2(new_n727), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT48), .ZN(new_n798));
  INV_X1    g612(.A(new_n715), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n701), .A2(new_n595), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n675), .ZN(new_n801));
  INV_X1    g615(.A(new_n722), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n668), .A2(new_n801), .A3(new_n634), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n681), .A2(new_n651), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n607), .B1(new_n669), .B2(new_n403), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n353), .A3(new_n596), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n592), .A2(new_n293), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n583), .A2(new_n636), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n711), .A2(new_n692), .A3(new_n699), .A4(new_n695), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n726), .A2(new_n729), .A3(new_n733), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n669), .B(new_n643), .C1(new_n621), .C2(new_n622), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n580), .A2(new_n299), .A3(new_n402), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n723), .A2(new_n708), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n634), .B(new_n760), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n715), .B1(new_n647), .B2(new_n650), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n681), .A4(new_n803), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n805), .A2(new_n811), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n809), .A2(new_n812), .A3(new_n817), .A4(new_n810), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n821), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n826), .A3(KEYINPUT54), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT54), .B1(new_n824), .B2(new_n826), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n796), .B(new_n798), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(G952), .A2(G953), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT120), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n775), .A2(KEYINPUT49), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n668), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n775), .A2(KEYINPUT49), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n654), .A2(new_n591), .A3(new_n735), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n300), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n833), .A2(new_n838), .ZN(G75));
  XNOR2_X1  g653(.A(new_n330), .B(new_n336), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT55), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n286), .B1(new_n824), .B2(new_n826), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(new_n350), .ZN(new_n843));
  XOR2_X1   g657(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n500), .B(new_n286), .C1(new_n824), .C2(new_n826), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n841), .B1(new_n846), .B2(KEYINPUT56), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n273), .A2(G952), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(G51));
  NAND2_X1  g664(.A1(new_n824), .A2(new_n826), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n718), .B(KEYINPUT122), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT57), .Z(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n827), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n284), .A3(new_n280), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n842), .A2(new_n749), .A3(new_n747), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n848), .B1(new_n857), .B2(new_n858), .ZN(G54));
  NAND3_X1  g673(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n391), .A3(new_n383), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .A4(new_n392), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n861), .A2(new_n849), .A3(new_n862), .ZN(G60));
  XNOR2_X1  g677(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n603), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n853), .A2(new_n827), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n598), .A2(new_n600), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n853), .A2(new_n867), .A3(new_n827), .A4(new_n865), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n869), .A2(new_n849), .A3(new_n870), .ZN(G63));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n428), .A2(new_n286), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n824), .B2(new_n826), .ZN(new_n877));
  INV_X1    g691(.A(new_n632), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n849), .B1(new_n877), .B2(new_n466), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n872), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n877), .A2(new_n466), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(KEYINPUT61), .A3(new_n849), .A4(new_n879), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(G66));
  INV_X1    g699(.A(new_n811), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n273), .B1(new_n442), .B2(G224), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n886), .A2(new_n273), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  OAI221_X1 g704(.A(new_n324), .B1(G898), .B2(new_n273), .C1(new_n329), .C2(new_n323), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(G69));
  AOI22_X1  g706(.A1(new_n741), .A2(new_n757), .B1(new_n765), .B2(new_n764), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n819), .A2(new_n894), .A3(new_n681), .A4(new_n672), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n819), .A2(new_n672), .A3(new_n681), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT62), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n573), .A2(new_n582), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n656), .A3(new_n724), .A4(new_n806), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n895), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n273), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n534), .B(new_n387), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(G900), .A2(G953), .ZN(new_n907));
  INV_X1    g721(.A(new_n727), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n754), .A2(new_n908), .A3(new_n800), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n812), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n893), .A2(new_n681), .A3(new_n819), .A4(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n906), .B(new_n907), .C1(new_n911), .C2(G953), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n901), .A2(KEYINPUT126), .A3(new_n902), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n915), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n905), .A2(new_n917), .A3(new_n912), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(G72));
  NAND2_X1  g733(.A1(G472), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT63), .Z(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n911), .B2(new_n886), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n522), .A3(new_n661), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n509), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n562), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n851), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n900), .B2(new_n886), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n662), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n849), .A2(new_n923), .A3(new_n927), .A4(new_n929), .ZN(G57));
endmodule


