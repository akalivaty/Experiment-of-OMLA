//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(KEYINPUT66), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT23), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n203), .A2(new_n204), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT24), .B1(new_n221), .B2(KEYINPUT67), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n214), .A2(new_n215), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n230), .A2(new_n231), .A3(new_n218), .A4(new_n219), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n228), .B1(new_n233), .B2(new_n214), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT27), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT68), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  AOI21_X1  g039(.A(G190gat), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT28), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n238), .A2(new_n243), .A3(G190gat), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n212), .A2(KEYINPUT26), .A3(new_n209), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n221), .B1(new_n205), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n226), .A2(new_n234), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(KEYINPUT69), .B2(KEYINPUT1), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n252), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n249), .B1(new_n242), .B2(new_n244), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n211), .A2(new_n213), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n227), .B1(new_n259), .B2(new_n232), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n260), .B2(new_n225), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n255), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT34), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT32), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n257), .A2(new_n264), .A3(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT70), .A4(new_n264), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT33), .B1(new_n271), .B2(new_n272), .ZN(new_n274));
  XOR2_X1   g073(.A(G15gat), .B(G43gat), .Z(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  AOI221_X4 g078(.A(new_n268), .B1(KEYINPUT33), .B2(new_n277), .C1(new_n271), .C2(new_n272), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n202), .B(new_n267), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n274), .A2(new_n278), .ZN(new_n282));
  INV_X1    g081(.A(new_n273), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n265), .B(KEYINPUT34), .ZN(new_n285));
  INV_X1    g084(.A(new_n280), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G1gat), .B(G29gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT0), .ZN(new_n290));
  XNOR2_X1  g089(.A(G57gat), .B(G85gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n290), .B(new_n291), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(KEYINPUT78), .Z(new_n295));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT75), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G148gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT76), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n297), .A2(new_n303), .A3(new_n307), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT77), .B(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G141gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n300), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n296), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n304), .B1(new_n314), .B2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n316), .A3(new_n255), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n306), .A2(new_n308), .B1(new_n313), .B2(new_n315), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(new_n255), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n295), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(KEYINPUT4), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n323), .A3(new_n255), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(KEYINPUT79), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n295), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n319), .A2(new_n328), .A3(new_n323), .A4(new_n255), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n256), .B1(new_n319), .B2(new_n330), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n327), .B(new_n329), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(KEYINPUT5), .B(new_n321), .C1(new_n326), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n327), .C1(new_n332), .C2(new_n333), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n340), .A3(new_n323), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n324), .A2(KEYINPUT80), .ZN(new_n342));
  AOI211_X1 g141(.A(KEYINPUT81), .B(new_n323), .C1(new_n319), .C2(new_n255), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n317), .B2(KEYINPUT4), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT6), .B(new_n293), .C1(new_n336), .C2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n293), .B1(new_n336), .B2(new_n347), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT6), .ZN(new_n350));
  INV_X1    g149(.A(new_n346), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n335), .B(new_n292), .C1(new_n351), .C2(new_n338), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G211gat), .B(G218gat), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT22), .ZN(new_n361));
  INV_X1    g160(.A(G211gat), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n364), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n358), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n261), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT74), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n261), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n369), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n370), .B1(new_n250), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n368), .B1(new_n381), .B2(new_n372), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n357), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n378), .B1(new_n375), .B2(new_n373), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n384), .B2(new_n368), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n356), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(KEYINPUT30), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n388), .A3(new_n356), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n348), .A2(new_n353), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G22gat), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT3), .B1(new_n368), .B2(new_n374), .ZN(new_n395));
  OAI211_X1 g194(.A(G228gat), .B(G233gat), .C1(new_n319), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n380), .B1(new_n319), .B2(new_n330), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n368), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n368), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT84), .B1(new_n401), .B2(new_n396), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n380), .B1(new_n365), .B2(new_n367), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n319), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n409), .A2(new_n410), .B1(new_n399), .B2(new_n368), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n408), .ZN(new_n412));
  INV_X1    g211(.A(new_n319), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n404), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n394), .B1(new_n403), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n393), .B1(new_n417), .B2(KEYINPUT85), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n402), .A3(new_n400), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n394), .A3(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n420), .A2(KEYINPUT85), .A3(new_n421), .A4(new_n393), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n267), .B1(new_n279), .B2(new_n280), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT72), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n288), .A2(new_n390), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n423), .A2(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n287), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n353), .A2(new_n348), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n387), .A2(new_n389), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n332), .A2(new_n333), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n327), .B1(new_n346), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n318), .A2(new_n320), .A3(new_n295), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT86), .B1(new_n444), .B2(new_n292), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n446), .B(new_n293), .C1(new_n440), .C2(new_n441), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT40), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI221_X1 g250(.A(new_n443), .B1(new_n449), .B2(KEYINPUT40), .C1(new_n445), .C2(new_n447), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n387), .A2(new_n349), .A3(new_n389), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n356), .B1(new_n385), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT88), .B(KEYINPUT38), .Z(new_n458));
  AOI21_X1  g257(.A(new_n368), .B1(new_n376), .B2(new_n378), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n381), .A2(new_n372), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT37), .B1(new_n460), .B2(new_n369), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n458), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n386), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n385), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n465), .B2(new_n456), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n433), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n469), .A3(new_n425), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n426), .A2(new_n287), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n427), .A2(new_n281), .A3(new_n287), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(KEYINPUT36), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n425), .A2(new_n390), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n438), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G57gat), .B(G64gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G71gat), .ZN(new_n481));
  INV_X1    g280(.A(G78gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT9), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n484), .B(new_n483), .C1(new_n479), .C2(new_n486), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT21), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G231gat), .A2(G233gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G127gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT16), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(G1gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(G1gat), .B2(new_n496), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G8gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n491), .B2(new_n490), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n495), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n504));
  INV_X1    g303(.A(G155gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G183gat), .B(G211gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n509), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT99), .ZN(new_n514));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n524));
  INV_X1    g323(.A(G85gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT97), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT97), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G85gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n524), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n531), .A2(new_n532), .B1(new_n515), .B2(KEYINPUT8), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n523), .A2(new_n530), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n530), .A2(new_n533), .A3(new_n516), .A4(new_n522), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT100), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT91), .B(G36gat), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G43gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G50gat), .ZN(new_n544));
  INV_X1    g343(.A(G50gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G43gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT15), .ZN(new_n547));
  OR3_X1    g346(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n542), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT92), .B1(new_n545), .B2(G43gat), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n543), .B2(G50gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(KEYINPUT92), .A3(G43gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT15), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n549), .A2(KEYINPUT90), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(KEYINPUT90), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n548), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n542), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n547), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n556), .B2(new_n562), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n540), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n563), .A2(new_n539), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n574));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n569), .B1(new_n567), .B2(new_n571), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n573), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n512), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n556), .A2(new_n562), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT93), .B1(new_n583), .B2(new_n501), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n563), .A2(new_n585), .A3(new_n500), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n501), .B1(new_n564), .B2(new_n566), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n587), .A2(KEYINPUT18), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n501), .ZN(new_n591));
  INV_X1    g390(.A(new_n586), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n585), .B1(new_n563), .B2(new_n500), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(new_n589), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n587), .A2(new_n589), .A3(new_n588), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(G169gat), .B(G197gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n599), .B(new_n602), .C1(new_n603), .C2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n598), .A3(new_n603), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n600), .A2(new_n601), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n590), .A2(new_n598), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n612), .B(new_n609), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n490), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n537), .A2(new_n534), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n537), .A2(new_n534), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n536), .A2(new_n490), .A3(new_n538), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT101), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n629), .A3(new_n625), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n621), .A2(new_n623), .ZN(new_n632));
  INV_X1    g431(.A(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT102), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n631), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n628), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n634), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n638), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n582), .A2(new_n617), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n478), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n468), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  INV_X1    g449(.A(new_n434), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G8gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n647), .A2(new_n434), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT42), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n655), .B1(new_n661), .B2(new_n662), .ZN(G1325gat));
  OR3_X1    g462(.A1(new_n647), .A2(G15gat), .A3(new_n431), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647), .B2(new_n474), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n647), .A2(new_n425), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  AOI21_X1  g468(.A(new_n581), .B1(new_n438), .B2(new_n477), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n617), .A2(new_n512), .A3(new_n645), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(G29gat), .A3(new_n433), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT45), .Z(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n467), .A2(new_n468), .B1(new_n424), .B2(new_n423), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n475), .B1(new_n676), .B2(new_n454), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n677), .A2(new_n474), .B1(new_n429), .B2(new_n437), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n678), .B2(new_n581), .ZN(new_n679));
  INV_X1    g478(.A(new_n581), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n478), .A2(KEYINPUT44), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n671), .B(KEYINPUT105), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n433), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n674), .A2(new_n685), .ZN(G1328gat));
  NOR3_X1   g485(.A1(new_n672), .A2(new_n434), .A3(new_n541), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT46), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n541), .B1(new_n684), .B2(new_n434), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(new_n474), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n679), .A2(new_n681), .A3(new_n691), .A4(new_n683), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G43gat), .ZN(new_n693));
  INV_X1    g492(.A(new_n672), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n431), .A2(G43gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT47), .B1(new_n697), .B2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n699), .B(new_n700), .C1(new_n693), .C2(new_n696), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n701), .ZN(G1330gat));
  OAI21_X1  g501(.A(new_n545), .B1(new_n672), .B2(new_n425), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n425), .A2(new_n545), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n684), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT48), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n708), .B(new_n703), .C1(new_n684), .C2(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1331gat));
  NAND2_X1  g509(.A1(new_n617), .A2(new_n645), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n582), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n478), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n433), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT107), .B(G57gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n434), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT108), .ZN(G1333gat));
  NOR3_X1   g521(.A1(new_n713), .A2(G71gat), .A3(new_n431), .ZN(new_n723));
  INV_X1    g522(.A(new_n713), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n691), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(G71gat), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g526(.A1(new_n713), .A2(new_n425), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n482), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n512), .A2(new_n616), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n670), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT51), .B1(new_n670), .B2(new_n730), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT109), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n526), .A2(new_n528), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n433), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n733), .A2(new_n645), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n711), .A2(new_n512), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n682), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(new_n433), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(G1336gat));
  NAND4_X1  g540(.A1(new_n679), .A2(new_n681), .A3(new_n651), .A4(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n524), .A2(new_n529), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n645), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n434), .A2(G92gat), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT110), .Z(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n731), .B2(new_n732), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g549(.A1(new_n431), .A2(G99gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n645), .A3(new_n734), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G99gat), .B1(new_n739), .B2(new_n474), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1338gat));
  NAND4_X1  g553(.A1(new_n679), .A2(new_n681), .A3(new_n430), .A4(new_n738), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G106gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n425), .A2(G106gat), .A3(new_n745), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT111), .Z(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n731), .B2(new_n732), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g560(.A(new_n512), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n624), .A2(new_n633), .A3(new_n625), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(KEYINPUT54), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n631), .A2(new_n764), .ZN(new_n765));
  AOI211_X1 g564(.A(KEYINPUT54), .B(new_n633), .C1(new_n624), .C2(new_n625), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(new_n767), .A3(new_n639), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n626), .A2(new_n769), .A3(new_n628), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT112), .B1(new_n770), .B2(new_n638), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n641), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n767), .B1(new_n766), .B2(new_n639), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n770), .A2(KEYINPUT112), .A3(new_n638), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n776), .A2(new_n777), .B1(new_n631), .B2(new_n764), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n640), .B1(new_n778), .B2(KEYINPUT55), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n772), .A2(new_n773), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n775), .A2(new_n781), .A3(new_n616), .A4(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n594), .B2(new_n597), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n587), .A2(KEYINPUT114), .A3(new_n591), .A4(new_n596), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n587), .A2(new_n588), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n589), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n608), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n599), .A2(new_n610), .A3(new_n602), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n645), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n680), .B1(new_n783), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n781), .A3(new_n782), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n680), .A2(new_n789), .A3(new_n790), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n762), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n617), .A2(new_n512), .A3(new_n581), .A4(new_n745), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n651), .A2(new_n433), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n432), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(G113gat), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n800), .A2(new_n801), .A3(new_n617), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n433), .B1(new_n796), .B2(new_n797), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n288), .A2(new_n425), .A3(new_n427), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT115), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n434), .A3(new_n616), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n802), .B1(new_n808), .B2(new_n801), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n800), .A2(new_n810), .A3(new_n745), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n434), .A3(new_n645), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n810), .ZN(G1341gat));
  OAI21_X1  g612(.A(G127gat), .B1(new_n800), .B2(new_n762), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n807), .A2(new_n434), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n762), .A2(G127gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(G1342gat));
  OAI21_X1  g616(.A(G134gat), .B1(new_n800), .B2(new_n581), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT116), .Z(new_n819));
  NOR2_X1   g618(.A1(new_n651), .A2(new_n581), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(G134gat), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n807), .A2(KEYINPUT56), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n807), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(G1343gat));
  OAI21_X1  g624(.A(KEYINPUT117), .B1(new_n778), .B2(KEYINPUT55), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n772), .A2(new_n827), .A3(new_n773), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n779), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n826), .A2(new_n779), .A3(new_n828), .A4(KEYINPUT118), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n616), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n680), .B1(new_n833), .B2(new_n791), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n762), .B1(new_n834), .B2(new_n795), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n797), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT57), .A4(new_n430), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n474), .A2(new_n799), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n840), .B(new_n425), .C1(new_n835), .C2(new_n797), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n425), .B1(new_n796), .B2(new_n797), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT119), .B1(new_n842), .B2(KEYINPUT57), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n838), .B(new_n839), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G141gat), .B1(new_n844), .B2(new_n617), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n691), .A2(new_n425), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n803), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n651), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n617), .A2(G141gat), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT58), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n845), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n310), .A2(KEYINPUT59), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n844), .B2(new_n745), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n839), .A2(KEYINPUT122), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n839), .A2(KEYINPUT122), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n745), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n842), .A2(KEYINPUT57), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n425), .B1(new_n835), .B2(new_n797), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n299), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n857), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n310), .A3(new_n645), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT121), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1345gat));
  OAI21_X1  g668(.A(G155gat), .B1(new_n844), .B2(new_n762), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n848), .A2(new_n505), .A3(new_n512), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1346gat));
  OAI21_X1  g671(.A(G162gat), .B1(new_n844), .B2(new_n581), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n821), .A2(G162gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n847), .B2(new_n874), .ZN(G1347gat));
  NAND2_X1  g674(.A1(new_n798), .A2(new_n432), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n468), .A2(new_n434), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT123), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n203), .B1(new_n879), .B2(new_n616), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT124), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n798), .A2(new_n877), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(new_n805), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n203), .A3(new_n616), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1348gat));
  INV_X1    g684(.A(new_n879), .ZN(new_n886));
  OAI21_X1  g685(.A(G176gat), .B1(new_n886), .B2(new_n745), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n204), .A3(new_n645), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1349gat));
  NOR2_X1   g688(.A1(new_n762), .A2(new_n238), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n883), .A2(new_n890), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n891));
  OAI21_X1  g690(.A(G183gat), .B1(new_n886), .B2(new_n762), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT126), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n893), .B(new_n895), .ZN(G1350gat));
  AOI21_X1  g695(.A(new_n217), .B1(new_n879), .B2(new_n680), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT61), .Z(new_n898));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n217), .A3(new_n680), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1351gat));
  INV_X1    g699(.A(G197gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n878), .A2(new_n691), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n864), .A2(new_n616), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n903), .B2(KEYINPUT127), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(KEYINPUT127), .B2(new_n903), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n882), .A2(new_n846), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n901), .A3(new_n616), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1352gat));
  INV_X1    g707(.A(G204gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n906), .A2(new_n909), .A3(new_n645), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT62), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n864), .A2(new_n902), .ZN(new_n912));
  OAI21_X1  g711(.A(G204gat), .B1(new_n912), .B2(new_n745), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(KEYINPUT62), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n906), .A2(new_n362), .A3(new_n512), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n864), .A2(new_n512), .A3(new_n902), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT63), .B1(new_n917), .B2(G211gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1354gat));
  OAI21_X1  g719(.A(G218gat), .B1(new_n912), .B2(new_n581), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n363), .A3(new_n680), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1355gat));
endmodule


