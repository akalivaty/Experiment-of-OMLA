//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT65), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n204), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NOR3_X1   g0019(.A1(new_n207), .A2(new_n211), .A3(new_n219), .ZN(G361));
  XNOR2_X1  g0020(.A(G238), .B(G244), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT2), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n225), .B(new_n228), .Z(G358));
  XOR2_X1   g0029(.A(G68), .B(G77), .Z(new_n230));
  XNOR2_X1  g0030(.A(G50), .B(G58), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XNOR2_X1  g0033(.A(G107), .B(G116), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G351));
  XNOR2_X1  g0036(.A(KEYINPUT3), .B(G33), .ZN(new_n237));
  NAND2_X1  g0037(.A1(G238), .A2(G1698), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n237), .B(new_n238), .C1(new_n224), .C2(G1698), .ZN(new_n239));
  NAND2_X1  g0039(.A1(G33), .A2(G41), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n240), .A2(G1), .A3(G13), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  OAI211_X1 g0042(.A(new_n239), .B(new_n242), .C1(G107), .C2(new_n237), .ZN(new_n243));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(new_n241), .A3(G274), .ZN(new_n247));
  INV_X1    g0047(.A(G244), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n243), .B(new_n247), .C1(new_n248), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G169), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G179), .B2(new_n252), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n210), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n249), .B2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G77), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(new_n209), .A3(G1), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(G77), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT15), .B(G87), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(new_n209), .A3(G33), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n269), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n263), .B1(new_n272), .B2(new_n257), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n255), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n252), .A2(G200), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(new_n275), .C1(new_n276), .C2(new_n252), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT69), .Z(new_n279));
  INV_X1    g0079(.A(KEYINPUT12), .ZN(new_n280));
  OAI21_X1  g0080(.A(G68), .B1(new_n258), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n280), .A2(new_n260), .A3(G1), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n262), .A2(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n257), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n209), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  INV_X1    g0091(.A(new_n270), .ZN(new_n292));
  INV_X1    g0092(.A(G50), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n283), .B1(new_n290), .B2(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n287), .B1(KEYINPUT11), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(KEYINPUT11), .B2(new_n295), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G226), .A2(G1698), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n224), .B2(G1698), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n237), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n242), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n299), .A2(new_n237), .B1(G33), .B2(G97), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT70), .B1(new_n305), .B2(new_n241), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G238), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n247), .B1(new_n308), .B2(new_n251), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT71), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n247), .B(new_n311), .C1(new_n308), .C2(new_n251), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n304), .A2(new_n306), .B1(new_n310), .B2(new_n312), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n297), .B1(new_n319), .B2(G200), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n321), .A3(KEYINPUT13), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT72), .B1(new_n316), .B2(new_n317), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(G190), .A4(new_n318), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n316), .A2(new_n317), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT14), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n253), .B1(new_n315), .B2(new_n318), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n322), .A2(new_n323), .A3(G179), .A4(new_n318), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n297), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G50), .A2(G58), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n209), .B1(new_n337), .B2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n268), .A2(new_n290), .B1(new_n339), .B2(new_n292), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n289), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n257), .B(KEYINPUT67), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n262), .ZN(new_n343));
  OAI21_X1  g0143(.A(G50), .B1(new_n209), .B2(G1), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n341), .B1(G50), .B2(new_n262), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT9), .ZN(new_n346));
  INV_X1    g0146(.A(G222), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n237), .B1(new_n347), .B2(G1698), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  OR2_X1    g0149(.A1(KEYINPUT66), .A2(G223), .ZN(new_n350));
  NAND2_X1  g0150(.A1(KEYINPUT66), .A2(G223), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n242), .B1(G77), .B2(new_n237), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n251), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G226), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n353), .A2(new_n247), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G190), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n346), .B(new_n357), .C1(new_n358), .C2(new_n356), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT10), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n345), .C1(G169), .C2(new_n356), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n279), .A2(new_n336), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n343), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n268), .B1(new_n249), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n366), .B1(new_n261), .B2(new_n268), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n257), .ZN(new_n369));
  XNOR2_X1  g0169(.A(G58), .B(G68), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(G20), .B1(G159), .B2(new_n270), .ZN(new_n371));
  INV_X1    g0171(.A(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G33), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT7), .B1(new_n376), .B2(new_n209), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(G20), .ZN(new_n379));
  OR2_X1    g0179(.A1(KEYINPUT73), .A2(G33), .ZN(new_n380));
  NAND2_X1  g0180(.A1(KEYINPUT73), .A2(G33), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT3), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n374), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n385));
  AOI21_X1  g0185(.A(G33), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n379), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT76), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n385), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n372), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(KEYINPUT73), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT73), .A2(G33), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n374), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT76), .A3(new_n379), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n377), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n371), .B1(new_n398), .B2(new_n282), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n369), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n371), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n380), .A2(KEYINPUT3), .A3(new_n381), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n384), .A2(G33), .A3(new_n385), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n209), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n282), .B1(new_n406), .B2(KEYINPUT7), .ZN(new_n407));
  AOI211_X1 g0207(.A(KEYINPUT7), .B(G20), .C1(new_n403), .C2(new_n404), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n402), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(G20), .B1(new_n403), .B2(new_n404), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n413), .B2(new_n378), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT16), .B(new_n371), .C1(new_n414), .C2(new_n408), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n368), .B1(new_n401), .B2(new_n417), .ZN(new_n418));
  MUX2_X1   g0218(.A(G223), .B(G226), .S(G1698), .Z(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n403), .A3(new_n404), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n241), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n247), .B1(new_n224), .B2(new_n251), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n361), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n253), .B1(new_n422), .B2(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n427), .B(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT18), .B1(new_n418), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n415), .B(new_n411), .ZN(new_n431));
  INV_X1    g0231(.A(new_n377), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT76), .B1(new_n396), .B2(new_n379), .ZN(new_n433));
  INV_X1    g0233(.A(new_n379), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n388), .B(new_n434), .C1(new_n392), .C2(new_n395), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n402), .B1(new_n436), .B2(G68), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n257), .B1(new_n437), .B2(KEYINPUT16), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n367), .B1(new_n431), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n427), .B(KEYINPUT77), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n430), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n424), .A2(G190), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n358), .B2(new_n424), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n367), .B(new_n447), .C1(new_n431), .C2(new_n438), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n364), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT19), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n209), .B1(new_n301), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT84), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n209), .C1(new_n301), .C2(new_n452), .ZN(new_n456));
  INV_X1    g0256(.A(G87), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n452), .B1(new_n290), .B2(new_n458), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n282), .A2(G20), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n403), .A2(new_n404), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n257), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n264), .B(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n261), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n372), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n266), .A2(new_n262), .A3(new_n342), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n249), .A2(G45), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G250), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n242), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n245), .A2(G1), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n241), .A2(G274), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  AND2_X1   g0281(.A1(G1), .A2(G13), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n240), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n478), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n477), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G238), .A2(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n248), .B2(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n403), .A2(new_n488), .A3(new_n404), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n380), .A2(new_n381), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G116), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(G179), .B(new_n486), .C1(new_n492), .C2(new_n241), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n484), .B1(new_n483), .B2(new_n478), .ZN(new_n494));
  AND4_X1   g0294(.A1(new_n484), .A2(new_n241), .A3(G274), .A4(new_n478), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n494), .A2(new_n495), .B1(new_n242), .B2(new_n476), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n241), .B1(new_n489), .B2(new_n491), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n493), .B1(new_n498), .B2(new_n253), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT85), .A4(new_n468), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n474), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n466), .A2(new_n468), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n498), .A2(G190), .ZN(new_n503));
  OAI21_X1  g0303(.A(G200), .B1(new_n496), .B2(new_n497), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n342), .A2(new_n262), .A3(new_n470), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n505), .A2(new_n457), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT86), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n501), .A2(new_n507), .A3(KEYINPUT86), .ZN(new_n511));
  INV_X1    g0311(.A(G257), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G1698), .ZN(new_n513));
  INV_X1    g0313(.A(G250), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n349), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n403), .A2(new_n404), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n490), .A2(G294), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n241), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT88), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT79), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n244), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n478), .B(new_n527), .C1(KEYINPUT5), .C2(new_n244), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT78), .B1(new_n529), .B2(new_n475), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n526), .A2(new_n528), .A3(new_n530), .A4(new_n483), .ZN(new_n531));
  AOI21_X1  g0331(.A(G41), .B1(new_n522), .B2(new_n524), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n478), .B1(KEYINPUT5), .B2(new_n244), .ZN(new_n533));
  OAI211_X1 g0333(.A(G264), .B(new_n241), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n520), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n518), .A2(new_n519), .ZN(new_n538));
  OAI21_X1  g0338(.A(G169), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n516), .A2(new_n517), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n242), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT89), .B1(new_n542), .B2(new_n361), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n535), .A2(new_n518), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT89), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(G179), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n539), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n505), .A2(new_n459), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n261), .A2(new_n459), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n549), .B(KEYINPUT25), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n457), .A2(G20), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n376), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n490), .A2(new_n209), .A3(G116), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n557));
  OR3_X1    g0357(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT22), .A4(new_n553), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT87), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT22), .B1(new_n237), .B2(new_n553), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n557), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT87), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n565), .A2(new_n560), .A3(new_n566), .A4(new_n556), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n562), .A2(KEYINPUT24), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n257), .B1(new_n562), .B2(KEYINPUT24), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n551), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n547), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G270), .B(new_n241), .C1(new_n532), .C2(new_n533), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n531), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n349), .A2(G264), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n512), .A2(new_n349), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n403), .A2(new_n404), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n376), .A2(G303), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n242), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n369), .A2(new_n262), .A3(G116), .A4(new_n470), .ZN(new_n581));
  INV_X1    g0381(.A(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n261), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n256), .A2(new_n210), .B1(G20), .B2(new_n582), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n209), .C1(G33), .C2(new_n458), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT20), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n581), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n580), .A2(G169), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n573), .A2(new_n579), .A3(G179), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n589), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n580), .A2(KEYINPUT21), .A3(G169), .A4(new_n589), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n531), .A2(new_n572), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n241), .B1(new_n576), .B2(new_n577), .ZN(new_n598));
  OAI21_X1  g0398(.A(G200), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n589), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n599), .B(new_n600), .C1(new_n580), .C2(new_n276), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n592), .A2(new_n595), .A3(new_n596), .A4(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n510), .A2(new_n511), .A3(new_n571), .A4(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n403), .A2(new_n404), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT4), .B1(new_n604), .B2(G244), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n349), .A2(KEYINPUT4), .A3(G244), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n237), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT4), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n237), .B2(G250), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n585), .C1(new_n610), .C2(new_n349), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n242), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n241), .C1(new_n532), .C2(new_n533), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n531), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(G190), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n612), .A2(KEYINPUT82), .A3(G190), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n262), .A2(G97), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n505), .B2(new_n458), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT6), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n624), .A2(new_n458), .A3(G107), .ZN(new_n625));
  XNOR2_X1  g0425(.A(G97), .B(G107), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n624), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n627), .A2(new_n209), .B1(new_n291), .B2(new_n292), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n398), .B2(new_n459), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n623), .B1(new_n630), .B2(new_n257), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n531), .A2(new_n613), .A3(KEYINPUT80), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT80), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n614), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n612), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT81), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(G200), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n635), .B2(G200), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n620), .B(new_n631), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n541), .A2(KEYINPUT88), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n536), .A3(new_n520), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n641), .A2(G190), .B1(G200), .B2(new_n544), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n642), .B(new_n551), .C1(new_n568), .C2(new_n569), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n612), .A2(new_n361), .A3(new_n634), .A4(new_n632), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n585), .B1(new_n376), .B2(new_n606), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT4), .B1(new_n376), .B2(new_n514), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(G1698), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n609), .B1(new_n405), .B2(new_n248), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n241), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n253), .B1(new_n649), .B2(new_n614), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n623), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n628), .B1(new_n436), .B2(G107), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n369), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n639), .A2(new_n643), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n603), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n451), .A2(new_n657), .ZN(G372));
  INV_X1    g0458(.A(KEYINPUT92), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n418), .A2(new_n429), .A3(KEYINPUT18), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n430), .A2(new_n442), .A3(KEYINPUT92), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n448), .B(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n326), .A2(new_n274), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n335), .A2(new_n297), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n360), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n363), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n651), .A2(new_n673), .A3(new_n654), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n644), .A2(new_n650), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT91), .B1(new_n631), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n571), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n570), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n679), .B1(new_n684), .B2(new_n656), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n507), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n499), .A2(new_n472), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n501), .A2(new_n507), .A3(KEYINPUT86), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT86), .B1(new_n501), .B2(new_n507), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n631), .A2(new_n675), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n688), .B1(new_n693), .B2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n451), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n672), .A2(new_n696), .ZN(G369));
  NAND3_X1  g0497(.A1(new_n249), .A2(new_n209), .A3(G13), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(G213), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n570), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n643), .A2(new_n571), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n703), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n680), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n682), .A2(new_n683), .A3(new_n706), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n589), .A2(new_n703), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT93), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n680), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n592), .A2(new_n595), .A3(new_n596), .A4(new_n601), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n705), .B1(new_n571), .B2(new_n706), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n205), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n460), .A2(G116), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n722), .A2(new_n249), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n208), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n722), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n639), .A2(new_n643), .A3(new_n655), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n547), .A2(new_n570), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n714), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n730), .A2(new_n691), .A3(new_n732), .A4(new_n706), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  INV_X1    g0534(.A(new_n534), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n518), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n612), .A2(new_n498), .A3(new_n736), .A4(new_n615), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n737), .B2(new_n593), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n498), .A2(new_n736), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n649), .A2(new_n614), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n594), .A3(KEYINPUT30), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n498), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n635), .A2(new_n742), .A3(new_n542), .A4(new_n580), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n738), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n703), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(KEYINPUT94), .B(new_n729), .C1(new_n733), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n733), .A2(new_n749), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(G330), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n703), .B1(new_n686), .B2(new_n694), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n507), .A2(new_n687), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n731), .B2(new_n680), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n656), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n510), .A2(new_n678), .A3(new_n692), .A4(new_n511), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n674), .B2(new_n676), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n761), .B(new_n687), .C1(new_n762), .C2(new_n678), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT96), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n762), .A2(new_n678), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(KEYINPUT96), .A3(new_n687), .A4(new_n761), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n703), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT29), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n750), .B(new_n753), .C1(new_n756), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n728), .B1(new_n770), .B2(G1), .ZN(G364));
  NOR2_X1   g0571(.A1(new_n260), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n249), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n722), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n717), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n715), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT98), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n210), .B1(G20), .B2(new_n253), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n232), .A2(new_n245), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n721), .A2(new_n604), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n784), .B(new_n786), .C1(new_n245), .C2(new_n726), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n205), .A2(new_n237), .ZN(new_n788));
  INV_X1    g0588(.A(G355), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n788), .A2(new_n789), .B1(G116), .B2(new_n205), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n783), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n209), .B1(new_n792), .B2(G190), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n458), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n209), .A2(G190), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n792), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n799));
  XNOR2_X1  g0599(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n276), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n794), .B(new_n800), .C1(G50), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n361), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n795), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n801), .A2(G190), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n237), .B1(new_n805), .B2(new_n291), .C1(new_n807), .C2(new_n282), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n209), .A2(new_n276), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n358), .A2(G179), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G87), .ZN(new_n813));
  INV_X1    g0613(.A(G58), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n809), .A2(new_n804), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n795), .A2(new_n810), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n808), .B(new_n816), .C1(G107), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G303), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n811), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n822), .A2(new_n817), .B1(new_n805), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n796), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n821), .B(new_n824), .C1(G329), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G322), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n376), .B1(new_n815), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT33), .B(G317), .Z(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n807), .A2(new_n829), .B1(new_n830), .B2(new_n793), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n828), .B(new_n831), .C1(G326), .C2(new_n802), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n803), .A2(new_n819), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n782), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n791), .B(new_n776), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT100), .ZN(new_n836));
  INV_X1    g0636(.A(new_n781), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n715), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n778), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  OR2_X1    g0640(.A1(new_n782), .A2(new_n779), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n776), .B1(G77), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT101), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n237), .B(new_n794), .C1(G107), .C2(new_n812), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G87), .A2(new_n818), .B1(new_n825), .B2(G311), .ZN(new_n845));
  INV_X1    g0645(.A(new_n815), .ZN(new_n846));
  INV_X1    g0646(.A(new_n805), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G294), .A2(new_n846), .B1(new_n847), .B2(G116), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G283), .A2(new_n806), .B1(new_n802), .B2(G303), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n844), .A2(new_n845), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G68), .A2(new_n818), .B1(new_n825), .B2(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n293), .B2(new_n811), .ZN(new_n852));
  INV_X1    g0652(.A(new_n793), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n405), .B(new_n852), .C1(G58), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT102), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G143), .A2(new_n846), .B1(new_n847), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(new_n802), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n857), .B2(new_n858), .C1(new_n339), .C2(new_n807), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT34), .Z(new_n860));
  OAI21_X1  g0660(.A(new_n850), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n782), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n274), .A2(new_n703), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n277), .B1(new_n273), .B2(new_n706), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n274), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n843), .B(new_n862), .C1(new_n867), .C2(new_n780), .ZN(new_n868));
  INV_X1    g0668(.A(new_n507), .ZN(new_n869));
  INV_X1    g0669(.A(new_n680), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n570), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT90), .B1(new_n547), .B2(new_n570), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n730), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n869), .B1(new_n874), .B2(new_n679), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n693), .A2(KEYINPUT26), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n687), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n706), .B(new_n867), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n866), .B(KEYINPUT103), .Z(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n754), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n753), .A2(new_n750), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT105), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n776), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n881), .A2(new_n886), .A3(new_n882), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(KEYINPUT105), .A3(new_n882), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n881), .B2(new_n882), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n868), .B1(new_n885), .B2(new_n890), .ZN(G384));
  INV_X1    g0691(.A(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n627), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(G20), .A3(G116), .A4(new_n482), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT106), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n894), .A2(new_n895), .B1(new_n892), .B2(new_n627), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  XOR2_X1   g0697(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n726), .B(G77), .C1(new_n814), .C2(new_n282), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n293), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n249), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  INV_X1    g0704(.A(new_n701), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n289), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n431), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n368), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n667), .B2(new_n443), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n439), .A2(new_n441), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n701), .B(KEYINPUT108), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n439), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n914), .A3(new_n448), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n368), .B(new_n446), .C1(new_n401), .C2(new_n417), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n916), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n441), .A2(new_n905), .B1(new_n907), .B2(new_n368), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n915), .A2(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n910), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n448), .B(KEYINPUT92), .C1(new_n418), .C2(new_n912), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n915), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n401), .A2(new_n417), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n912), .B1(new_n925), .B2(new_n367), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n917), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(new_n659), .A3(KEYINPUT37), .A4(new_n911), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n662), .A2(new_n449), .A3(new_n663), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n904), .B(new_n921), .C1(new_n931), .C2(KEYINPUT38), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT38), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n908), .B1(new_n444), .B2(new_n449), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n915), .A2(new_n916), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n918), .A2(new_n919), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n933), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n921), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n335), .A2(new_n297), .A3(new_n706), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n297), .A2(new_n703), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n669), .A2(new_n325), .A3(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n297), .B(new_n703), .C1(new_n326), .C2(new_n335), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n878), .B2(new_n863), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n950), .A2(new_n939), .B1(new_n665), .B2(new_n912), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n756), .A2(new_n451), .A3(new_n769), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n672), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n921), .B1(new_n931), .B2(KEYINPUT38), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n866), .B1(new_n946), .B2(new_n947), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(new_n752), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n958), .A2(KEYINPUT40), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n920), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n910), .B2(new_n920), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n963));
  AOI22_X1  g0763(.A1(new_n956), .A2(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n451), .A3(new_n752), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(G330), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n451), .B2(new_n752), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n955), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n249), .B2(new_n772), .C1(new_n955), .C2(new_n968), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n903), .B1(new_n971), .B2(new_n972), .ZN(G367));
  OAI211_X1 g0773(.A(new_n639), .B(new_n655), .C1(new_n631), .C2(new_n706), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n692), .A2(new_n703), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(new_n708), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n974), .A2(new_n571), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n703), .B1(new_n980), .B2(new_n655), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n978), .B2(KEYINPUT42), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n502), .A2(new_n506), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n703), .ZN(new_n984));
  MUX2_X1   g0784(.A(new_n688), .B(new_n758), .S(new_n984), .Z(new_n985));
  AOI22_X1  g0785(.A1(new_n979), .A2(new_n982), .B1(KEYINPUT43), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n719), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n976), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n988), .B(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n722), .B(KEYINPUT41), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n710), .A2(new_n976), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT45), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n976), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT44), .B1(new_n710), .B2(new_n976), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n994), .A2(new_n997), .A3(KEYINPUT111), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT111), .B1(new_n994), .B2(new_n997), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n989), .A3(new_n999), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n994), .A2(new_n997), .A3(new_n989), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(KEYINPUT112), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n717), .A2(KEYINPUT113), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n716), .B(KEYINPUT113), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n707), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n708), .B1(new_n718), .B2(new_n1005), .ZN(new_n1006));
  MUX2_X1   g0806(.A(new_n1003), .B(new_n1004), .S(new_n1006), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n770), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1002), .B(new_n1009), .C1(KEYINPUT112), .C2(new_n1000), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n992), .B1(new_n1010), .B2(new_n770), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n991), .B1(new_n1011), .B2(new_n774), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n783), .B1(new_n205), .B2(new_n467), .C1(new_n786), .C2(new_n228), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n776), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n812), .A2(G116), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT46), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(new_n1016), .B1(new_n802), .B2(G311), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n1016), .B2(new_n1015), .C1(new_n459), .C2(new_n793), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n458), .A2(new_n817), .B1(new_n805), .B2(new_n822), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n815), .A2(new_n820), .B1(new_n796), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n405), .B1(new_n807), .B2(new_n830), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n853), .A2(G68), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n237), .C1(new_n293), .C2(new_n805), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n811), .A2(new_n814), .B1(new_n796), .B2(new_n858), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n815), .A2(new_n339), .B1(new_n817), .B2(new_n291), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n802), .A2(G143), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n807), .B2(new_n797), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1023), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1014), .B1(new_n985), .B2(new_n837), .C1(new_n1032), .C2(new_n834), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1012), .A2(new_n1033), .ZN(G387));
  NOR2_X1   g0834(.A1(new_n770), .A2(new_n1007), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1008), .A2(new_n722), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(KEYINPUT115), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT115), .B2(new_n1036), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n718), .A2(new_n837), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n788), .A2(new_n723), .B1(G107), .B2(new_n205), .ZN(new_n1040));
  AOI211_X1 g0840(.A(G45), .B(new_n724), .C1(G68), .C2(G77), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1046), .A2(new_n785), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n225), .A2(G45), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n783), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n776), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n811), .A2(new_n830), .B1(new_n793), .B2(new_n822), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G317), .A2(new_n846), .B1(new_n847), .B2(G303), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n857), .B2(new_n827), .C1(new_n823), .C2(new_n807), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G116), .A2(new_n818), .B1(new_n825), .B2(G326), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1059), .A2(new_n405), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n805), .A2(new_n282), .B1(new_n796), .B2(new_n339), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G50), .B2(new_n846), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n266), .A2(new_n853), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n811), .A2(new_n291), .B1(new_n817), .B2(new_n458), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n405), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n269), .A2(new_n806), .B1(G159), .B2(new_n802), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1051), .B1(new_n1070), .B2(new_n782), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1007), .A2(new_n774), .B1(new_n1039), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1038), .A2(new_n1072), .ZN(G393));
  NOR2_X1   g0873(.A1(new_n994), .A2(new_n997), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n719), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1008), .B1(new_n1075), .B2(new_n1001), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1010), .A2(new_n722), .A3(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1075), .A2(new_n773), .A3(new_n1001), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n977), .A2(new_n781), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n783), .B1(new_n458), .B2(new_n205), .C1(new_n786), .C2(new_n235), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n776), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT116), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n853), .A2(G77), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n604), .A2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G87), .A2(new_n818), .B1(new_n825), .B2(G143), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n282), .B2(new_n811), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n807), .A2(new_n293), .B1(new_n805), .B2(new_n268), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1084), .B(new_n1086), .C1(KEYINPUT117), .C2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n857), .A2(new_n339), .B1(new_n815), .B2(new_n797), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(KEYINPUT117), .C2(new_n1087), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n376), .B1(new_n817), .B2(new_n459), .C1(new_n807), .C2(new_n820), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G116), .B2(new_n853), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n857), .A2(new_n1020), .B1(new_n815), .B2(new_n823), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n805), .A2(new_n830), .B1(new_n796), .B2(new_n827), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G283), .B2(new_n812), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1082), .B1(new_n1102), .B2(new_n782), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1078), .B1(new_n1079), .B2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1077), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n747), .A2(new_n748), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n657), .B2(new_n706), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT94), .B1(new_n1108), .B2(new_n729), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n752), .A2(new_n751), .A3(G330), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n866), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n948), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n863), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n768), .B2(new_n865), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n752), .A2(G330), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n949), .B1(new_n1115), .B2(new_n879), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1115), .A2(new_n866), .A3(new_n949), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n867), .B1(new_n753), .B2(new_n750), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n949), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1113), .B1(new_n754), .B2(new_n867), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT120), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1115), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n957), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1111), .B2(new_n948), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT120), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1121), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1117), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n451), .A2(new_n1123), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n953), .A2(new_n672), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n932), .B(new_n940), .C1(new_n943), .C2(new_n950), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n942), .B(KEYINPUT119), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n956), .B(new_n1135), .C1(new_n1114), .C2(new_n949), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n1112), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n904), .B1(new_n938), .B2(new_n921), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n930), .A2(new_n926), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n927), .A2(new_n911), .B1(new_n922), .B2(KEYINPUT37), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n448), .B1(new_n418), .B2(new_n912), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n418), .A2(new_n429), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT92), .A4(new_n916), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n960), .B1(new_n1145), .B2(new_n933), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1138), .B1(new_n1146), .B2(new_n904), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n942), .B1(new_n1121), .B2(new_n949), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n933), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1134), .B1(new_n1149), .B2(new_n921), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n865), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n703), .B(new_n1151), .C1(new_n765), .C2(new_n767), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n948), .B1(new_n1152), .B2(new_n1113), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1147), .A2(new_n1148), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1137), .B1(new_n1154), .B2(new_n1124), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n722), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n776), .B1(new_n269), .B2(new_n841), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n811), .A2(new_n339), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n825), .A2(G125), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n847), .A2(new_n1165), .B1(new_n818), .B2(G50), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n376), .B1(new_n846), .B2(G132), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n802), .B1(new_n806), .B2(G137), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n797), .C2(new_n793), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G116), .A2(new_n846), .B1(new_n825), .B2(G294), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n282), .B2(new_n817), .C1(new_n458), .C2(new_n805), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G107), .A2(new_n806), .B1(new_n802), .B2(G283), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n813), .A2(new_n1173), .A3(new_n1083), .A4(new_n376), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1167), .A2(new_n1170), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1160), .B1(new_n782), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n941), .B2(new_n780), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1155), .B2(new_n773), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT121), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1159), .B1(new_n1180), .B2(new_n1181), .ZN(G378));
  INV_X1    g0982(.A(new_n1131), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1155), .B2(new_n1129), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n360), .A2(new_n363), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1185), .B(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n345), .A3(new_n905), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1185), .B(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n345), .A2(new_n905), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n964), .B2(G330), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n962), .A2(new_n963), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT38), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1196));
  OAI211_X1 g0996(.A(KEYINPUT40), .B(new_n958), .C1(new_n1196), .C2(new_n960), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1193), .A2(new_n1195), .A3(new_n1197), .A4(G330), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n952), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1195), .A2(new_n1197), .A3(G330), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1202), .A2(new_n944), .A3(new_n951), .A4(new_n1198), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1184), .A2(new_n1204), .A3(KEYINPUT57), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1204), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n722), .B(new_n1205), .C1(new_n1206), .C2(KEYINPUT125), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT125), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(KEYINPUT57), .C1(new_n1184), .C2(new_n1204), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1193), .A2(new_n780), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n776), .B1(G50), .B2(new_n841), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1024), .B1(new_n857), .B2(new_n582), .C1(new_n458), .C2(new_n807), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G41), .B(new_n604), .C1(G77), .C2(new_n812), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT122), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(KEYINPUT122), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G107), .A2(new_n846), .B1(new_n825), .B2(G283), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n814), .B2(new_n817), .C1(new_n467), .C2(new_n805), .ZN(new_n1219));
  OR4_X1    g1019(.A1(new_n1213), .A2(new_n1216), .A3(new_n1217), .A4(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n244), .B1(new_n405), .B2(new_n372), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1220), .A2(new_n1221), .B1(new_n293), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n853), .A2(G150), .B1(G125), .B2(new_n802), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT124), .ZN(new_n1225));
  INV_X1    g1025(.A(G128), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1226), .A2(new_n815), .B1(new_n811), .B2(new_n1164), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT123), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n847), .A2(G137), .B1(G132), .B2(new_n806), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n372), .B(new_n244), .C1(new_n817), .C2(new_n797), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G124), .B2(new_n825), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1223), .B1(new_n1221), .B2(new_n1220), .C1(new_n1231), .C2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1212), .B1(new_n1236), .B2(new_n782), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1204), .A2(new_n774), .B1(new_n1211), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1210), .A2(new_n1238), .ZN(G375));
  INV_X1    g1039(.A(new_n1129), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1183), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n992), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n949), .A2(new_n779), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n776), .B1(G68), .B2(new_n841), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n376), .B1(new_n817), .B2(new_n291), .C1(new_n857), .C2(new_n830), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G116), .B2(new_n806), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G107), .A2(new_n847), .B1(new_n825), .B2(G303), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G97), .A2(new_n812), .B1(new_n846), .B2(G283), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1248), .A2(new_n1065), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n811), .A2(new_n797), .B1(new_n796), .B2(new_n1226), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT127), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n805), .A2(new_n339), .B1(new_n793), .B2(new_n293), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT126), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n815), .A2(new_n858), .B1(new_n817), .B2(new_n814), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n405), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1165), .A2(new_n806), .B1(G132), .B2(new_n802), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1253), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n834), .B1(new_n1251), .B2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1246), .A2(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1240), .A2(new_n774), .B1(new_n1245), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1244), .A2(new_n1262), .ZN(G381));
  NAND3_X1  g1063(.A1(new_n1012), .A2(new_n1105), .A3(new_n1033), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1038), .A2(new_n839), .A3(new_n1072), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1264), .A2(G384), .A3(G381), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G375), .ZN(new_n1267));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(G407));
  NOR2_X1   g1069(.A1(new_n1266), .A2(new_n702), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1271));
  OAI21_X1  g1071(.A(G213), .B1(new_n1270), .B2(new_n1271), .ZN(G409));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  INV_X1    g1073(.A(G213), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G343), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1238), .C1(new_n1207), .C2(new_n1209), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1184), .A2(new_n1204), .A3(new_n1242), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1238), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1268), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1275), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1243), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1241), .A3(new_n722), .A4(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G384), .A3(new_n1262), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1286), .B2(new_n1262), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1282), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1287), .A3(new_n1281), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1273), .B1(new_n1280), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1275), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1296), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1265), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n839), .B1(new_n1038), .B2(new_n1072), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1012), .A2(new_n1105), .A3(new_n1033), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1105), .B1(new_n1012), .B2(new_n1033), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G387), .A2(G390), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1305), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1264), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1295), .A2(new_n1302), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1280), .A2(new_n1315), .A3(new_n1300), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1280), .B2(new_n1300), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1316), .A2(new_n1294), .A3(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1314), .B1(new_n1318), .B2(new_n1312), .ZN(G405));
  INV_X1    g1119(.A(new_n1312), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1268), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1301), .A3(new_n1276), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1301), .B1(new_n1321), .B2(new_n1276), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1320), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1324), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(new_n1312), .A3(new_n1322), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(G402));
endmodule


