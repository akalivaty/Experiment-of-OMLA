//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n224));
  AND4_X1   g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G238), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n210), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT1), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n215), .B1(new_n217), .B2(new_n220), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n231), .A2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G68), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n246), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT21), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n216), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI211_X1 g0060(.A(G257), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT78), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT78), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(G257), .A4(new_n258), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n259), .A2(new_n260), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n269), .A2(G264), .B1(new_n270), .B2(G303), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n257), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT75), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT5), .A2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT5), .A2(G41), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  OAI21_X1  g0081(.A(G274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n273), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n216), .B2(new_n256), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT5), .B(G41), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT75), .A4(new_n275), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n286), .A2(new_n275), .B1(new_n216), .B2(new_n256), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G270), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n272), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G283), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n293), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  INV_X1    g0096(.A(G116), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n294), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n296), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G116), .ZN(new_n305));
  INV_X1    g0105(.A(new_n304), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G1), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n306), .A2(new_n296), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n305), .B1(new_n309), .B2(G116), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n255), .B1(new_n292), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT80), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT80), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n255), .C1(new_n292), .C2(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n283), .A2(new_n287), .B1(new_n289), .B2(G270), .ZN(new_n318));
  OAI211_X1 g0118(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n319));
  INV_X1    g0119(.A(G303), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n265), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n267), .B2(new_n262), .ZN(new_n322));
  OAI211_X1 g0122(.A(G179), .B(new_n318), .C1(new_n322), .C2(new_n257), .ZN(new_n323));
  INV_X1    g0123(.A(new_n311), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n318), .B1(new_n322), .B2(new_n257), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n303), .B2(new_n310), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(KEYINPUT21), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT79), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n326), .A2(KEYINPUT79), .A3(new_n328), .A4(KEYINPUT21), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n325), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n311), .B1(new_n326), .B2(G200), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n326), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n317), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n307), .A2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G20), .A2(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G150), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n201), .B2(new_n209), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n296), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT68), .B(new_n296), .C1(new_n341), .C2(new_n344), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n304), .A2(G50), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n296), .B1(new_n208), .B2(G20), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(G50), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n347), .A2(KEYINPUT9), .A3(new_n348), .A4(new_n351), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n269), .A2(G223), .B1(new_n270), .B2(G77), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n265), .A2(G222), .A3(new_n258), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT67), .ZN(new_n359));
  INV_X1    g0159(.A(new_n257), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT67), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n361), .A3(new_n357), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G274), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n257), .A2(new_n364), .ZN(new_n367));
  INV_X1    g0167(.A(G226), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n354), .B(new_n355), .C1(new_n371), .C2(new_n335), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n257), .B1(new_n358), .B2(KEYINPUT67), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(new_n362), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n354), .A2(new_n355), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n371), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n374), .A2(G190), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n371), .A2(G179), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n352), .B1(new_n374), .B2(G169), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n339), .B1(G20), .B2(G77), .ZN(new_n390));
  INV_X1    g0190(.A(new_n338), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n342), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n390), .A2(new_n392), .B1(new_n281), .B2(new_n295), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n350), .A2(G77), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G77), .B2(new_n304), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G244), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n366), .B1(new_n367), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n269), .A2(G238), .B1(new_n270), .B2(G107), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n265), .A2(G232), .A3(new_n258), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n360), .ZN(new_n403));
  INV_X1    g0203(.A(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n397), .B(new_n405), .C1(G169), .C2(new_n403), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(G190), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n396), .C1(new_n375), .C2(new_n403), .ZN(new_n408));
  AND4_X1   g0208(.A1(new_n383), .A2(new_n387), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT69), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n342), .A2(G50), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT71), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n227), .A2(new_n209), .B1(new_n202), .B2(new_n340), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n296), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n227), .B2(new_n304), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n420), .A2(new_n422), .B1(new_n350), .B2(G68), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n367), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(G238), .B1(G274), .B2(new_n365), .ZN(new_n427));
  OAI211_X1 g0227(.A(G232), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n428));
  OAI211_X1 g0228(.A(G226), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT70), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n431), .A2(new_n432), .A3(new_n360), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n431), .B2(new_n360), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n427), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n427), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(G179), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n327), .B1(new_n436), .B2(new_n438), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI211_X1 g0242(.A(KEYINPUT14), .B(new_n327), .C1(new_n436), .C2(new_n438), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n425), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n436), .A2(new_n438), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G190), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n424), .C1(new_n375), .C2(new_n445), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n411), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n338), .A2(new_n304), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n350), .B2(new_n338), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n263), .A2(new_n209), .A3(new_n264), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT7), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT7), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n263), .A2(new_n453), .A3(new_n209), .A4(new_n264), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(G68), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G58), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n219), .B1(new_n226), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n342), .A2(G159), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n455), .A2(new_n458), .A3(KEYINPUT16), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n296), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n457), .A2(G20), .B1(G159), .B2(new_n342), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n227), .A3(new_n454), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT16), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n450), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n257), .A2(G232), .A3(new_n364), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n366), .ZN(new_n467));
  OR2_X1    g0267(.A1(G223), .A2(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n368), .A2(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G87), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n470), .A2(new_n270), .B1(new_n307), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n467), .A2(KEYINPUT73), .B1(new_n472), .B2(new_n360), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT73), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n466), .A2(new_n366), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(G179), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n467), .A2(KEYINPUT73), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n360), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n477), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(new_n327), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n465), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT18), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT18), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n465), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n375), .B1(new_n473), .B2(new_n475), .ZN(new_n487));
  AND4_X1   g0287(.A1(G190), .A2(new_n477), .A3(new_n478), .A4(new_n475), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n462), .A2(new_n463), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT16), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n296), .A3(new_n460), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n489), .A2(KEYINPUT17), .A3(new_n493), .A4(new_n450), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT17), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n473), .A2(G190), .A3(new_n475), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n479), .B2(new_n375), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n465), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n486), .B(new_n499), .C1(new_n409), .C2(new_n410), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n448), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n452), .A2(G107), .A3(new_n454), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n342), .A2(G77), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n204), .A3(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n504), .B1(new_n508), .B2(new_n209), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n296), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n304), .A2(G97), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n309), .B2(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G250), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT74), .ZN(new_n515));
  OAI211_X1 g0315(.A(G244), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(new_n293), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n360), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n283), .A2(new_n287), .B1(new_n289), .B2(G257), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(G179), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n327), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n513), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n209), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n265), .A2(new_n528), .A3(new_n209), .A4(G87), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n209), .A2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n531), .A2(new_n532), .B1(G20), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT81), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n531), .A2(new_n537), .A3(new_n532), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n530), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n530), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n296), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XOR2_X1   g0343(.A(KEYINPUT82), .B(KEYINPUT25), .Z(new_n544));
  NOR2_X1   g0344(.A1(new_n304), .A2(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(G107), .B2(new_n309), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n265), .A2(G250), .A3(new_n258), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G294), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n360), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n289), .A2(G264), .ZN(new_n553));
  AND4_X1   g0353(.A1(new_n335), .A2(new_n552), .A3(new_n288), .A4(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n551), .A2(new_n360), .B1(G264), .B2(new_n289), .ZN(new_n555));
  AOI21_X1  g0355(.A(G200), .B1(new_n555), .B2(new_n288), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n543), .B(new_n547), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n521), .A2(G190), .A3(new_n522), .ZN(new_n558));
  INV_X1    g0358(.A(new_n512), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n502), .B(new_n504), .C1(new_n209), .C2(new_n508), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n296), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n289), .A2(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n288), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n516), .A2(new_n517), .B1(G33), .B2(G283), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT74), .B1(new_n269), .B2(G250), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT74), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n514), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n519), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n563), .B1(new_n360), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n558), .B(new_n561), .C1(new_n569), .C2(new_n375), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n525), .A2(new_n557), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n573));
  OAI211_X1 g0373(.A(G238), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n533), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT76), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT76), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n573), .A2(new_n574), .A3(new_n577), .A4(new_n533), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n360), .ZN(new_n580));
  INV_X1    g0380(.A(new_n275), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G250), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n582), .A2(new_n360), .B1(new_n284), .B2(new_n581), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n404), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n257), .B1(new_n576), .B2(new_n578), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n583), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT77), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n404), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n340), .B2(new_n204), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n265), .A2(new_n209), .A3(G68), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n209), .B1(new_n430), .B2(new_n591), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G87), .B2(new_n206), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n296), .B1(new_n306), .B2(new_n388), .ZN(new_n597));
  INV_X1    g0397(.A(new_n309), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n388), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n327), .B1(new_n587), .B2(new_n583), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n586), .A2(new_n590), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n543), .A2(new_n547), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n555), .A2(new_n404), .A3(new_n288), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n555), .A2(new_n288), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n327), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n580), .A2(G190), .A3(new_n584), .ZN(new_n607));
  OAI21_X1  g0407(.A(G200), .B1(new_n587), .B2(new_n583), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n309), .A2(G87), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n597), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n601), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n337), .A2(new_n501), .A3(new_n572), .A4(new_n612), .ZN(G372));
  NAND2_X1  g0413(.A1(new_n521), .A2(new_n522), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n513), .B1(G200), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n521), .A2(G179), .A3(new_n522), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n569), .B2(new_n327), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n615), .A2(new_n558), .B1(new_n617), .B2(new_n513), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n585), .A2(new_n599), .A3(new_n600), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n618), .A2(new_n620), .A3(KEYINPUT83), .A4(new_n557), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n611), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n571), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n317), .A2(new_n333), .A3(new_n606), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(KEYINPUT84), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT84), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n616), .B(new_n628), .C1(new_n569), .C2(new_n327), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n513), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n627), .A2(KEYINPUT85), .A3(new_n629), .A4(new_n513), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n620), .A4(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n619), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n601), .A2(new_n513), .A3(new_n617), .A4(new_n611), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n626), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n501), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n447), .A2(new_n499), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n406), .B2(new_n444), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n383), .B1(new_n642), .B2(new_n485), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n387), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(G369));
  NAND3_X1  g0445(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n317), .B2(new_n333), .ZN(new_n652));
  INV_X1    g0452(.A(new_n557), .ZN(new_n653));
  INV_X1    g0453(.A(new_n651), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n543), .B2(new_n547), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n606), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n606), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n652), .A2(new_n656), .B1(new_n657), .B2(new_n654), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n317), .A2(new_n333), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n311), .A2(new_n651), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT86), .Z(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n337), .A2(KEYINPUT87), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(new_n661), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n337), .A2(KEYINPUT87), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n657), .A2(new_n654), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n656), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(G330), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT88), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n666), .A2(new_n672), .A3(G330), .A4(new_n668), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n658), .B1(new_n671), .B2(new_n674), .ZN(G399));
  NOR2_X1   g0475(.A1(new_n212), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n220), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(new_n555), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n323), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n569), .A4(new_n588), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n580), .A2(new_n521), .A3(new_n522), .A4(new_n584), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n268), .A2(new_n271), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n360), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(G179), .A3(new_n555), .A4(new_n318), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n685), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(G179), .B1(new_n688), .B2(new_n318), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n580), .A2(new_n584), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n614), .A4(new_n604), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n684), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n694), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT31), .B1(new_n694), .B2(new_n651), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n337), .A2(new_n572), .A3(new_n612), .A4(new_n654), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n639), .A2(new_n654), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n632), .A2(KEYINPUT26), .A3(new_n620), .A4(new_n634), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n637), .A2(new_n633), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(KEYINPUT89), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n571), .A2(new_n623), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n636), .B1(new_n707), .B2(new_n625), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n704), .B2(KEYINPUT89), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT29), .B(new_n654), .C1(new_n706), .C2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n701), .B1(new_n703), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n681), .B1(new_n711), .B2(G1), .ZN(G364));
  AOI21_X1  g0512(.A(new_n281), .B1(G20), .B2(new_n327), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n209), .A2(G190), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G179), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT92), .Z(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G329), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n209), .A2(new_n335), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n375), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n404), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(G303), .A2(new_n722), .B1(new_n725), .B2(G311), .ZN(new_n726));
  INV_X1    g0526(.A(G283), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n714), .A2(new_n720), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n718), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n209), .B1(new_n715), .B2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(G294), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n719), .A2(new_n723), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n270), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n404), .A2(new_n375), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n714), .ZN(new_n737));
  XOR2_X1   g0537(.A(KEYINPUT33), .B(G317), .Z(new_n738));
  NAND2_X1  g0538(.A1(new_n719), .A2(new_n736), .ZN(new_n739));
  INV_X1    g0539(.A(G326), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n729), .A2(new_n732), .A3(new_n735), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT93), .Z(new_n743));
  XNOR2_X1  g0543(.A(new_n730), .B(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G97), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n739), .A2(new_n247), .B1(new_n737), .B2(new_n249), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(G87), .B2(new_n722), .ZN(new_n747));
  INV_X1    g0547(.A(G159), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n716), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT32), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n733), .A2(new_n456), .B1(new_n724), .B2(new_n202), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n728), .A2(new_n205), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n751), .A2(new_n270), .A3(new_n752), .ZN(new_n753));
  AND4_X1   g0553(.A1(new_n745), .A2(new_n747), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n713), .B1(new_n743), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n211), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n208), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n676), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n713), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT90), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(new_n270), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n297), .B2(new_n212), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n253), .A2(new_n274), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n212), .A2(new_n265), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G45), .B2(new_n220), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n760), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n763), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n755), .B(new_n773), .C1(new_n666), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n666), .A2(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n760), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n666), .A2(G330), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n397), .A2(new_n651), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n406), .A2(new_n408), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT95), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n406), .A2(new_n408), .A3(new_n783), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n639), .A2(new_n654), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n406), .A2(new_n654), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n782), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n702), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n759), .B1(new_n790), .B2(new_n700), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n700), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n713), .A2(new_n761), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n759), .B1(G77), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n733), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G143), .A2(new_n796), .B1(new_n725), .B2(G159), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  INV_X1    g0598(.A(G150), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n739), .C1(new_n799), .C2(new_n737), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT34), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n728), .A2(new_n249), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n265), .B1(new_n721), .B2(new_n247), .ZN(new_n803));
  INV_X1    g0603(.A(new_n730), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n802), .B(new_n803), .C1(G58), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  INV_X1    g0606(.A(new_n717), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT94), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n727), .A2(new_n737), .B1(new_n733), .B2(new_n731), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n739), .A2(new_n320), .B1(new_n724), .B2(new_n297), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n270), .B1(new_n721), .B2(new_n205), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n728), .A2(new_n471), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n745), .C1(new_n816), .C2(new_n807), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n809), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n810), .B2(new_n817), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n795), .B1(new_n819), .B2(new_n713), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n789), .B2(new_n762), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n792), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  NAND3_X1  g0623(.A1(new_n703), .A2(new_n501), .A3(new_n710), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n644), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n406), .A2(new_n651), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n786), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n482), .A2(new_n484), .A3(new_n494), .A4(new_n498), .ZN(new_n830));
  INV_X1    g0630(.A(new_n649), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT16), .B1(new_n462), .B2(new_n455), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n450), .B1(new_n461), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n487), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n493), .A2(new_n835), .A3(new_n450), .A4(new_n496), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n465), .A2(new_n831), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n836), .A2(new_n481), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n465), .A2(new_n497), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n480), .A2(new_n831), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n833), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n839), .B1(new_n842), .B2(new_n838), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n834), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n834), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n425), .A2(new_n651), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n444), .A2(new_n447), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n425), .B(new_n651), .C1(new_n442), .C2(new_n443), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n829), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT98), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n486), .A2(new_n831), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n837), .B2(KEYINPUT99), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n836), .A2(new_n481), .A3(new_n837), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n830), .A2(new_n465), .A3(new_n831), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n834), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n846), .A2(KEYINPUT39), .A3(new_n847), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n444), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n654), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n857), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n854), .B1(new_n853), .B2(new_n856), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n826), .B(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n501), .A2(new_n699), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n788), .B1(new_n850), .B2(new_n851), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n877), .B(new_n699), .C1(new_n863), .C2(new_n864), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT40), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n877), .A2(new_n699), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT40), .B1(new_n846), .B2(new_n847), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n876), .A2(new_n883), .ZN(new_n885));
  INV_X1    g0685(.A(G330), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n875), .A2(new_n887), .B1(new_n208), .B2(new_n756), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n875), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n217), .A2(new_n297), .ZN(new_n890));
  INV_X1    g0690(.A(new_n508), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(KEYINPUT35), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT96), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(KEYINPUT35), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT36), .Z(new_n898));
  INV_X1    g0698(.A(new_n220), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n899), .B(G77), .C1(new_n456), .C2(new_n226), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n208), .B(G13), .C1(new_n900), .C2(new_n248), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n889), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT101), .ZN(G367));
  INV_X1    g0703(.A(new_n770), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n764), .B1(new_n213), .B2(new_n388), .C1(new_n242), .C2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n759), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n610), .A2(new_n654), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n636), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n623), .B2(new_n907), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n270), .B1(new_n722), .B2(G58), .ZN(new_n910));
  INV_X1    g0710(.A(G143), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n910), .B1(new_n911), .B2(new_n739), .C1(new_n748), .C2(new_n737), .ZN(new_n912));
  INV_X1    g0712(.A(new_n744), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n249), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n724), .A2(new_n247), .B1(new_n716), .B2(new_n798), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n733), .A2(new_n799), .B1(new_n728), .B2(new_n202), .ZN(new_n916));
  NOR4_X1   g0716(.A1(new_n912), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G303), .A2(new_n796), .B1(new_n725), .B2(G283), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n731), .B2(new_n737), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n722), .A2(KEYINPUT46), .A3(G116), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT46), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n721), .B2(new_n297), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(new_n922), .C1(new_n205), .C2(new_n730), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n270), .B1(new_n739), .B2(new_n816), .ZN(new_n924));
  INV_X1    g0724(.A(G317), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n728), .A2(new_n204), .B1(new_n716), .B2(new_n925), .ZN(new_n926));
  NOR4_X1   g0726(.A1(new_n919), .A2(new_n923), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n917), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT47), .ZN(new_n929));
  INV_X1    g0729(.A(new_n713), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n906), .B1(new_n909), .B2(new_n774), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n676), .B(KEYINPUT41), .Z(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n670), .A2(new_n933), .A3(new_n673), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT44), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n630), .A2(new_n654), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n618), .B1(new_n561), .B2(new_n654), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n935), .B1(new_n939), .B2(new_n658), .ZN(new_n940));
  INV_X1    g0740(.A(new_n658), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n938), .A3(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n658), .A3(KEYINPUT45), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n941), .B2(new_n938), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n934), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n668), .B(new_n652), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n776), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n670), .A2(new_n933), .A3(new_n673), .A4(new_n948), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n932), .B1(new_n954), .B2(new_n711), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n758), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n671), .A2(new_n674), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n939), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n525), .B1(new_n938), .B2(new_n606), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n654), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n668), .A2(new_n652), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n938), .A2(new_n961), .A3(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT42), .B1(new_n938), .B2(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n909), .B(KEYINPUT43), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n960), .A2(new_n962), .A3(new_n963), .A4(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n968), .A2(KEYINPUT102), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(KEYINPUT102), .ZN(new_n970));
  OAI211_X1 g0770(.A(KEYINPUT103), .B(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n962), .A2(new_n963), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT102), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n973), .A2(new_n974), .A3(new_n960), .A4(new_n967), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n968), .A2(KEYINPUT102), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT103), .B1(new_n977), .B2(new_n966), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n958), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT103), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n982), .A2(new_n957), .A3(new_n939), .A4(new_n971), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n931), .B1(new_n956), .B2(new_n984), .ZN(G387));
  AOI21_X1  g0785(.A(new_n677), .B1(new_n952), .B2(new_n711), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n711), .B2(new_n952), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n952), .A2(new_n758), .ZN(new_n988));
  INV_X1    g0788(.A(new_n678), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n767), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(G107), .B2(new_n213), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n239), .A2(new_n274), .ZN(new_n992));
  AOI211_X1 g0792(.A(G45), .B(new_n989), .C1(G68), .C2(G77), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n338), .A2(G50), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT50), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n904), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n991), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n759), .B1(new_n997), .B2(new_n765), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n744), .A2(new_n389), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n247), .A2(new_n733), .B1(new_n737), .B2(new_n338), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n721), .A2(new_n202), .B1(new_n716), .B2(new_n799), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n728), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n270), .B1(new_n1003), .B2(G97), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n739), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1005), .A2(G159), .B1(new_n725), .B2(G68), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n999), .A2(new_n1002), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n739), .A2(new_n734), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n733), .A2(new_n925), .B1(new_n724), .B2(new_n320), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n737), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1009), .C1(G311), .C2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT48), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT48), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n722), .A2(G294), .B1(new_n804), .B2(G283), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT49), .Z(new_n1016));
  OAI221_X1 g0816(.A(new_n270), .B1(new_n716), .B2(new_n740), .C1(new_n297), .C2(new_n728), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n998), .B1(new_n1018), .B2(new_n713), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n668), .B2(new_n774), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n987), .A2(new_n988), .A3(new_n1020), .ZN(G393));
  AOI21_X1  g0821(.A(new_n677), .B1(new_n950), .B2(new_n953), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n711), .A3(new_n952), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n957), .A2(new_n948), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n949), .B1(new_n671), .B2(new_n674), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n986), .C2(new_n758), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n764), .B1(new_n204), .B2(new_n213), .C1(new_n246), .C2(new_n904), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n759), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n739), .A2(new_n799), .B1(new_n733), .B2(new_n748), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n721), .A2(new_n226), .B1(new_n724), .B2(new_n338), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n737), .A2(new_n247), .B1(new_n716), .B2(new_n911), .ZN(new_n1032));
  NOR4_X1   g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n270), .A4(new_n814), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n744), .A2(G77), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n739), .A2(new_n925), .B1(new_n733), .B2(new_n816), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  AOI211_X1 g0837(.A(new_n265), .B(new_n752), .C1(G116), .C2(new_n804), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G303), .A2(new_n1010), .B1(new_n725), .B2(G294), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n716), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G283), .A2(new_n722), .B1(new_n1040), .B2(G322), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1035), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1028), .B1(new_n1043), .B2(new_n713), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n939), .B2(new_n774), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1023), .A2(new_n1026), .A3(new_n1045), .ZN(G390));
  OAI21_X1  g0846(.A(new_n759), .B1(new_n391), .B2(new_n794), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n802), .B1(new_n717), .B2(G294), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT107), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n265), .B1(new_n722), .B2(G87), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n739), .A2(new_n727), .B1(new_n737), .B2(new_n205), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n733), .A2(new_n297), .B1(new_n724), .B2(new_n204), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1034), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT108), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G132), .A2(new_n796), .B1(new_n1003), .B2(G50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n270), .B1(new_n1005), .B2(G128), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n798), .C2(new_n737), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G159), .B2(new_n744), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n717), .A2(G125), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n721), .A2(new_n799), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT53), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT54), .B(G143), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT106), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n725), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT109), .B1(new_n1055), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(new_n930), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1055), .A2(KEYINPUT109), .A3(new_n1066), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1047), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n867), .B2(new_n762), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n701), .A2(new_n877), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n829), .A2(new_n852), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n867), .B1(new_n1074), .B2(new_n869), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n869), .B1(new_n863), .B2(new_n864), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n654), .B(new_n785), .C1(new_n706), .C2(new_n709), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n827), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1078), .B2(new_n852), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n865), .A2(new_n866), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n852), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n786), .B2(new_n828), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1083), .B2(new_n870), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1082), .B1(new_n1077), .B2(new_n827), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1072), .C1(new_n1085), .C2(new_n1076), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1071), .B1(new_n1087), .B2(new_n757), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n448), .A2(new_n700), .A3(new_n500), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n825), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1082), .B1(new_n700), .B2(new_n788), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1072), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n829), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1078), .B2(new_n1092), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT105), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(new_n1087), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n677), .B1(new_n1095), .B2(new_n1087), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1088), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(G378));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT115), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n352), .A2(new_n831), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n383), .B2(new_n387), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n383), .A2(new_n387), .A3(new_n1103), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1102), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1103), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1108), .B(new_n386), .C1(new_n377), .C2(new_n382), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1102), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1104), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1101), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1105), .A2(new_n1106), .A3(new_n1102), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1110), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(KEYINPUT115), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n883), .A2(new_n1100), .A3(new_n1116), .A4(G330), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(KEYINPUT40), .A2(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n886), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n886), .B1(new_n879), .B2(new_n882), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1100), .B1(new_n1122), .B2(new_n1116), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n874), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  AOI221_X4 g0925(.A(new_n1082), .B1(new_n847), .B2(new_n846), .C1(new_n786), .C2(new_n828), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT98), .B1(new_n1126), .B2(new_n855), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n857), .A3(new_n871), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n1123), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1080), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1125), .A2(new_n1130), .B1(new_n1090), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT117), .B1(new_n1132), .B2(KEYINPUT57), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n677), .B1(new_n1132), .B2(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1090), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n872), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1121), .A2(new_n1124), .B1(new_n1136), .B2(new_n1127), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1128), .A2(new_n1129), .A3(new_n1123), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1133), .A2(new_n1134), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n758), .ZN(new_n1145));
  AOI211_X1 g0945(.A(G33), .B(G41), .C1(new_n1040), .C2(G124), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n744), .A2(G150), .B1(G125), .B2(new_n1005), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT113), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n1064), .A2(new_n722), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT112), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(KEYINPUT112), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n733), .A2(new_n1152), .B1(new_n724), .B2(new_n798), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G132), .B2(new_n1010), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .A4(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n1156));
  OAI221_X1 g0956(.A(new_n1146), .B1(new_n748), .B2(new_n728), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n247), .B1(new_n259), .B2(G41), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n733), .A2(new_n205), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT110), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n807), .B2(new_n727), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G41), .B(new_n265), .C1(new_n722), .C2(G77), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G116), .A2(new_n1005), .B1(new_n1010), .B2(G97), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1003), .A2(G58), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n725), .A2(new_n389), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1162), .A2(new_n914), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1159), .B1(new_n1168), .B2(KEYINPUT58), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(KEYINPUT111), .B1(KEYINPUT58), .B2(new_n1168), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(KEYINPUT111), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n713), .B1(new_n1158), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n760), .B1(new_n247), .B2(new_n793), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n1116), .C2(new_n762), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1145), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1143), .A2(new_n1176), .ZN(G375));
  NAND2_X1  g0977(.A1(new_n1094), .A2(new_n758), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n760), .B1(new_n249), .B2(new_n793), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n204), .A2(new_n721), .B1(new_n737), .B2(new_n297), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n265), .B(new_n1180), .C1(G77), .C2(new_n1003), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n717), .A2(G303), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n739), .A2(new_n731), .B1(new_n724), .B2(new_n205), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G283), .B2(new_n796), .ZN(new_n1184));
  AND4_X1   g0984(.A1(new_n999), .A2(new_n1181), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1165), .A2(new_n265), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT118), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n721), .A2(new_n748), .B1(new_n724), .B2(new_n799), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n717), .B2(G128), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n247), .C2(new_n913), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT119), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n739), .A2(new_n806), .B1(new_n733), .B2(new_n798), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1064), .B2(new_n1010), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1185), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1179), .B1(new_n930), .B2(new_n1194), .C1(new_n852), .C2(new_n762), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1178), .A2(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n932), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(G381));
  NAND3_X1  g1001(.A1(new_n1143), .A2(new_n1098), .A3(new_n1176), .ZN(new_n1202));
  INV_X1    g1002(.A(G390), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1203), .A2(new_n1200), .A3(new_n822), .A4(new_n1204), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1202), .A2(G387), .A3(new_n1205), .ZN(G407));
  AND2_X1   g1006(.A1(G407), .A2(G213), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n650), .A2(G213), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT120), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT121), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT121), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1207), .B(new_n1215), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(G409));
  INV_X1    g1017(.A(new_n932), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1144), .A2(new_n1218), .A3(new_n1135), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1098), .B1(new_n1175), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT122), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT122), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1098), .B(new_n1222), .C1(new_n1175), .C2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1143), .A2(G378), .A3(new_n1176), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1208), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1199), .B1(new_n1197), .B2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1090), .A2(new_n1094), .A3(new_n1227), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n677), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1196), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(new_n822), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n650), .A2(G213), .A3(G2897), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT124), .Z(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1231), .B(G384), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1226), .B2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1221), .B(new_n1223), .C1(G375), .C2(new_n1098), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT62), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1208), .A4(new_n1232), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1208), .B(new_n1232), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT62), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1203), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G390), .B(new_n931), .C1(new_n956), .C2(new_n984), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G393), .B(G396), .ZN(new_n1250));
  AND4_X1   g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(KEYINPUT125), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1252), .A2(new_n1250), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1246), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1244), .B2(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1244), .A2(new_n1258), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1226), .A2(KEYINPUT123), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1239), .B1(new_n1226), .B2(KEYINPUT123), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1259), .B(new_n1260), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1263), .ZN(G405));
  AND3_X1   g1064(.A1(new_n1143), .A2(new_n1098), .A3(new_n1176), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1098), .B1(new_n1143), .B2(new_n1176), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1236), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1236), .B(KEYINPUT127), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n1202), .A3(new_n1232), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1232), .A4(new_n1202), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1271), .A2(new_n1277), .A3(new_n1254), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1254), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G402));
endmodule


