

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770;

  XOR2_X1 U386 ( .A(G137), .B(G140), .Z(n537) );
  AND2_X4 U387 ( .A1(n647), .A2(n468), .ZN(n425) );
  XNOR2_X2 U388 ( .A(n527), .B(G469), .ZN(n614) );
  NOR2_X1 U389 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U390 ( .A1(n682), .A2(n646), .ZN(n468) );
  XNOR2_X1 U391 ( .A(n760), .B(KEYINPUT72), .ZN(n426) );
  NOR2_X1 U392 ( .A1(n770), .A2(n580), .ZN(n581) );
  XNOR2_X1 U393 ( .A(n431), .B(n430), .ZN(n769) );
  XNOR2_X1 U394 ( .A(n379), .B(n460), .ZN(n766) );
  XNOR2_X1 U395 ( .A(n458), .B(KEYINPUT101), .ZN(n670) );
  NOR2_X1 U396 ( .A1(n614), .A2(n692), .ZN(n594) );
  NOR2_X1 U397 ( .A1(n596), .A2(n410), .ZN(n409) );
  AND2_X1 U398 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U399 ( .A(n368), .B(n476), .ZN(n531) );
  INV_X2 U400 ( .A(G125), .ZN(n414) );
  XNOR2_X1 U401 ( .A(n724), .B(n725), .ZN(n726) );
  NAND2_X1 U402 ( .A1(n629), .A2(n705), .ZN(n623) );
  NAND2_X1 U403 ( .A1(n365), .A2(n384), .ZN(n383) );
  XNOR2_X1 U404 ( .A(n634), .B(KEYINPUT77), .ZN(n384) );
  XNOR2_X1 U405 ( .A(n522), .B(n521), .ZN(n532) );
  XNOR2_X1 U406 ( .A(G131), .B(G134), .ZN(n521) );
  XNOR2_X1 U407 ( .A(n532), .B(n537), .ZN(n752) );
  XNOR2_X1 U408 ( .A(n595), .B(n373), .ZN(n636) );
  NOR2_X1 U409 ( .A1(n622), .A2(n623), .ZN(n420) );
  INV_X1 U410 ( .A(n569), .ZN(n403) );
  INV_X1 U411 ( .A(n555), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n429), .B(n428), .ZN(n639) );
  INV_X1 U413 ( .A(KEYINPUT46), .ZN(n428) );
  NOR2_X1 U414 ( .A1(n766), .A2(n769), .ZN(n429) );
  XNOR2_X1 U415 ( .A(n673), .B(n408), .ZN(n380) );
  INV_X1 U416 ( .A(n679), .ZN(n454) );
  NAND2_X1 U417 ( .A1(n639), .A2(KEYINPUT48), .ZN(n450) );
  XNOR2_X1 U418 ( .A(G143), .B(G131), .ZN(n508) );
  XNOR2_X1 U419 ( .A(G101), .B(KEYINPUT3), .ZN(n476) );
  XNOR2_X1 U420 ( .A(n456), .B(G104), .ZN(n507) );
  INV_X1 U421 ( .A(G122), .ZN(n456) );
  NOR2_X1 U422 ( .A1(n709), .A2(n708), .ZN(n637) );
  INV_X1 U423 ( .A(KEYINPUT0), .ZN(n436) );
  NAND2_X1 U424 ( .A1(n610), .A2(n487), .ZN(n437) );
  NAND2_X2 U425 ( .A1(n394), .A2(n392), .ZN(n629) );
  NAND2_X1 U426 ( .A1(n485), .A2(n488), .ZN(n393) );
  AND2_X1 U427 ( .A1(n386), .A2(n593), .ZN(n632) );
  AND2_X1 U428 ( .A1(n594), .A2(n387), .ZN(n386) );
  INV_X1 U429 ( .A(KEYINPUT30), .ZN(n591) );
  XOR2_X1 U430 ( .A(n514), .B(n513), .Z(n572) );
  INV_X1 U431 ( .A(KEYINPUT121), .ZN(n463) );
  NAND2_X1 U432 ( .A1(n413), .A2(n641), .ZN(n647) );
  XNOR2_X1 U433 ( .A(n752), .B(n465), .ZN(n731) );
  XNOR2_X1 U434 ( .A(n526), .B(n523), .ZN(n465) );
  XNOR2_X1 U435 ( .A(n525), .B(n375), .ZN(n526) );
  NOR2_X1 U436 ( .A1(n761), .A2(G952), .ZN(n740) );
  INV_X1 U437 ( .A(KEYINPUT83), .ZN(n408) );
  NAND2_X1 U438 ( .A1(n404), .A2(n401), .ZN(n400) );
  NAND2_X1 U439 ( .A1(n399), .A2(n367), .ZN(n398) );
  OR2_X1 U440 ( .A1(G237), .A2(G902), .ZN(n486) );
  INV_X1 U441 ( .A(n689), .ZN(n410) );
  XNOR2_X1 U442 ( .A(G128), .B(G119), .ZN(n538) );
  XNOR2_X1 U443 ( .A(G110), .B(KEYINPUT97), .ZN(n539) );
  XOR2_X1 U444 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n498) );
  XOR2_X1 U445 ( .A(KEYINPUT69), .B(G110), .Z(n524) );
  NOR2_X1 U446 ( .A1(n451), .A2(n449), .ZN(n644) );
  NAND2_X1 U447 ( .A1(n450), .A2(n454), .ZN(n449) );
  NOR2_X2 U448 ( .A1(n670), .A2(n668), .ZN(n710) );
  NAND2_X1 U449 ( .A1(n706), .A2(n705), .ZN(n709) );
  XNOR2_X1 U450 ( .A(n629), .B(n427), .ZN(n706) );
  INV_X1 U451 ( .A(KEYINPUT38), .ZN(n427) );
  XNOR2_X1 U452 ( .A(n556), .B(n377), .ZN(n577) );
  INV_X1 U453 ( .A(KEYINPUT71), .ZN(n377) );
  NAND2_X1 U454 ( .A1(n397), .A2(n646), .ZN(n395) );
  INV_X1 U455 ( .A(n596), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n467), .B(n529), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n531), .B(n366), .ZN(n390) );
  XNOR2_X1 U459 ( .A(G953), .B(KEYINPUT64), .ZN(n587) );
  AND2_X2 U460 ( .A1(n644), .A2(n677), .ZN(n760) );
  XNOR2_X1 U461 ( .A(n418), .B(G128), .ZN(n492) );
  INV_X1 U462 ( .A(G143), .ZN(n418) );
  XNOR2_X1 U463 ( .A(G134), .B(G122), .ZN(n494) );
  XNOR2_X1 U464 ( .A(n457), .B(n455), .ZN(n512) );
  XNOR2_X1 U465 ( .A(n507), .B(n508), .ZN(n455) );
  XNOR2_X1 U466 ( .A(n511), .B(n370), .ZN(n457) );
  XNOR2_X1 U467 ( .A(n524), .B(n376), .ZN(n375) );
  INV_X1 U468 ( .A(KEYINPUT96), .ZN(n376) );
  XOR2_X1 U469 ( .A(G107), .B(G104), .Z(n520) );
  XNOR2_X1 U470 ( .A(G101), .B(G146), .ZN(n519) );
  XNOR2_X1 U471 ( .A(n492), .B(n417), .ZN(n522) );
  INV_X1 U472 ( .A(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n479), .B(n412), .ZN(n481) );
  XNOR2_X1 U474 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n479) );
  XNOR2_X1 U475 ( .A(KEYINPUT89), .B(KEYINPUT91), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n477), .B(n478), .ZN(n741) );
  INV_X1 U477 ( .A(KEYINPUT80), .ZN(n416) );
  NAND2_X1 U478 ( .A1(G234), .A2(G237), .ZN(n469) );
  INV_X1 U479 ( .A(KEYINPUT35), .ZN(n432) );
  INV_X1 U480 ( .A(KEYINPUT22), .ZN(n517) );
  INV_X1 U481 ( .A(KEYINPUT95), .ZN(n435) );
  INV_X1 U482 ( .A(KEYINPUT124), .ZN(n440) );
  INV_X1 U483 ( .A(G953), .ZN(n757) );
  INV_X1 U484 ( .A(KEYINPUT42), .ZN(n430) );
  OR2_X1 U485 ( .A1(n704), .A2(n638), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n461), .B(KEYINPUT110), .ZN(n460) );
  NAND2_X1 U487 ( .A1(n636), .A2(n668), .ZN(n379) );
  INV_X1 U488 ( .A(KEYINPUT40), .ZN(n461) );
  NAND2_X1 U489 ( .A1(n381), .A2(n625), .ZN(n673) );
  XNOR2_X1 U490 ( .A(n420), .B(n466), .ZN(n381) );
  XNOR2_X1 U491 ( .A(n385), .B(KEYINPUT108), .ZN(n768) );
  NAND2_X1 U492 ( .A1(n632), .A2(n631), .ZN(n385) );
  XNOR2_X1 U493 ( .A(n441), .B(n438), .ZN(G69) );
  XNOR2_X1 U494 ( .A(n751), .B(n439), .ZN(n438) );
  NAND2_X1 U495 ( .A1(n750), .A2(n749), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n440), .B(KEYINPUT125), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n464), .B(n462), .ZN(n739) );
  XNOR2_X1 U498 ( .A(n738), .B(n463), .ZN(n462) );
  INV_X1 U499 ( .A(KEYINPUT60), .ZN(n442) );
  INV_X1 U500 ( .A(n740), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n729), .B(n421), .ZN(n732) );
  XNOR2_X1 U502 ( .A(n731), .B(n730), .ZN(n421) );
  XNOR2_X1 U503 ( .A(G902), .B(KEYINPUT15), .ZN(n488) );
  AND2_X1 U504 ( .A1(n620), .A2(n619), .ZN(n365) );
  XNOR2_X1 U505 ( .A(G146), .B(G116), .ZN(n366) );
  AND2_X1 U506 ( .A1(n767), .A2(n405), .ZN(n367) );
  XOR2_X1 U507 ( .A(G113), .B(G119), .Z(n368) );
  AND2_X1 U508 ( .A1(n406), .A2(n400), .ZN(n369) );
  XNOR2_X1 U509 ( .A(n584), .B(n583), .ZN(n683) );
  INV_X1 U510 ( .A(n485), .ZN(n397) );
  AND2_X1 U511 ( .A1(G214), .A2(n530), .ZN(n370) );
  AND2_X1 U512 ( .A1(n569), .A2(n555), .ZN(n371) );
  AND2_X1 U513 ( .A1(n682), .A2(n681), .ZN(n372) );
  XNOR2_X1 U514 ( .A(KEYINPUT39), .B(KEYINPUT84), .ZN(n373) );
  XNOR2_X1 U515 ( .A(n422), .B(n741), .ZN(n724) );
  XOR2_X1 U516 ( .A(n734), .B(n733), .Z(n374) );
  NAND2_X1 U517 ( .A1(n369), .A2(n398), .ZN(n562) );
  NAND2_X1 U518 ( .A1(n645), .A2(n644), .ZN(n682) );
  NOR2_X1 U519 ( .A1(n383), .A2(n635), .ZN(n382) );
  NAND2_X1 U520 ( .A1(n577), .A2(n557), .ZN(n558) );
  NAND2_X1 U521 ( .A1(n565), .A2(n378), .ZN(n582) );
  NAND2_X1 U522 ( .A1(n765), .A2(n564), .ZN(n378) );
  XNOR2_X2 U523 ( .A(n614), .B(KEYINPUT1), .ZN(n691) );
  XNOR2_X1 U524 ( .A(n433), .B(n432), .ZN(n563) );
  NOR2_X1 U525 ( .A1(n714), .A2(n560), .ZN(n561) );
  NAND2_X1 U526 ( .A1(n382), .A2(n380), .ZN(n640) );
  XNOR2_X1 U527 ( .A(n532), .B(n388), .ZN(n648) );
  NAND2_X1 U528 ( .A1(n391), .A2(n516), .ZN(n518) );
  XNOR2_X1 U529 ( .A(n391), .B(n435), .ZN(n575) );
  NAND2_X1 U530 ( .A1(n701), .A2(n391), .ZN(n578) );
  XNOR2_X2 U531 ( .A(n437), .B(n436), .ZN(n391) );
  OR2_X1 U532 ( .A1(n724), .A2(n393), .ZN(n392) );
  NAND2_X1 U533 ( .A1(n724), .A2(n397), .ZN(n396) );
  XNOR2_X2 U534 ( .A(n623), .B(KEYINPUT19), .ZN(n610) );
  NAND2_X1 U535 ( .A1(n407), .A2(n371), .ZN(n406) );
  XNOR2_X2 U536 ( .A(n535), .B(KEYINPUT65), .ZN(n407) );
  NAND2_X1 U537 ( .A1(n407), .A2(n569), .ZN(n663) );
  INV_X1 U538 ( .A(n407), .ZN(n399) );
  NAND2_X1 U539 ( .A1(n767), .A2(n402), .ZN(n401) );
  NAND2_X1 U540 ( .A1(n403), .A2(n405), .ZN(n402) );
  OR2_X1 U541 ( .A1(n767), .A2(n555), .ZN(n404) );
  NAND2_X1 U542 ( .A1(n425), .A2(G210), .ZN(n727) );
  NAND2_X1 U543 ( .A1(n425), .A2(G472), .ZN(n650) );
  NAND2_X1 U544 ( .A1(n411), .A2(n409), .ZN(n597) );
  INV_X1 U545 ( .A(n688), .ZN(n411) );
  XNOR2_X1 U546 ( .A(n484), .B(n482), .ZN(n422) );
  NAND2_X1 U547 ( .A1(n426), .A2(n745), .ZN(n413) );
  XNOR2_X2 U548 ( .A(n414), .B(G146), .ZN(n505) );
  XNOR2_X2 U549 ( .A(n506), .B(KEYINPUT67), .ZN(n753) );
  AND2_X1 U550 ( .A1(n415), .A2(n372), .ZN(n686) );
  XNOR2_X1 U551 ( .A(n684), .B(n416), .ZN(n415) );
  XNOR2_X1 U552 ( .A(n419), .B(n544), .ZN(n738) );
  XNOR2_X1 U553 ( .A(n753), .B(n543), .ZN(n419) );
  NAND2_X1 U554 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U555 ( .A(n423), .B(n654), .ZN(G57) );
  NOR2_X2 U556 ( .A1(n651), .A2(n740), .ZN(n423) );
  XNOR2_X1 U557 ( .A(n424), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U558 ( .A1(n728), .A2(n740), .ZN(n424) );
  NAND2_X1 U559 ( .A1(n425), .A2(G469), .ZN(n729) );
  NAND2_X1 U560 ( .A1(n425), .A2(G475), .ZN(n446) );
  NAND2_X1 U561 ( .A1(n425), .A2(G478), .ZN(n735) );
  NAND2_X1 U562 ( .A1(n425), .A2(G217), .ZN(n464) );
  INV_X1 U563 ( .A(n563), .ZN(n765) );
  NAND2_X1 U564 ( .A1(n434), .A2(n630), .ZN(n433) );
  XNOR2_X1 U565 ( .A(n561), .B(KEYINPUT34), .ZN(n434) );
  XNOR2_X1 U566 ( .A(n443), .B(n442), .ZN(G60) );
  NAND2_X1 U567 ( .A1(n445), .A2(n444), .ZN(n443) );
  XNOR2_X1 U568 ( .A(n446), .B(n374), .ZN(n445) );
  NAND2_X1 U569 ( .A1(n448), .A2(n447), .ZN(n453) );
  NOR2_X1 U570 ( .A1(n639), .A2(KEYINPUT48), .ZN(n447) );
  INV_X1 U571 ( .A(n640), .ZN(n448) );
  NAND2_X1 U572 ( .A1(n640), .A2(KEYINPUT48), .ZN(n452) );
  INV_X1 U573 ( .A(n573), .ZN(n459) );
  NAND2_X1 U574 ( .A1(n459), .A2(n572), .ZN(n458) );
  INV_X1 U575 ( .A(n572), .ZN(n574) );
  INV_X1 U576 ( .A(n683), .ZN(n745) );
  XNOR2_X1 U577 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U578 ( .A(n727), .B(n726), .ZN(n728) );
  INV_X1 U579 ( .A(n688), .ZN(n569) );
  XNOR2_X1 U580 ( .A(n522), .B(n483), .ZN(n484) );
  XOR2_X1 U581 ( .A(n624), .B(KEYINPUT112), .Z(n466) );
  AND2_X1 U582 ( .A1(n530), .A2(G210), .ZN(n467) );
  XNOR2_X1 U583 ( .A(n554), .B(KEYINPUT87), .ZN(n555) );
  XNOR2_X1 U584 ( .A(n597), .B(KEYINPUT68), .ZN(n612) );
  NOR2_X1 U585 ( .A1(n738), .A2(G902), .ZN(n549) );
  INV_X1 U586 ( .A(KEYINPUT63), .ZN(n652) );
  XNOR2_X1 U587 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U588 ( .A(n587), .ZN(n761) );
  XNOR2_X1 U589 ( .A(n469), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U590 ( .A1(G952), .A2(n472), .ZN(n470) );
  XNOR2_X1 U591 ( .A(KEYINPUT92), .B(n470), .ZN(n720) );
  NOR2_X1 U592 ( .A1(n720), .A2(G953), .ZN(n471) );
  XNOR2_X1 U593 ( .A(n471), .B(KEYINPUT93), .ZN(n588) );
  NOR2_X1 U594 ( .A1(G898), .A2(n757), .ZN(n743) );
  NAND2_X1 U595 ( .A1(G902), .A2(n472), .ZN(n585) );
  INV_X1 U596 ( .A(n585), .ZN(n473) );
  NAND2_X1 U597 ( .A1(n743), .A2(n473), .ZN(n474) );
  NAND2_X1 U598 ( .A1(n588), .A2(n474), .ZN(n475) );
  XNOR2_X1 U599 ( .A(KEYINPUT94), .B(n475), .ZN(n487) );
  XOR2_X1 U600 ( .A(G116), .B(G107), .Z(n493) );
  XOR2_X1 U601 ( .A(KEYINPUT16), .B(n493), .Z(n478) );
  XNOR2_X1 U602 ( .A(n531), .B(n507), .ZN(n477) );
  XNOR2_X1 U603 ( .A(n524), .B(n505), .ZN(n480) );
  XNOR2_X1 U604 ( .A(n481), .B(n480), .ZN(n482) );
  AND2_X1 U605 ( .A1(G224), .A2(n761), .ZN(n483) );
  INV_X1 U606 ( .A(n488), .ZN(n646) );
  NAND2_X1 U607 ( .A1(G210), .A2(n486), .ZN(n485) );
  NAND2_X1 U608 ( .A1(G214), .A2(n486), .ZN(n705) );
  XOR2_X1 U609 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n491) );
  NAND2_X1 U610 ( .A1(G234), .A2(n488), .ZN(n489) );
  XNOR2_X1 U611 ( .A(KEYINPUT20), .B(n489), .ZN(n545) );
  NAND2_X1 U612 ( .A1(G221), .A2(n545), .ZN(n490) );
  XNOR2_X1 U613 ( .A(n491), .B(n490), .ZN(n689) );
  XNOR2_X1 U614 ( .A(n492), .B(KEYINPUT9), .ZN(n496) );
  XNOR2_X1 U615 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U616 ( .A(n496), .B(n495), .ZN(n502) );
  XOR2_X1 U617 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n500) );
  NAND2_X1 U618 ( .A1(G234), .A2(n761), .ZN(n497) );
  XNOR2_X1 U619 ( .A(n498), .B(n497), .ZN(n536) );
  NAND2_X1 U620 ( .A1(n536), .A2(G217), .ZN(n499) );
  XNOR2_X1 U621 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U622 ( .A(n502), .B(n501), .ZN(n736) );
  NOR2_X1 U623 ( .A1(G902), .A2(n736), .ZN(n504) );
  XNOR2_X1 U624 ( .A(KEYINPUT100), .B(G478), .ZN(n503) );
  XNOR2_X1 U625 ( .A(n504), .B(n503), .ZN(n573) );
  XNOR2_X1 U626 ( .A(n505), .B(KEYINPUT10), .ZN(n506) );
  XOR2_X1 U627 ( .A(G140), .B(KEYINPUT11), .Z(n510) );
  XNOR2_X1 U628 ( .A(G113), .B(KEYINPUT12), .ZN(n509) );
  XNOR2_X1 U629 ( .A(n510), .B(n509), .ZN(n511) );
  NOR2_X1 U630 ( .A1(G953), .A2(G237), .ZN(n530) );
  XNOR2_X1 U631 ( .A(n512), .B(n753), .ZN(n734) );
  NOR2_X1 U632 ( .A1(G902), .A2(n734), .ZN(n514) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(G475), .ZN(n513) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n708) );
  INV_X1 U635 ( .A(n708), .ZN(n515) );
  AND2_X1 U636 ( .A1(n689), .A2(n515), .ZN(n516) );
  XNOR2_X2 U637 ( .A(n518), .B(n517), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n520), .B(n519), .ZN(n523) );
  NAND2_X1 U639 ( .A1(G227), .A2(n761), .ZN(n525) );
  NOR2_X1 U640 ( .A1(n731), .A2(G902), .ZN(n527) );
  NAND2_X1 U641 ( .A1(n566), .A2(n691), .ZN(n528) );
  XNOR2_X1 U642 ( .A(n528), .B(KEYINPUT103), .ZN(n534) );
  XNOR2_X1 U643 ( .A(KEYINPUT5), .B(G137), .ZN(n529) );
  NOR2_X1 U644 ( .A1(n648), .A2(G902), .ZN(n533) );
  XNOR2_X2 U645 ( .A(n533), .B(G472), .ZN(n611) );
  NAND2_X1 U646 ( .A1(n534), .A2(n611), .ZN(n535) );
  AND2_X1 U647 ( .A1(G221), .A2(n536), .ZN(n544) );
  XNOR2_X1 U648 ( .A(n538), .B(n537), .ZN(n542) );
  XOR2_X1 U649 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n540) );
  XNOR2_X1 U650 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U651 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U652 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n547) );
  NAND2_X1 U653 ( .A1(n545), .A2(G217), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X2 U655 ( .A(n549), .B(n548), .ZN(n688) );
  XOR2_X1 U656 ( .A(KEYINPUT6), .B(n611), .Z(n598) );
  INV_X1 U657 ( .A(n598), .ZN(n557) );
  OR2_X1 U658 ( .A1(n688), .A2(n691), .ZN(n550) );
  NOR2_X1 U659 ( .A1(n557), .A2(n550), .ZN(n551) );
  XNOR2_X1 U660 ( .A(KEYINPUT74), .B(n551), .ZN(n552) );
  NAND2_X1 U661 ( .A1(n552), .A2(n566), .ZN(n553) );
  XNOR2_X1 U662 ( .A(n553), .B(KEYINPUT32), .ZN(n767) );
  INV_X1 U663 ( .A(KEYINPUT44), .ZN(n564) );
  NAND2_X1 U664 ( .A1(n564), .A2(KEYINPUT86), .ZN(n554) );
  XOR2_X1 U665 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n559) );
  NAND2_X1 U666 ( .A1(n689), .A2(n688), .ZN(n692) );
  NOR2_X1 U667 ( .A1(n691), .A2(n692), .ZN(n556) );
  XNOR2_X1 U668 ( .A(n559), .B(n558), .ZN(n714) );
  INV_X1 U669 ( .A(n575), .ZN(n560) );
  NOR2_X1 U670 ( .A1(n572), .A2(n573), .ZN(n630) );
  NAND2_X1 U671 ( .A1(n562), .A2(n563), .ZN(n565) );
  AND2_X1 U672 ( .A1(n566), .A2(n598), .ZN(n567) );
  XNOR2_X1 U673 ( .A(n567), .B(KEYINPUT85), .ZN(n568) );
  NOR2_X1 U674 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U675 ( .A1(n570), .A2(n691), .ZN(n571) );
  XOR2_X1 U676 ( .A(KEYINPUT102), .B(n571), .Z(n770) );
  NAND2_X1 U677 ( .A1(n574), .A2(n573), .ZN(n601) );
  INV_X1 U678 ( .A(n601), .ZN(n668) );
  INV_X1 U679 ( .A(n611), .ZN(n698) );
  NAND2_X1 U680 ( .A1(n594), .A2(n575), .ZN(n576) );
  NOR2_X1 U681 ( .A1(n698), .A2(n576), .ZN(n658) );
  AND2_X1 U682 ( .A1(n698), .A2(n577), .ZN(n701) );
  XNOR2_X1 U683 ( .A(n578), .B(KEYINPUT31), .ZN(n671) );
  NOR2_X1 U684 ( .A1(n658), .A2(n671), .ZN(n579) );
  NOR2_X1 U685 ( .A1(n710), .A2(n579), .ZN(n580) );
  NAND2_X1 U686 ( .A1(n582), .A2(n581), .ZN(n584) );
  XOR2_X1 U687 ( .A(KEYINPUT45), .B(KEYINPUT82), .Z(n583) );
  NOR2_X1 U688 ( .A1(G900), .A2(n585), .ZN(n586) );
  NAND2_X1 U689 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U690 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U691 ( .A(n590), .B(KEYINPUT75), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n698), .A2(n705), .ZN(n592) );
  XNOR2_X1 U693 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U694 ( .A1(n632), .A2(n706), .ZN(n595) );
  NAND2_X1 U695 ( .A1(n670), .A2(n636), .ZN(n677) );
  XOR2_X1 U696 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n605) );
  NOR2_X1 U697 ( .A1(n612), .A2(n598), .ZN(n599) );
  XNOR2_X1 U698 ( .A(n599), .B(KEYINPUT105), .ZN(n600) );
  NOR2_X2 U699 ( .A1(n601), .A2(n600), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n621), .A2(n705), .ZN(n602) );
  XOR2_X1 U701 ( .A(KEYINPUT106), .B(n602), .Z(n603) );
  NAND2_X1 U702 ( .A1(n603), .A2(n691), .ZN(n604) );
  XOR2_X1 U703 ( .A(n605), .B(n604), .Z(n606) );
  NOR2_X1 U704 ( .A1(n629), .A2(n606), .ZN(n679) );
  XOR2_X1 U705 ( .A(KEYINPUT70), .B(n710), .Z(n608) );
  INV_X1 U706 ( .A(KEYINPUT47), .ZN(n607) );
  NAND2_X1 U707 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U708 ( .A1(n609), .A2(KEYINPUT78), .ZN(n618) );
  INV_X1 U709 ( .A(n610), .ZN(n617) );
  NOR2_X1 U710 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U711 ( .A(n613), .B(KEYINPUT28), .ZN(n616) );
  XNOR2_X1 U712 ( .A(n614), .B(KEYINPUT109), .ZN(n615) );
  NAND2_X1 U713 ( .A1(n616), .A2(n615), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n617), .A2(n638), .ZN(n666) );
  NAND2_X1 U715 ( .A1(n618), .A2(n666), .ZN(n620) );
  OR2_X1 U716 ( .A1(KEYINPUT47), .A2(KEYINPUT78), .ZN(n619) );
  XNOR2_X1 U717 ( .A(KEYINPUT111), .B(n621), .ZN(n622) );
  INV_X1 U718 ( .A(KEYINPUT36), .ZN(n624) );
  INV_X1 U719 ( .A(n691), .ZN(n625) );
  NAND2_X1 U720 ( .A1(KEYINPUT70), .A2(n666), .ZN(n626) );
  NAND2_X1 U721 ( .A1(KEYINPUT78), .A2(n626), .ZN(n627) );
  NOR2_X1 U722 ( .A1(n607), .A2(n627), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n710), .A2(KEYINPUT47), .ZN(n628) );
  XOR2_X1 U724 ( .A(KEYINPUT79), .B(n628), .Z(n633) );
  AND2_X1 U725 ( .A1(n629), .A2(n630), .ZN(n631) );
  NAND2_X1 U726 ( .A1(n633), .A2(n768), .ZN(n634) );
  XNOR2_X1 U727 ( .A(n637), .B(KEYINPUT41), .ZN(n704) );
  INV_X1 U728 ( .A(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U729 ( .A1(KEYINPUT2), .A2(n677), .ZN(n642) );
  XNOR2_X1 U730 ( .A(KEYINPUT76), .B(n642), .ZN(n643) );
  NOR2_X1 U731 ( .A1(n683), .A2(n643), .ZN(n645) );
  XNOR2_X1 U732 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  XNOR2_X1 U733 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n653) );
  XOR2_X1 U734 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n656) );
  NAND2_X1 U735 ( .A1(n658), .A2(n668), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U737 ( .A(G104), .B(n657), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n660) );
  NAND2_X1 U739 ( .A1(n658), .A2(n670), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n662) );
  XOR2_X1 U741 ( .A(G107), .B(KEYINPUT27), .Z(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(G9) );
  XNOR2_X1 U743 ( .A(n663), .B(G110), .ZN(G12) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n670), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n665), .B(n664), .ZN(G30) );
  NAND2_X1 U747 ( .A1(n666), .A2(n668), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n667), .B(G146), .ZN(G48) );
  NAND2_X1 U749 ( .A1(n671), .A2(n668), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(G113), .ZN(G15) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(G116), .ZN(G18) );
  INV_X1 U753 ( .A(n673), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n674), .B(KEYINPUT37), .ZN(n675) );
  XNOR2_X1 U755 ( .A(n675), .B(KEYINPUT116), .ZN(n676) );
  XNOR2_X1 U756 ( .A(G125), .B(n676), .ZN(G27) );
  XOR2_X1 U757 ( .A(G134), .B(n677), .Z(n678) );
  XNOR2_X1 U758 ( .A(n678), .B(KEYINPUT117), .ZN(G36) );
  XOR2_X1 U759 ( .A(G140), .B(n679), .Z(G42) );
  NOR2_X1 U760 ( .A1(n760), .A2(KEYINPUT2), .ZN(n680) );
  XNOR2_X1 U761 ( .A(n680), .B(KEYINPUT81), .ZN(n681) );
  NOR2_X1 U762 ( .A1(KEYINPUT2), .A2(n745), .ZN(n684) );
  NOR2_X1 U763 ( .A1(n714), .A2(n704), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U765 ( .A1(n687), .A2(n757), .ZN(n722) );
  NOR2_X1 U766 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U767 ( .A(KEYINPUT49), .B(n690), .ZN(n696) );
  NAND2_X1 U768 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U769 ( .A(n693), .B(KEYINPUT50), .ZN(n694) );
  XNOR2_X1 U770 ( .A(KEYINPUT118), .B(n694), .ZN(n695) );
  NAND2_X1 U771 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U772 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U773 ( .A(KEYINPUT119), .B(n699), .Z(n700) );
  NOR2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U775 ( .A(KEYINPUT51), .B(n702), .Z(n703) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n716) );
  NOR2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  XNOR2_X1 U784 ( .A(KEYINPUT120), .B(n718), .ZN(n719) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(n723), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U787 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n725) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n730) );
  NOR2_X1 U789 ( .A1(n740), .A2(n732), .ZN(G54) );
  INV_X1 U790 ( .A(KEYINPUT59), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U792 ( .A1(n740), .A2(n737), .ZN(G63) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(G66) );
  XOR2_X1 U794 ( .A(n741), .B(G110), .Z(n742) );
  XNOR2_X1 U795 ( .A(KEYINPUT123), .B(n742), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n757), .A2(n745), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n746), .B(KEYINPUT122), .ZN(n750) );
  NAND2_X1 U799 ( .A1(G953), .A2(G224), .ZN(n747) );
  XNOR2_X1 U800 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n748), .A2(G898), .ZN(n749) );
  XOR2_X1 U802 ( .A(n752), .B(n753), .Z(n759) );
  XOR2_X1 U803 ( .A(G227), .B(n759), .Z(n754) );
  NAND2_X1 U804 ( .A1(n754), .A2(G900), .ZN(n755) );
  XOR2_X1 U805 ( .A(KEYINPUT126), .B(n755), .Z(n756) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(KEYINPUT127), .ZN(n764) );
  XNOR2_X1 U808 ( .A(n760), .B(n759), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U811 ( .A(G122), .B(n765), .Z(G24) );
  XOR2_X1 U812 ( .A(G131), .B(n766), .Z(G33) );
  XNOR2_X1 U813 ( .A(G119), .B(n767), .ZN(G21) );
  XNOR2_X1 U814 ( .A(G143), .B(n768), .ZN(G45) );
  XOR2_X1 U815 ( .A(G137), .B(n769), .Z(G39) );
  XOR2_X1 U816 ( .A(G101), .B(n770), .Z(G3) );
endmodule

