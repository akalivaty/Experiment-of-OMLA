//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(G71gat), .ZN(new_n203));
  INV_X1    g002(.A(G78gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n206), .A2(G71gat), .A3(G78gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209));
  OAI22_X1  g008(.A1(new_n209), .A2(new_n206), .B1(new_n203), .B2(new_n204), .ZN(new_n210));
  NOR2_X1   g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT101), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n208), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT102), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT21), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  AOI21_X1  g018(.A(G1gat), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(G8gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n218), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT98), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n221), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(G183gat), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT103), .B(KEYINPUT21), .Z(new_n227));
  OR2_X1    g026(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n226), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n229), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G127gat), .B(G155gat), .ZN(new_n233));
  INV_X1    g032(.A(G211gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G231gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g038(.A(new_n232), .B(new_n239), .Z(new_n240));
  XOR2_X1   g039(.A(G43gat), .B(G50gat), .Z(new_n241));
  INV_X1    g040(.A(KEYINPUT15), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT95), .ZN(new_n244));
  NAND2_X1  g043(.A1(G29gat), .A2(G36gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT94), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n242), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT96), .ZN(new_n249));
  NOR2_X1   g048(.A1(G29gat), .A2(G36gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT95), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(new_n241), .B2(new_n242), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n248), .A2(new_n249), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n251), .B(KEYINPUT93), .ZN(new_n256));
  INV_X1    g055(.A(new_n246), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n243), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n244), .A2(new_n246), .A3(new_n254), .A4(new_n247), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT96), .B1(new_n259), .B2(new_n251), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT97), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(KEYINPUT97), .A3(new_n262), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n255), .A2(KEYINPUT17), .A3(new_n260), .A4(new_n258), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n267), .A2(KEYINPUT99), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(KEYINPUT99), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n265), .B(new_n266), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G85gat), .A2(G92gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT7), .ZN(new_n272));
  INV_X1    g071(.A(G99gat), .ZN(new_n273));
  INV_X1    g072(.A(G106gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT8), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n275), .C1(G85gat), .C2(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G99gat), .B(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G232gat), .A2(G233gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n261), .A2(new_n278), .B1(KEYINPUT41), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G190gat), .B(G218gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n279), .B2(new_n281), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n280), .A2(KEYINPUT41), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT106), .ZN(new_n288));
  XOR2_X1   g087(.A(G134gat), .B(G162gat), .Z(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n285), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n279), .A2(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n294), .B2(new_n284), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n240), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT78), .ZN(new_n299));
  XNOR2_X1  g098(.A(G64gat), .B(G92gat), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n299), .B(new_n300), .Z(new_n301));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n302));
  NOR2_X1   g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT67), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(G169gat), .A3(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n310), .A3(new_n311), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AND4_X1   g118(.A1(KEYINPUT25), .A2(new_n309), .A3(new_n315), .A4(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n304), .A3(new_n307), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT66), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n312), .A2(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n303), .B1(new_n306), .B2(new_n305), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n323), .A4(new_n322), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n320), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT27), .B(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n334), .B2(G190gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  OR3_X1    g135(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n315), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n335), .A2(new_n338), .A3(new_n305), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n302), .B1(new_n332), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT22), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G211gat), .A2(G218gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G197gat), .B(G204gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n355));
  NOR2_X1   g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n350), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n350), .ZN(new_n360));
  INV_X1    g159(.A(new_n350), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n355), .B1(new_n361), .B2(new_n356), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n360), .A2(new_n362), .A3(new_n352), .A4(new_n353), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(G226gat), .B(G233gat), .C1(new_n332), .C2(new_n343), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n346), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n346), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n301), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n364), .ZN(new_n373));
  INV_X1    g172(.A(new_n301), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n346), .A2(new_n365), .A3(new_n366), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT30), .B(new_n301), .C1(new_n367), .C2(new_n368), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n371), .A2(KEYINPUT87), .A3(new_n376), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT68), .ZN(new_n383));
  INV_X1    g182(.A(G134gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(G127gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(G127gat), .ZN(new_n386));
  INV_X1    g185(.A(G127gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G120gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G113gat), .ZN(new_n391));
  INV_X1    g190(.A(G113gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G120gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT1), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT69), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT71), .ZN(new_n401));
  OR2_X1    g200(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n390), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n391), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n403), .ZN(new_n407));
  NOR2_X1   g206(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n408));
  OAI21_X1  g207(.A(G120gat), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(KEYINPUT71), .A3(new_n391), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT1), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n406), .A2(new_n410), .A3(new_n411), .A4(new_n386), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n384), .A2(G127gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n400), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT2), .ZN(new_n418));
  INV_X1    g217(.A(G155gat), .ZN(new_n419));
  INV_X1    g218(.A(G162gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G141gat), .B(G148gat), .Z(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n419), .A3(new_n420), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n430), .B2(new_n417), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT80), .B(new_n416), .C1(new_n428), .C2(new_n429), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n423), .B1(new_n418), .B2(new_n416), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n425), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n415), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n429), .ZN(new_n438));
  NOR3_X1   g237(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n417), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT80), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n430), .A2(new_n426), .A3(new_n417), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n434), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n424), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n443), .B2(new_n424), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n436), .B(new_n437), .C1(new_n448), .C2(new_n415), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n449), .A2(KEYINPUT39), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT3), .B1(new_n446), .B2(new_n447), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n453), .A3(new_n424), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n452), .A2(new_n414), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n443), .A2(new_n424), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT4), .B1(new_n414), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n410), .A2(new_n411), .ZN(new_n458));
  INV_X1    g257(.A(new_n413), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n386), .A3(new_n459), .A4(new_n406), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n435), .A3(new_n461), .A4(new_n400), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n450), .B(new_n451), .C1(new_n465), .C2(new_n437), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n449), .A2(KEYINPUT39), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n414), .B(new_n454), .C1(new_n448), .C2(new_n453), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n437), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n469), .B2(KEYINPUT89), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT82), .B(KEYINPUT0), .Z(new_n471));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G57gat), .B(G85gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT88), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT40), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(new_n437), .A3(new_n463), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n436), .B1(new_n448), .B2(new_n415), .ZN(new_n479));
  INV_X1    g278(.A(new_n437), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT5), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n470), .A3(new_n476), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n382), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT90), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT29), .B1(new_n435), .B2(new_n453), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n364), .ZN(new_n496));
  AND2_X1   g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n359), .A2(new_n302), .A3(new_n363), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n359), .A2(new_n363), .A3(new_n500), .A4(new_n302), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n453), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n497), .B1(new_n502), .B2(new_n456), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n364), .B1(new_n454), .B2(new_n302), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n496), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n447), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n507), .A2(new_n445), .B1(new_n453), .B2(new_n498), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n497), .B1(new_n508), .B2(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(G22gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(KEYINPUT84), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n516), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n511), .A2(KEYINPUT84), .A3(new_n513), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G78gat), .B(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n521), .A3(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n373), .A2(new_n527), .A3(new_n375), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n373), .B2(new_n375), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n526), .B(new_n374), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n528), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n535), .A2(KEYINPUT91), .A3(new_n526), .A4(new_n374), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n374), .B1(new_n373), .B2(new_n375), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n374), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(KEYINPUT38), .ZN(new_n540));
  INV_X1    g339(.A(new_n475), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n483), .A2(new_n541), .A3(new_n485), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n485), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n484), .B1(new_n478), .B2(new_n481), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n475), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n487), .A2(new_n547), .A3(new_n543), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n537), .A2(new_n540), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n382), .A2(new_n488), .A3(new_n550), .A4(new_n491), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n493), .A2(new_n525), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT75), .ZN(new_n554));
  NAND2_X1  g353(.A1(G227gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT64), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n330), .A2(new_n331), .ZN(new_n558));
  INV_X1    g357(.A(new_n320), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n560), .A2(new_n342), .B1(new_n460), .B2(new_n400), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n414), .A2(new_n332), .A3(new_n343), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT32), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(G71gat), .B(G99gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(KEYINPUT33), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n560), .A2(new_n400), .A3(new_n460), .A4(new_n342), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n414), .B1(new_n332), .B2(new_n343), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n556), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT72), .B1(new_n575), .B2(KEYINPUT33), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n572), .A2(new_n576), .A3(new_n567), .A4(new_n564), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT73), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n579));
  INV_X1    g378(.A(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n571), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(KEYINPUT72), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n573), .A2(new_n574), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT33), .B1(new_n583), .B2(new_n557), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n584), .A2(new_n570), .B1(KEYINPUT32), .B2(new_n563), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n579), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n554), .B(new_n569), .C1(new_n578), .C2(new_n586), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n583), .A2(KEYINPUT34), .A3(new_n557), .ZN(new_n588));
  INV_X1    g387(.A(new_n555), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT34), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT73), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n582), .A2(new_n585), .A3(new_n579), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n568), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n554), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n595), .A2(new_n554), .A3(new_n591), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n553), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n595), .B(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n603), .A2(new_n553), .ZN(new_n604));
  INV_X1    g403(.A(new_n525), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n542), .A2(new_n547), .A3(new_n543), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n544), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n378), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n552), .A2(new_n599), .A3(new_n604), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n382), .B1(new_n523), .B2(new_n524), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT35), .B1(new_n544), .B2(new_n548), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n597), .C2(new_n598), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n595), .A2(new_n602), .ZN(new_n615));
  AOI211_X1 g414(.A(new_n568), .B(new_n601), .C1(new_n593), .C2(new_n594), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n517), .A2(new_n521), .A3(new_n519), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n521), .B1(new_n517), .B2(new_n519), .ZN(new_n618));
  OAI22_X1  g417(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT35), .B1(new_n619), .B2(new_n609), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n297), .B1(new_n611), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  INV_X1    g422(.A(new_n224), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n261), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n270), .B2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n623), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n268), .A2(new_n269), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n224), .A3(new_n265), .A4(new_n266), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n631), .A2(KEYINPUT18), .A3(new_n627), .A4(new_n625), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT100), .B1(new_n624), .B2(new_n261), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n625), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n627), .B(KEYINPUT13), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n629), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G169gat), .B(G197gat), .Z(new_n638));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n643), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n629), .A2(new_n632), .A3(new_n636), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n278), .B(new_n208), .C1(new_n210), .C2(new_n213), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n216), .B2(new_n278), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(G230gat), .A3(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n216), .A2(new_n278), .A3(KEYINPUT10), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT107), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(KEYINPUT107), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n649), .B(new_n659), .C1(new_n216), .C2(new_n278), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n661), .A2(KEYINPUT108), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT108), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n651), .B(new_n655), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n655), .B1(new_n667), .B2(new_n651), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n648), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n622), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n607), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n382), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT109), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  OAI22_X1  g479(.A1(new_n677), .A2(new_n679), .B1(new_n680), .B2(G8gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n676), .B2(new_n682), .ZN(G1325gat));
  OR2_X1    g482(.A1(new_n597), .A2(new_n598), .ZN(new_n684));
  AOI21_X1  g483(.A(G15gat), .B1(new_n672), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n604), .A2(new_n599), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n685), .B1(G15gat), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n671), .A2(new_n525), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n692), .B(new_n296), .C1(new_n611), .C2(new_n621), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n614), .A2(new_n620), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n614), .B2(new_n620), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n611), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n296), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n693), .B1(new_n699), .B2(new_n692), .ZN(new_n700));
  INV_X1    g499(.A(new_n240), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n670), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT111), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n697), .B2(new_n698), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n705), .A2(new_n706), .A3(new_n693), .A4(new_n702), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n607), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n296), .B(new_n702), .C1(new_n621), .C2(new_n611), .ZN(new_n710));
  INV_X1    g509(.A(G29gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n673), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(G1328gat));
  OAI21_X1  g513(.A(new_n382), .B1(new_n704), .B2(new_n707), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT112), .B(new_n382), .C1(new_n704), .C2(new_n707), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(G36gat), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(G36gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n710), .A2(new_n720), .A3(new_n382), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n710), .A2(new_n724), .A3(new_n684), .ZN(new_n725));
  INV_X1    g524(.A(new_n700), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(new_n686), .A3(new_n702), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT47), .B(new_n725), .C1(new_n727), .C2(new_n724), .ZN(new_n728));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  INV_X1    g528(.A(new_n686), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n704), .B2(new_n707), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(G43gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n728), .B1(new_n732), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n710), .A2(new_n734), .A3(new_n605), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT114), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n726), .A2(new_n525), .A3(new_n702), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n736), .B(KEYINPUT48), .C1(new_n737), .C2(new_n734), .ZN(new_n738));
  INV_X1    g537(.A(new_n735), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n605), .B1(new_n704), .B2(new_n707), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(G50gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(G1331gat));
  AND2_X1   g542(.A1(new_n697), .A2(new_n648), .ZN(new_n744));
  INV_X1    g543(.A(new_n669), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n297), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n673), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n746), .ZN(new_n750));
  INV_X1    g549(.A(new_n382), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n750), .A2(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n747), .A2(new_n382), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT49), .B(G64gat), .Z(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT115), .ZN(G1333gat));
  NAND3_X1  g555(.A1(new_n747), .A2(new_n203), .A3(new_n684), .ZN(new_n757));
  OAI21_X1  g556(.A(G71gat), .B1(new_n750), .B2(new_n686), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g559(.A1(new_n750), .A2(new_n525), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT116), .B(G78gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n240), .A2(new_n647), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n669), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT117), .Z(new_n766));
  AND2_X1   g565(.A1(new_n700), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(G85gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n697), .A2(new_n698), .A3(new_n764), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n673), .A3(new_n669), .ZN(new_n772));
  INV_X1    g571(.A(G85gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n768), .A2(new_n673), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  NOR3_X1   g573(.A1(new_n745), .A2(G92gat), .A3(new_n751), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT119), .Z(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n700), .A2(new_n382), .A3(new_n766), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n777), .B(new_n779), .C1(new_n781), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n273), .A3(new_n669), .A4(new_n684), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n700), .A2(new_n730), .A3(new_n766), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G99gat), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n787), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1338gat));
  NOR2_X1   g592(.A1(new_n525), .A2(G106gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n669), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n767), .A2(new_n605), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n274), .ZN(new_n798));
  INV_X1    g597(.A(new_n796), .ZN(new_n799));
  INV_X1    g598(.A(new_n795), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n274), .B1(new_n767), .B2(new_n605), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(G1339gat));
  NAND4_X1  g602(.A1(new_n240), .A2(new_n648), .A3(new_n745), .A4(new_n296), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n661), .A2(new_n662), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT54), .B(new_n805), .C1(new_n663), .C2(new_n664), .ZN(new_n806));
  XOR2_X1   g605(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n807));
  NAND3_X1  g606(.A1(new_n661), .A2(new_n662), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n654), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n654), .A4(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n665), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n627), .B1(new_n631), .B2(new_n625), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n634), .A2(new_n635), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n642), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n646), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n296), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n669), .A2(new_n646), .A3(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n648), .B2(new_n813), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n296), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n804), .B1(new_n821), .B2(new_n240), .ZN(new_n822));
  INV_X1    g621(.A(new_n619), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n607), .A2(new_n382), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n647), .C1(new_n408), .C2(new_n407), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n822), .A2(new_n673), .A3(new_n612), .A4(new_n684), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n648), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1340gat));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n390), .A3(new_n669), .ZN(new_n830));
  OAI21_X1  g629(.A(G120gat), .B1(new_n827), .B2(new_n745), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n825), .B2(new_n240), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n827), .A2(new_n387), .A3(new_n701), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(G1342gat));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n384), .A3(new_n698), .ZN(new_n836));
  XOR2_X1   g635(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n837));
  XNOR2_X1  g636(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n827), .B2(new_n296), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1343gat));
  INV_X1    g639(.A(G141gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n686), .A2(new_n824), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n647), .A2(new_n665), .A3(new_n811), .A4(new_n812), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n698), .B1(new_n843), .B2(new_n819), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n818), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n820), .A2(new_n296), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT124), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n240), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n804), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT57), .B(new_n605), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n822), .A2(new_n605), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n842), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n841), .B1(new_n855), .B2(new_n647), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n852), .A2(new_n842), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n841), .A3(new_n647), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT58), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n648), .B(new_n842), .C1(new_n851), .C2(new_n854), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n861), .B(new_n858), .C1(new_n862), .C2(new_n841), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(G1344gat));
  INV_X1    g663(.A(G148gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n865), .A3(new_n669), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT125), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  INV_X1    g667(.A(new_n842), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n605), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n822), .B2(new_n605), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n669), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n605), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n745), .B1(new_n854), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(KEYINPUT126), .A3(new_n869), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n868), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g677(.A(KEYINPUT59), .B(new_n865), .C1(new_n855), .C2(new_n669), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n867), .B1(new_n878), .B2(new_n879), .ZN(G1345gat));
  AOI21_X1  g679(.A(G155gat), .B1(new_n857), .B2(new_n240), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n701), .A2(new_n419), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n855), .B2(new_n882), .ZN(G1346gat));
  AOI21_X1  g682(.A(G162gat), .B1(new_n857), .B2(new_n698), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n296), .A2(new_n420), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n855), .B2(new_n885), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n673), .A2(new_n751), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n822), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n823), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n310), .A3(new_n647), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n525), .A3(new_n684), .ZN(new_n891));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n648), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n889), .B2(new_n669), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n891), .A2(new_n311), .A3(new_n745), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n889), .A2(new_n333), .A3(new_n240), .ZN(new_n897));
  OAI21_X1  g696(.A(G183gat), .B1(new_n891), .B2(new_n701), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n889), .A2(new_n340), .A3(new_n698), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n888), .A2(new_n525), .A3(new_n684), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n340), .B1(new_n902), .B2(new_n698), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n686), .A2(new_n887), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n852), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G197gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n911), .A3(new_n647), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n909), .B1(new_n854), .B2(new_n875), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n647), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(new_n911), .ZN(G1352gat));
  INV_X1    g714(.A(new_n909), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n876), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G204gat), .ZN(new_n918));
  INV_X1    g717(.A(G204gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n822), .A2(new_n919), .A3(new_n605), .A4(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT62), .B1(new_n920), .B2(new_n745), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n920), .A2(KEYINPUT62), .A3(new_n745), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n918), .A2(KEYINPUT127), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n876), .B2(new_n916), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n921), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n234), .A3(new_n240), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n240), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n910), .B2(new_n698), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n698), .A2(G218gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n913), .B2(new_n935), .ZN(G1355gat));
endmodule


