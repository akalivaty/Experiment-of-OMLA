//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(G125), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n467), .B1(new_n473), .B2(new_n465), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT68), .Z(G160));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n472), .B2(G112), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n460), .A2(new_n462), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n481), .B2(new_n472), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n470), .A2(new_n483), .A3(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(G124), .B2(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n472), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n472), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n470), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n472), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n494), .A2(new_n496), .A3(G2104), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G75), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n501), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT5), .B(G543), .Z(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G166));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(new_n503), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  OAI211_X1 g096(.A(G543), .B(new_n520), .C1(new_n510), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n523), .B2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n520), .B(new_n518), .C1(new_n510), .C2(new_n521), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n524), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  NAND2_X1  g109(.A1(new_n523), .A2(G52), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT73), .B(G90), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n507), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n523), .A2(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n507), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n527), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NOR2_X1   g128(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n522), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT74), .B(KEYINPUT9), .Z(new_n557));
  NAND4_X1  g132(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n513), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n508), .A2(G91), .A3(new_n518), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n556), .A2(new_n558), .A3(new_n562), .A4(new_n563), .ZN(G299));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n533), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n524), .A2(new_n532), .A3(KEYINPUT75), .A4(new_n526), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(G286));
  OR2_X1    g143(.A1(new_n512), .A2(new_n516), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI221_X1 g147(.A(new_n570), .B1(new_n527), .B2(new_n571), .C1(new_n572), .C2(new_n522), .ZN(G288));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n522), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n507), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n528), .A2(G86), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G60), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n513), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n523), .A2(G47), .B1(new_n583), .B2(new_n510), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n528), .A2(G85), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n527), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n508), .A2(KEYINPUT10), .A3(G92), .A4(new_n518), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n513), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n590), .A2(new_n591), .B1(G651), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n523), .A2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n599), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n587), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n587), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G286), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n602), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n610), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n613), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT78), .B1(new_n613), .B2(new_n605), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n547), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g192(.A1(new_n481), .A2(G2105), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(G135), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT79), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n485), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2443), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT81), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT17), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n655), .B(new_n656), .C1(new_n654), .C2(new_n650), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  INV_X1    g243(.A(new_n662), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  AOI22_X1  g245(.A1(new_n666), .A2(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n662), .A3(new_n665), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n673), .C1(new_n666), .C2(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT84), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G6), .ZN(new_n683));
  INV_X1    g258(.A(G305), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n682), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(G1971), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n686), .B(new_n683), .C1(new_n684), .C2(new_n682), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(G1971), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n688), .A2(new_n691), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n570), .B1(new_n527), .B2(new_n571), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G49), .B2(new_n523), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(KEYINPUT86), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n699));
  NAND2_X1  g274(.A1(G288), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G16), .B2(G23), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT87), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n708));
  INV_X1    g283(.A(new_n705), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n703), .B(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n710), .B2(new_n694), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G290), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(new_n682), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n682), .B2(G24), .ZN(new_n717));
  INV_X1    g292(.A(G1986), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n707), .A2(new_n711), .A3(KEYINPUT34), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n618), .A2(G131), .ZN(new_n723));
  OR2_X1    g298(.A1(G95), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G119), .B2(new_n485), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n722), .B1(new_n727), .B2(new_n721), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT85), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT35), .B(G1991), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI22_X1  g306(.A1(new_n729), .A2(new_n731), .B1(new_n717), .B2(new_n718), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n731), .B2(new_n729), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n714), .A2(new_n719), .A3(new_n720), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n736), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(G34), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n742), .A2(new_n743), .A3(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G160), .B2(G29), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G2084), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n682), .A2(G19), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n546), .B2(G16), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n747), .B(new_n748), .S(KEYINPUT91), .Z(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G5), .B2(G16), .ZN(new_n753));
  OR3_X1    g328(.A1(new_n752), .A2(G5), .A3(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(G301), .C2(new_n682), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n746), .B(new_n750), .C1(new_n751), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n721), .A2(G26), .ZN(new_n757));
  INV_X1    g332(.A(G140), .ZN(new_n758));
  NOR2_X1   g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(new_n472), .B2(G116), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n476), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G128), .B2(new_n485), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(new_n721), .ZN(new_n763));
  MUX2_X1   g338(.A(new_n757), .B(new_n763), .S(KEYINPUT28), .Z(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT92), .B(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n682), .A2(G4), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n602), .B2(new_n682), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT90), .B(G1348), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n756), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G21), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G168), .B2(G16), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT95), .B(G1966), .Z(new_n774));
  XOR2_X1   g349(.A(new_n773), .B(new_n774), .Z(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NOR2_X1   g351(.A1(new_n755), .A2(new_n751), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n628), .A2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G28), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n779), .B2(KEYINPUT30), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT30), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT97), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n485), .A2(G129), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT26), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n618), .A2(G141), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n785), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G32), .B(new_n790), .S(G29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT27), .B(G1996), .Z(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT25), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n618), .A2(G139), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n797), .B(new_n798), .C1(new_n472), .C2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G33), .B(new_n800), .S(G29), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2072), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n721), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n721), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2078), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n794), .A2(new_n795), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n721), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n721), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT29), .B(G2090), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AND4_X1   g385(.A1(new_n556), .A2(new_n558), .A3(new_n562), .A4(new_n563), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT23), .B1(new_n811), .B2(new_n682), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n682), .A2(G20), .ZN(new_n813));
  MUX2_X1   g388(.A(KEYINPUT23), .B(new_n812), .S(new_n813), .Z(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(G1956), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(G1956), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n806), .A2(new_n810), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n771), .A2(new_n784), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n745), .A2(G2084), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n720), .A2(new_n733), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n821), .A2(new_n737), .A3(new_n719), .A4(new_n714), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n740), .A2(new_n818), .A3(new_n820), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NOR2_X1   g399(.A1(new_n601), .A2(new_n610), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n528), .A2(G93), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n523), .A2(G55), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n828), .C1(new_n507), .C2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(new_n546), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n836), .B(new_n837), .C1(new_n833), .C2(new_n832), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n830), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT37), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(G145));
  INV_X1    g417(.A(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n476), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G130), .B2(new_n485), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n620), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n727), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n790), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n762), .B(G164), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(new_n850), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n851), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G162), .ZN(new_n858));
  XNOR2_X1  g433(.A(G160), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n628), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n860), .C1(new_n851), .C2(new_n855), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n849), .A2(KEYINPUT102), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(new_n855), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n855), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n861), .B(new_n862), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n869));
  NAND2_X1  g444(.A1(G303), .A2(new_n715), .ZN(new_n870));
  NAND2_X1  g445(.A1(G166), .A2(G290), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n698), .A2(new_n873), .A3(new_n700), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n698), .B2(new_n700), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n871), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n874), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n877), .A2(new_n684), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n684), .B1(new_n877), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n869), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n877), .A2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G305), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(new_n684), .A3(new_n880), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT106), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n881), .A2(new_n882), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(KEYINPUT42), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n612), .B(new_n831), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n595), .A2(new_n596), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(G299), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(KEYINPUT103), .A3(G299), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n597), .B2(new_n811), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(KEYINPUT104), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n897), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n893), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n900), .A2(new_n896), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n904), .B2(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n893), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n892), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n910), .A3(new_n892), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n891), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(new_n888), .B2(KEYINPUT42), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n915), .A2(new_n917), .A3(new_n911), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n830), .A2(new_n605), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(G331));
  AND2_X1   g497(.A1(new_n883), .A2(new_n887), .ZN(new_n923));
  AOI21_X1  g498(.A(G301), .B1(new_n566), .B2(new_n567), .ZN(new_n924));
  NOR2_X1   g499(.A1(G171), .A2(new_n533), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n831), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT109), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n831), .B(new_n928), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n924), .A2(new_n925), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n830), .B(new_n546), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(KEYINPUT108), .A3(new_n932), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n926), .A3(KEYINPUT110), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n931), .A2(KEYINPUT110), .A3(new_n932), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n937), .A2(new_n909), .B1(new_n904), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n923), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n943), .B(new_n896), .C1(new_n901), .C2(new_n903), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(new_n939), .A3(new_n938), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n937), .B2(new_n905), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n888), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n937), .A2(new_n909), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n940), .A2(new_n904), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n888), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT43), .B1(new_n942), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n942), .A2(new_n956), .A3(new_n948), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n942), .B2(new_n952), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n959), .ZN(G397));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n790), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n762), .B(G2067), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n727), .A2(new_n731), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n727), .A2(new_n731), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n474), .A2(G40), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n499), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n718), .A3(new_n715), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT48), .ZN(new_n977));
  INV_X1    g552(.A(G2067), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n762), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n964), .B2(new_n966), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n975), .A2(new_n977), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n963), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n974), .B1(new_n982), .B2(new_n790), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n984));
  INV_X1    g559(.A(new_n974), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(G1996), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n974), .A2(KEYINPUT46), .A3(new_n961), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n981), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G305), .B(G1981), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n463), .A2(new_n464), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n472), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(KEYINPUT67), .C1(new_n472), .C2(new_n471), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n999), .B2(new_n467), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n970), .A3(new_n499), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT112), .B(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n994), .A2(new_n995), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n697), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(G1981), .B2(G305), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n1004), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(G1976), .B2(new_n701), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1010), .B(new_n1011), .C1(G1976), .C2(new_n697), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1005), .B(new_n1012), .C1(new_n1011), .C2(new_n1010), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n973), .A2(G40), .A3(new_n474), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1016), .B2(new_n774), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n499), .A2(new_n1020), .A3(new_n970), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1019), .A2(G40), .A3(new_n474), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G2084), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(new_n1014), .A3(new_n774), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1026), .A2(new_n607), .A3(new_n1002), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1016), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1028), .A2(G1971), .B1(G2090), .B2(new_n1022), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(G166), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  NAND3_X1  g610(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1027), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT63), .B1(new_n1013), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1029), .A2(new_n1002), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(new_n1038), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT63), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1027), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1041), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1009), .B(new_n1040), .C1(new_n1049), .C2(new_n1013), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1002), .B1(new_n1026), .B2(new_n533), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n533), .A2(new_n1002), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT121), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1026), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1016), .A2(new_n1014), .A3(new_n774), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1059), .A2(new_n1017), .A3(new_n1023), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n1033), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1057), .B1(new_n1061), .B2(new_n1054), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1053), .B1(new_n1062), .B2(new_n1052), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1016), .A2(new_n1066), .A3(G2078), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1022), .A2(new_n751), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1016), .B2(G2078), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT62), .B(new_n1053), .C1(new_n1062), .C2(new_n1052), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1065), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT115), .B1(G299), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(G299), .A2(KEYINPUT115), .A3(new_n1075), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n811), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(G299), .B2(new_n1075), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1077), .A2(new_n1078), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1022), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1000), .A2(new_n1015), .A3(new_n973), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1082), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1028), .A2(new_n1085), .B1(new_n1083), .B2(new_n1022), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT116), .B1(new_n811), .B2(KEYINPUT57), .ZN(new_n1091));
  NOR3_X1   g666(.A1(G299), .A2(new_n1080), .A3(new_n1075), .ZN(new_n1092));
  AND3_X1   g667(.A1(G299), .A2(KEYINPUT115), .A3(new_n1075), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n1076), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT117), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n969), .A2(new_n971), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1098), .A2(new_n978), .B1(new_n1022), .B2(new_n769), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n601), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n601), .A2(KEYINPUT119), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n598), .A2(new_n1105), .A3(new_n600), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1104), .A2(new_n1099), .A3(KEYINPUT60), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1022), .A2(new_n769), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(KEYINPUT60), .C1(G2067), .C2(new_n1001), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(KEYINPUT119), .A3(new_n601), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1103), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n1097), .A3(KEYINPUT61), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n973), .A2(new_n1015), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n961), .A4(new_n1000), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT118), .B1(new_n1016), .B2(G1996), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1001), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n547), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1123), .B2(new_n547), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1115), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1101), .B1(new_n1113), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT120), .B(new_n1101), .C1(new_n1113), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1069), .A2(new_n1068), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1116), .A2(G2078), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1066), .B1(new_n969), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1000), .A2(KEYINPUT122), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1134), .A2(new_n1136), .A3(KEYINPUT123), .A4(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1133), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G301), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1067), .A2(G301), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT54), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT125), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1145), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1147), .B(new_n1148), .C1(G301), .C2(new_n1142), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1061), .A2(new_n1054), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT51), .B1(new_n1151), .B2(new_n1057), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1142), .A2(G301), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(KEYINPUT124), .A3(new_n1071), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1156), .A3(G301), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1150), .A2(new_n1152), .A3(new_n1158), .A4(new_n1053), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1074), .B1(new_n1132), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1041), .B(new_n1013), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1050), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n968), .ZN(new_n1163));
  XNOR2_X1  g738(.A(G290), .B(new_n718), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n985), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n991), .B1(new_n1162), .B2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g741(.A(G401), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n867), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(new_n1169), .ZN(new_n1170));
  INV_X1    g744(.A(G319), .ZN(new_n1171));
  OR3_X1    g745(.A1(G229), .A2(new_n1171), .A3(G227), .ZN(new_n1172));
  INV_X1    g746(.A(new_n1172), .ZN(new_n1173));
  OAI211_X1 g747(.A(new_n1170), .B(new_n1173), .C1(new_n957), .C2(new_n958), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


