//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n205), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n221), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n205), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n218), .A2(new_n219), .A3(new_n222), .A4(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT76), .ZN(new_n245));
  INV_X1    g0045(.A(G169), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT67), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT67), .A2(G45), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT75), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G232), .A3(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n255), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(new_n255), .B2(new_n261), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(G33), .B2(G41), .ZN(new_n266));
  OR2_X1    g0066(.A1(G223), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G226), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT74), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT74), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(new_n271), .A3(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n270), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n273), .A2(new_n207), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n246), .B1(new_n264), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n254), .ZN(new_n282));
  INV_X1    g0082(.A(new_n251), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT67), .A2(G45), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(new_n285), .B2(new_n250), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n258), .A2(G232), .A3(new_n260), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT75), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n255), .A2(new_n256), .A3(new_n261), .ZN(new_n289));
  AND4_X1   g0089(.A1(G179), .A2(new_n280), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n245), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G58), .ZN(new_n292));
  INV_X1    g0092(.A(G68), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(G20), .B1(new_n294), .B2(new_n201), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G159), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n273), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT3), .B(G33), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(KEYINPUT74), .ZN(new_n303));
  INV_X1    g0103(.A(G20), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n275), .A2(new_n300), .A3(new_n304), .A4(new_n277), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G68), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT16), .B(new_n299), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n300), .B1(new_n302), .B2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n272), .A2(new_n274), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT7), .A3(new_n304), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n293), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n313), .B2(new_n298), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT69), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n205), .B2(new_n273), .ZN(new_n316));
  NAND4_X1  g0116(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n265), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n308), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n316), .A2(new_n265), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n259), .B2(G20), .ZN(new_n324));
  INV_X1    g0124(.A(new_n320), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n322), .A2(new_n324), .B1(new_n325), .B2(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n280), .A2(new_n288), .A3(new_n289), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G169), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n264), .A2(G179), .A3(new_n280), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT76), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n291), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT18), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n291), .A2(new_n327), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT78), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n319), .A2(new_n326), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT77), .A2(G190), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT77), .A2(G190), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n280), .A2(new_n288), .A3(new_n289), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT17), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  AND4_X1   g0146(.A1(KEYINPUT17), .A2(new_n345), .A3(new_n319), .A4(new_n326), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n319), .A3(new_n326), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n338), .A2(KEYINPUT17), .A3(new_n345), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT78), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n336), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G222), .A2(G1698), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(G223), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n302), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n266), .C1(G77), .C2(new_n302), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n258), .A2(new_n260), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n255), .C1(new_n268), .C2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT68), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n246), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n361), .B(KEYINPUT68), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n259), .A2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n322), .A2(G50), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n304), .A2(G33), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  INV_X1    g0171(.A(new_n296), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n323), .A2(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G50), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n304), .B1(new_n201), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n318), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n369), .B(new_n376), .C1(G50), .C2(new_n320), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n364), .A2(new_n367), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n365), .A2(G190), .B1(new_n380), .B2(new_n377), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n377), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT10), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT70), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n365), .B2(new_n339), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n363), .A2(KEYINPUT70), .A3(G200), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n384), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT10), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n379), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G13), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(G1), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n304), .A2(G68), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT12), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n394), .B(new_n395), .C1(KEYINPUT73), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(KEYINPUT73), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n322), .A2(G68), .A3(new_n368), .ZN(new_n400));
  INV_X1    g0200(.A(G77), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n370), .A2(new_n401), .B1(new_n304), .B2(G68), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT72), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n374), .B2(new_n372), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n318), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n399), .B(new_n400), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n411));
  OAI21_X1  g0211(.A(G238), .B1(new_n360), .B2(KEYINPUT71), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G226), .A2(G1698), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n229), .B2(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n302), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n286), .B1(new_n418), .B2(new_n266), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n415), .A2(new_n302), .B1(G33), .B2(G97), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n255), .B1(new_n422), .B2(new_n258), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n411), .A2(new_n412), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT13), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G190), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n410), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n339), .B1(new_n421), .B2(new_n425), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(new_n425), .A3(G179), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n426), .A2(new_n434), .A3(G169), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n410), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G20), .A2(G77), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n439), .B1(new_n323), .B2(new_n372), .C1(new_n370), .C2(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(new_n318), .B1(new_n401), .B2(new_n325), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n322), .A2(G77), .A3(new_n368), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G244), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n255), .B1(new_n445), .B2(new_n360), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n302), .A2(G238), .A3(G1698), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n302), .A2(G232), .A3(new_n356), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n302), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n450), .B2(new_n266), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n444), .B1(G169), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n366), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n444), .B1(G190), .B2(new_n451), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AND4_X1   g0259(.A1(new_n354), .A2(new_n392), .A3(new_n438), .A4(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n248), .A2(G1), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G257), .A3(new_n258), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT5), .B(G41), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(G274), .A3(new_n258), .A4(new_n461), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n445), .A2(G1698), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n303), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n272), .A2(new_n274), .A3(G250), .A4(G1698), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT4), .A2(G244), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n272), .A2(new_n274), .A3(new_n478), .A4(new_n356), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n258), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n246), .B1(new_n472), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(G97), .A2(G107), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n485), .A2(new_n486), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(KEYINPUT6), .B2(new_n209), .ZN(new_n489));
  XNOR2_X1  g0289(.A(G97), .B(G107), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n491), .A2(new_n304), .B1(new_n401), .B2(new_n372), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n449), .B1(new_n310), .B2(new_n312), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n318), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n273), .A2(G1), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n321), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n325), .A2(new_n209), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n465), .A2(new_n470), .A3(new_n467), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n470), .B1(new_n465), .B2(new_n467), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n275), .A2(new_n277), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT4), .B1(new_n503), .B2(new_n474), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n266), .B1(new_n504), .B2(new_n481), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n366), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n484), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  AOI211_X1 g0307(.A(KEYINPUT81), .B(new_n339), .C1(new_n502), .C2(new_n505), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT81), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(new_n469), .A3(new_n471), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(G200), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n499), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n427), .B2(new_n510), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n507), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n440), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n496), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n440), .A2(new_n325), .ZN(new_n518));
  AOI21_X1  g0318(.A(G20), .B1(new_n275), .B2(new_n277), .ZN(new_n519));
  NOR3_X1   g0319(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n520));
  AOI21_X1  g0320(.A(G20), .B1(G33), .B2(G97), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT19), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR3_X1    g0322(.A1(new_n370), .A2(KEYINPUT19), .A3(new_n209), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n519), .A2(G68), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n318), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n517), .B(new_n518), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n503), .A2(new_n304), .A3(G68), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n522), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n318), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(KEYINPUT83), .A3(new_n518), .A4(new_n517), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT82), .A2(G250), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n461), .A2(new_n253), .A3(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(KEYINPUT82), .A2(new_n208), .B1(new_n248), .B2(G1), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n258), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n273), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n445), .A2(G1698), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G238), .B2(G1698), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n503), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G179), .B(new_n538), .C1(new_n544), .C2(new_n258), .ZN(new_n545));
  INV_X1    g0345(.A(new_n538), .ZN(new_n546));
  INV_X1    g0346(.A(new_n540), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n303), .B2(new_n542), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n266), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n545), .B1(new_n549), .B2(new_n246), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n534), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n210), .A2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(G250), .B2(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G294), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n303), .A2(new_n553), .B1(new_n273), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n266), .B1(new_n461), .B2(new_n466), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n555), .A2(new_n266), .B1(G264), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n366), .A3(new_n467), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n553), .B1(new_n277), .B2(new_n275), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n273), .A2(new_n554), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n266), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(G264), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n467), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n246), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n207), .A2(G20), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT22), .B1(new_n302), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT23), .B1(new_n304), .B2(G107), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n449), .A3(G20), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n304), .A2(G33), .A3(G116), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT90), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n567), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(KEYINPUT22), .A2(G87), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n503), .A2(new_n304), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n525), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n496), .A2(G107), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n320), .A2(G107), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n584), .B(KEYINPUT25), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n558), .B(new_n564), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n581), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n578), .B1(new_n574), .B2(new_n576), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n318), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n586), .ZN(new_n591));
  AOI21_X1  g0391(.A(G200), .B1(new_n557), .B2(new_n467), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n427), .A2(new_n561), .A3(new_n467), .A4(new_n562), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n496), .A2(G87), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(new_n518), .C1(new_n524), .C2(new_n525), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n542), .B1(new_n277), .B2(new_n275), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n266), .B1(new_n597), .B2(new_n540), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n339), .B1(new_n598), .B2(new_n538), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n549), .A2(KEYINPUT84), .A3(G190), .ZN(new_n601));
  OAI211_X1 g0401(.A(G190), .B(new_n538), .C1(new_n544), .C2(new_n258), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT84), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n551), .A2(new_n587), .A3(new_n594), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n515), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n556), .A2(G270), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n467), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT85), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n210), .A2(G1698), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n303), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G303), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n272), .B2(new_n274), .ZN(new_n615));
  AND2_X1   g0415(.A1(G264), .A2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n503), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n503), .A2(KEYINPUT85), .A3(new_n611), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n609), .B1(new_n619), .B2(new_n266), .ZN(new_n620));
  NAND2_X1  g0420(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n621));
  NOR2_X1   g0421(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(G20), .B2(new_n539), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n480), .B(new_n304), .C1(G33), .C2(new_n209), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n621), .B1(new_n525), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n621), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n318), .A2(new_n624), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(G116), .B1(new_n321), .B2(new_n495), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n320), .A2(new_n539), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n620), .A2(G179), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(KEYINPUT87), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(KEYINPUT87), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n619), .A2(new_n266), .ZN(new_n638));
  INV_X1    g0438(.A(new_n609), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(G169), .A3(new_n633), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n635), .A2(new_n636), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n626), .A2(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n620), .A2(new_n644), .A3(new_n246), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n637), .B1(new_n645), .B2(KEYINPUT88), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n643), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT21), .B1(new_n641), .B2(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(KEYINPUT88), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(KEYINPUT89), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n642), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n640), .A2(G200), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(new_n644), .C1(new_n343), .C2(new_n640), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n460), .A2(new_n607), .A3(new_n653), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n594), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n598), .A2(new_n538), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G200), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n531), .A2(new_n318), .B1(new_n325), .B2(new_n440), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(new_n595), .A4(new_n602), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n550), .A2(new_n526), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n664), .B(new_n507), .C1(new_n512), .C2(new_n514), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n653), .B2(new_n587), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT92), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n602), .B(KEYINPUT84), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n550), .A2(new_n534), .B1(new_n670), .B2(new_n600), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n484), .A2(new_n499), .A3(new_n506), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n600), .A2(new_n602), .B1(new_n550), .B2(new_n526), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n674), .A3(new_n669), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n550), .A2(new_n676), .A3(new_n526), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n550), .B2(new_n526), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n668), .B1(new_n673), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n551), .A2(new_n672), .A3(new_n605), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT26), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .A3(new_n675), .A4(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n667), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n460), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n348), .A2(new_n353), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n435), .A2(new_n433), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n434), .B1(new_n426), .B2(G169), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n437), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n455), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n430), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n329), .A2(new_n330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n327), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(new_n334), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n389), .A2(new_n391), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n379), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n689), .A2(new_n702), .ZN(G369));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n653), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n394), .A2(new_n304), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G213), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G343), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n633), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n711), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n653), .B(new_n655), .C1(new_n644), .C2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n704), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n587), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n657), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n711), .B1(new_n582), .B2(new_n586), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n711), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n653), .A2(new_n711), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n718), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n717), .A2(new_n713), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n723), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n223), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n520), .A2(new_n539), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n220), .B2(new_n731), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n515), .A2(new_n606), .A3(new_n711), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n653), .A2(new_n737), .A3(new_n655), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n549), .A2(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n640), .A2(KEYINPUT93), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n658), .A2(new_n366), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n620), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n510), .A2(new_n563), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n620), .A2(G179), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n502), .A2(new_n557), .A3(new_n549), .A4(new_n505), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n748), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n366), .B(new_n609), .C1(new_n619), .C2(new_n266), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT30), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n745), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n753), .B2(new_n711), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n704), .B1(new_n738), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n711), .B1(new_n667), .B2(new_n687), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT29), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT26), .B1(new_n663), .B2(new_n507), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n680), .B(new_n760), .C1(new_n683), .C2(KEYINPUT26), .ZN(new_n761));
  OAI211_X1 g0561(.A(KEYINPUT29), .B(new_n713), .C1(new_n666), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n757), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n736), .B1(new_n763), .B2(G1), .ZN(G364));
  NAND3_X1  g0564(.A1(new_n712), .A2(new_n704), .A3(new_n714), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n393), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n259), .B1(new_n766), .B2(G45), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n731), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n716), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n712), .A2(new_n714), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n769), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n302), .A2(new_n223), .ZN(new_n776));
  INV_X1    g0576(.A(G355), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(G116), .B2(new_n223), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n243), .A2(G45), .B1(new_n221), .B2(new_n285), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n503), .A2(new_n729), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n265), .B1(G20), .B2(new_n246), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n775), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n304), .A2(new_n366), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n339), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n343), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n304), .A2(G179), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(new_n427), .A3(G200), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n789), .A2(new_n292), .B1(new_n449), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n786), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n343), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n311), .B(new_n792), .C1(G50), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n793), .A2(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n787), .A2(G190), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n293), .B1(new_n799), .B2(new_n401), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n427), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n304), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n209), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n207), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n800), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n366), .A2(new_n427), .A3(new_n339), .A4(G20), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT32), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n810), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n795), .A2(new_n806), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  INV_X1    g0615(.A(new_n791), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n796), .A2(new_n815), .B1(new_n816), .B2(G283), .ZN(new_n817));
  INV_X1    g0617(.A(G326), .ZN(new_n818));
  INV_X1    g0618(.A(new_n794), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n554), .B2(new_n802), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n302), .B1(new_n788), .B2(G322), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n614), .B2(new_n804), .C1(new_n822), .C2(new_n799), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G329), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n810), .B(KEYINPUT96), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n814), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n785), .B1(new_n828), .B2(new_n782), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n774), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n770), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  INV_X1    g0632(.A(KEYINPUT100), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT99), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n452), .B2(new_n454), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n456), .A2(new_n246), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(KEYINPUT99), .A3(new_n444), .A4(new_n453), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n458), .A2(new_n457), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n444), .A2(new_n711), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n833), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n458), .A2(new_n457), .B1(new_n444), .B2(new_n711), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n843), .A2(KEYINPUT100), .A3(new_n835), .A4(new_n837), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n713), .B(new_n845), .C1(new_n666), .C2(new_n686), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n455), .A2(new_n711), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n842), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n846), .B1(new_n758), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n769), .B1(new_n851), .B2(new_n757), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n757), .B2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n782), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n772), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n775), .B1(G77), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(KEYINPUT97), .B(G283), .Z(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G294), .A2(new_n788), .B1(new_n796), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n816), .A2(G87), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n859), .B(new_n860), .C1(new_n539), .C2(new_n799), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n803), .B(new_n861), .C1(G303), .C2(new_n794), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n311), .B1(new_n804), .B2(new_n449), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT98), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(new_n864), .C1(new_n822), .C2(new_n826), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n802), .A2(new_n292), .B1(new_n791), .B2(new_n293), .ZN(new_n866));
  INV_X1    g0666(.A(new_n804), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n303), .B(new_n866), .C1(G50), .C2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n826), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(G143), .A2(new_n788), .B1(new_n796), .B2(G150), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n871), .B1(new_n872), .B2(new_n819), .C1(new_n811), .C2(new_n799), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT34), .Z(new_n874));
  OAI21_X1  g0674(.A(new_n865), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n856), .B1(new_n875), .B2(new_n782), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n849), .B2(new_n772), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT101), .Z(new_n878));
  NOR2_X1   g0678(.A1(new_n853), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  NOR3_X1   g0680(.A1(new_n265), .A2(new_n304), .A3(new_n539), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT35), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n491), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n882), .B2(new_n491), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT36), .ZN(new_n885));
  OR3_X1    g0685(.A1(new_n220), .A2(new_n401), .A3(new_n294), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n374), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n259), .B(G13), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n299), .B1(new_n305), .B2(new_n307), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n309), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n308), .A2(new_n318), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n326), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n709), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n697), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n349), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT37), .B1(new_n338), .B2(new_n345), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT102), .B1(new_n327), .B2(new_n894), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT102), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n901), .B(new_n709), .C1(new_n319), .C2(new_n326), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n899), .B(new_n332), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(KEYINPUT38), .B(new_n904), .C1(new_n354), .C2(new_n895), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n349), .B(new_n698), .C1(new_n900), .C2(new_n902), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n332), .A2(new_n908), .A3(new_n349), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n901), .B1(new_n338), .B2(new_n709), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n327), .A2(KEYINPUT102), .A3(new_n894), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(KEYINPUT37), .A2(new_n907), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n346), .A2(new_n347), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n699), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n906), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n905), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n437), .B(new_n711), .C1(new_n436), .C2(new_n430), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n428), .A2(new_n429), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n437), .A2(new_n711), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n693), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n848), .B1(new_n738), .B2(new_n756), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n336), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n895), .B1(new_n690), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n904), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n906), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT40), .B1(new_n929), .B2(new_n905), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n848), .B(new_n922), .C1(new_n738), .C2(new_n756), .ZN(new_n931));
  AOI22_X1  g0731(.A1(KEYINPUT40), .A2(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n738), .A2(new_n756), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n460), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n933), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n936), .A2(new_n937), .A3(new_n704), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n436), .A2(new_n437), .A3(new_n713), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n929), .B2(new_n905), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n905), .A2(new_n916), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n838), .A2(new_n713), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n846), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n929), .A2(new_n905), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(new_n923), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n699), .A2(new_n894), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n945), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n460), .B(new_n762), .C1(new_n758), .C2(KEYINPUT29), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n702), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n952), .B(new_n954), .Z(new_n955));
  OAI22_X1  g0755(.A1(new_n938), .A2(new_n955), .B1(new_n259), .B2(new_n766), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n938), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n889), .B1(new_n956), .B2(new_n957), .ZN(G367));
  AND2_X1   g0758(.A1(new_n236), .A2(new_n780), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n783), .B1(new_n223), .B2(new_n440), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n816), .A2(G97), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n797), .B2(new_n554), .C1(new_n614), .C2(new_n789), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n303), .B1(new_n819), .B2(new_n822), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n799), .A2(new_n857), .B1(new_n802), .B2(new_n449), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT46), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n804), .B2(new_n539), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n867), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n967), .B(new_n968), .C1(new_n810), .C2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n802), .A2(new_n293), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G143), .B2(new_n794), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n374), .B2(new_n799), .C1(new_n811), .C2(new_n797), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n867), .A2(G58), .B1(new_n816), .B2(G77), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n311), .B1(new_n788), .B2(G150), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n872), .C2(new_n810), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n965), .A2(new_n970), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n775), .B1(new_n959), .B2(new_n960), .C1(new_n979), .C2(new_n854), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT109), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n596), .A2(new_n711), .ZN(new_n982));
  MUX2_X1   g0782(.A(new_n680), .B(new_n663), .S(new_n982), .Z(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n773), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n515), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n499), .A2(new_n711), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n672), .A2(new_n711), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n723), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT105), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n984), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n994), .B(new_n996), .Z(new_n997));
  INV_X1    g0797(.A(new_n725), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n992), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n988), .A2(new_n717), .A3(new_n989), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n711), .B1(new_n1001), .B2(new_n507), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n999), .B2(KEYINPUT42), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1000), .A2(new_n1003), .B1(KEYINPUT43), .B2(new_n984), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n997), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n722), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n724), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n725), .B1(new_n1007), .B2(KEYINPUT106), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT106), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n998), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n715), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n716), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n763), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT107), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n763), .A3(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n992), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n727), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n992), .B1(new_n725), .B2(new_n726), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n723), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n723), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1022), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n763), .B1(new_n1019), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n730), .B(KEYINPUT41), .Z(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n767), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n987), .B1(new_n1005), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G387));
  OR2_X1    g0836(.A1(new_n1014), .A2(new_n763), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1018), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT107), .B1(new_n1014), .B2(new_n763), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n730), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n767), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1014), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT110), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1014), .A2(KEYINPUT110), .A3(new_n1041), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n722), .A2(new_n773), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n780), .B1(new_n232), .B2(new_n285), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n733), .B2(new_n776), .ZN(new_n1048));
  AOI21_X1  g0848(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n323), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1050), .A2(KEYINPUT50), .A3(new_n374), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT50), .B1(new_n1050), .B2(new_n374), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n733), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1048), .A2(new_n1053), .B1(new_n449), .B2(new_n729), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n775), .B1(new_n1054), .B2(new_n784), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n804), .A2(new_n401), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n961), .A2(new_n503), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(G159), .C2(new_n794), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n802), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n516), .A2(new_n1059), .B1(new_n788), .B2(G50), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G68), .A2(new_n798), .B1(new_n796), .B2(new_n1050), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n810), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(G150), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n503), .B1(G116), .B2(new_n816), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n802), .A2(new_n857), .B1(new_n804), .B2(new_n554), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT111), .B(G322), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G317), .A2(new_n788), .B1(new_n794), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n614), .B2(new_n799), .C1(new_n822), .C2(new_n797), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1065), .B1(new_n818), .B2(new_n810), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1055), .B1(new_n1076), .B2(new_n782), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1044), .A2(new_n1045), .B1(new_n1046), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1040), .A2(new_n1078), .ZN(G393));
  AND3_X1   g0879(.A1(new_n1022), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1027), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1041), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n780), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n783), .B1(new_n209), .B2(new_n223), .C1(new_n1084), .C2(new_n240), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT112), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(KEYINPUT113), .A3(new_n775), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT113), .B1(new_n1086), .B2(new_n775), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n797), .A2(new_n374), .B1(new_n293), .B2(new_n804), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n799), .A2(new_n323), .B1(new_n401), .B2(new_n802), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1062), .A2(G143), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1091), .A2(new_n503), .A3(new_n860), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G150), .A2(new_n794), .B1(new_n788), .B2(G159), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G311), .A2(new_n788), .B1(new_n794), .B2(G317), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1059), .A2(G116), .B1(new_n858), .B2(new_n867), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G294), .A2(new_n798), .B1(new_n796), .B2(G303), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n302), .B1(new_n816), .B2(G107), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1093), .A2(new_n1095), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1088), .B1(new_n782), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1087), .B(new_n1104), .C1(new_n992), .C2(new_n985), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1083), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1038), .A2(new_n1039), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT114), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT114), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1019), .A2(new_n1029), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n731), .B1(new_n1113), .B2(new_n1082), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(KEYINPUT115), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT115), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1116), .B2(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(new_n944), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n948), .A2(KEYINPUT39), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n922), .B1(new_n846), .B2(new_n946), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1119), .B(new_n1120), .C1(new_n1121), .C2(new_n940), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n940), .B1(new_n905), .B2(new_n916), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n713), .B(new_n845), .C1(new_n666), .C2(new_n761), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1124), .A2(new_n946), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n922), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n934), .A2(G330), .A3(new_n849), .A4(new_n923), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1122), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n924), .A2(G330), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n922), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1127), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n947), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT116), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n849), .B1(new_n757), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(KEYINPUT116), .B(new_n704), .C1(new_n738), .C2(new_n756), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n922), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1127), .A2(new_n946), .A3(new_n1124), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n460), .A2(new_n757), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n953), .A2(new_n702), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1129), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1122), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1144), .A2(new_n1150), .A3(new_n1151), .A4(new_n1147), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n730), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1130), .A2(new_n1041), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1119), .A2(new_n1120), .A3(new_n771), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n775), .B1(new_n1050), .B2(new_n855), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G97), .A2(new_n798), .B1(new_n796), .B2(G107), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT118), .Z(new_n1158));
  INV_X1    g0958(.A(G283), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n539), .A2(new_n789), .B1(new_n819), .B2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n802), .A2(new_n401), .B1(new_n791), .B2(new_n293), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1160), .A2(new_n302), .A3(new_n805), .A4(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1158), .B(new_n1162), .C1(new_n554), .C2(new_n826), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT119), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n788), .A2(G132), .B1(new_n816), .B2(G50), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n872), .B2(new_n797), .ZN(new_n1167));
  INV_X1    g0967(.A(G128), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n819), .A2(new_n1168), .B1(new_n799), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n302), .B1(new_n802), .B2(new_n811), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1167), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n804), .A2(new_n371), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT53), .ZN(new_n1174));
  INV_X1    g0974(.A(G125), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n1174), .C1(new_n1175), .C2(new_n826), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1165), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1156), .B1(new_n1178), .B2(new_n782), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1155), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1153), .A2(new_n1154), .A3(new_n1180), .ZN(G378));
  NAND2_X1  g0981(.A1(new_n925), .A2(KEYINPUT40), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n930), .A2(new_n931), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n704), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n952), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n950), .B1(new_n1121), .B2(new_n948), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n945), .B(new_n1186), .C1(new_n932), .C2(new_n704), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n377), .A2(new_n894), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n392), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n392), .A2(new_n1188), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  OR3_X1    g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1193), .A2(KEYINPUT121), .A3(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1185), .A2(new_n1187), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1146), .B1(new_n1130), .B2(new_n1144), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n730), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1195), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1185), .A2(new_n1187), .A3(new_n1195), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1152), .A2(new_n1147), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT123), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1208));
  OAI211_X1 g1008(.A(KEYINPUT122), .B(new_n730), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT123), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1211), .C1(new_n1212), .C2(new_n1199), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1202), .A2(new_n1208), .A3(new_n1209), .A4(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1193), .A2(new_n771), .A3(new_n1194), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n775), .B1(G50), .B2(new_n855), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n273), .B(new_n250), .C1(new_n791), .C2(new_n811), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1175), .A2(new_n819), .B1(new_n789), .B2(new_n1168), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n797), .A2(new_n869), .B1(new_n804), .B2(new_n1169), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n872), .B2(new_n799), .C1(new_n371), .C2(new_n802), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1217), .B(new_n1222), .C1(G124), .C2(new_n1062), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n303), .A2(new_n250), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G50), .B1(new_n273), .B2(new_n250), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1223), .A2(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n449), .A2(new_n789), .B1(new_n799), .B2(new_n440), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G116), .B2(new_n794), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n816), .A2(G58), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n797), .B2(new_n209), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1231), .A2(new_n971), .A3(new_n1056), .A4(new_n1225), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1229), .B(new_n1232), .C1(new_n1159), .C2(new_n826), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT58), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(KEYINPUT120), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n854), .B1(new_n1235), .B2(KEYINPUT120), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1216), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1215), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1212), .B2(new_n767), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1214), .A2(new_n1241), .ZN(G375));
  INV_X1    g1042(.A(new_n1135), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT117), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1139), .A2(new_n1141), .A3(new_n1140), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1243), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1146), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1148), .A3(new_n1032), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n922), .A2(new_n771), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n775), .B1(G68), .B2(new_n855), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n799), .A2(new_n371), .B1(new_n802), .B2(new_n374), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT124), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n869), .A2(new_n819), .B1(new_n789), .B2(new_n872), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n797), .A2(new_n1169), .B1(new_n811), .B2(new_n804), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1253), .A2(new_n1256), .A3(new_n503), .A4(new_n1230), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n826), .A2(new_n1168), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n826), .A2(new_n614), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G283), .A2(new_n788), .B1(new_n798), .B2(G107), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n516), .A2(new_n1059), .B1(new_n794), .B2(G294), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n796), .A2(G116), .B1(new_n867), .B2(G97), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n302), .B1(new_n816), .B2(G77), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1257), .A2(new_n1258), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1251), .B1(new_n1265), .B2(new_n782), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1250), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1247), .B2(new_n767), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1249), .A2(new_n1269), .ZN(G381));
  AND3_X1   g1070(.A1(new_n1040), .A2(new_n1078), .A3(new_n831), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1035), .A2(new_n879), .A3(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1108), .A2(KEYINPUT114), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1110), .B1(new_n1019), .B2(new_n1029), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1114), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT115), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1115), .ZN(new_n1278));
  INV_X1    g1078(.A(G378), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1107), .A3(new_n1279), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G375), .A2(new_n1272), .A3(new_n1280), .A4(G381), .ZN(G407));
  NAND2_X1  g1081(.A1(new_n710), .A2(G213), .ZN(new_n1282));
  OR3_X1    g1082(.A1(G375), .A2(G378), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(G409));
  NAND3_X1  g1084(.A1(new_n1214), .A2(G378), .A3(new_n1241), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1212), .A2(new_n1199), .A3(new_n1031), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1279), .B1(new_n1286), .B2(new_n1240), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(new_n1146), .A3(KEYINPUT60), .A4(new_n1135), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n730), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT60), .B1(new_n1247), .B2(new_n1146), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1248), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1296), .B2(new_n1269), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n879), .B(new_n1268), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1289), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(KEYINPUT60), .B2(new_n1148), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1269), .B1(new_n1301), .B2(new_n1292), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n879), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1296), .A2(G384), .A3(new_n1269), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(KEYINPUT125), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1299), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1288), .A2(new_n1282), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1308), .A2(KEYINPUT127), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1288), .A2(new_n1282), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n710), .A2(G213), .A3(G2897), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1306), .B2(new_n1312), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1288), .A2(new_n1282), .A3(new_n1306), .A4(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1310), .A2(new_n1315), .A3(new_n1317), .A4(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n831), .B1(new_n1040), .B2(new_n1078), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1271), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1278), .B2(new_n1107), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n1106), .B(new_n1321), .C1(new_n1277), .C2(new_n1115), .ZN(new_n1324));
  OAI21_X1  g1124(.A(G387), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G390), .A2(new_n1321), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1278), .A2(new_n1107), .A3(new_n1322), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n1035), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1319), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1307), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1325), .A2(new_n1328), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1307), .A2(new_n1331), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1332), .A2(new_n1334), .A3(new_n1315), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1330), .A2(new_n1336), .ZN(G405));
  INV_X1    g1137(.A(new_n1285), .ZN(new_n1338));
  AOI21_X1  g1138(.A(G378), .B1(new_n1214), .B2(new_n1241), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1306), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1341), .A2(new_n1329), .A3(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1329), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(G402));
endmodule


