//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(G125), .B(G140), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OAI211_X1 g008(.A(G146), .B(new_n189), .C1(new_n190), .C2(new_n191), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G110), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n199), .B(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n202), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  OAI221_X1 g020(.A(new_n196), .B1(new_n197), .B2(new_n203), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n197), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT76), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n204), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(KEYINPUT77), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G125), .B(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n193), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(KEYINPUT78), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n195), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT77), .B1(new_n209), .B2(new_n210), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n207), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT72), .A2(G953), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT72), .A2(G953), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XOR2_X1   g035(.A(new_n221), .B(KEYINPUT22), .Z(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n207), .B(new_n224), .C1(new_n215), .C2(new_n216), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n226), .A2(KEYINPUT25), .A3(new_n227), .A4(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(G234), .B2(new_n227), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n229), .A2(new_n235), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(G472), .A2(G902), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT74), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n193), .A2(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n193), .A3(G143), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n241), .A2(new_n244), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G137), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n257), .B2(G137), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n261), .C1(new_n257), .C2(G137), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n260), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n258), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n257), .A2(G137), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT67), .B1(new_n266), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n255), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n241), .A2(new_n244), .A3(KEYINPUT0), .A4(G128), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  OR2_X1    g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n247), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n259), .A2(new_n263), .A3(new_n265), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n266), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT68), .B(new_n255), .C1(new_n270), .C2(new_n271), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT2), .B(G113), .Z(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n201), .B2(G116), .ZN(new_n290));
  INV_X1    g104(.A(G116), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT70), .A3(G119), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n201), .A2(G116), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n288), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n294), .B2(new_n293), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n287), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n294), .ZN(new_n298));
  INV_X1    g112(.A(new_n288), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n293), .A3(new_n294), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(KEYINPUT71), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n286), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n255), .A2(new_n269), .A3(new_n266), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n284), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n303), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n286), .A2(new_n310), .A3(new_n304), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(G101), .ZN(new_n317));
  AOI21_X1  g131(.A(G237), .B1(new_n218), .B2(new_n219), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G210), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n240), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g136(.A(KEYINPUT74), .B(new_n320), .C1(new_n312), .C2(new_n314), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n286), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n307), .A2(KEYINPUT30), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n325), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n328), .A2(new_n304), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n308), .A3(new_n320), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT31), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n334), .A3(new_n308), .A4(new_n320), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n239), .B1(new_n324), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT32), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n333), .B(new_n335), .C1(new_n322), .C2(new_n323), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT32), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(new_n239), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n307), .B(new_n303), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n343), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n343), .A2(KEYINPUT28), .B1(KEYINPUT75), .B2(new_n314), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT29), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(KEYINPUT29), .B2(new_n315), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n227), .B1(new_n347), .B2(new_n321), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n331), .A2(new_n308), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n349), .A2(KEYINPUT29), .A3(new_n320), .ZN(new_n350));
  OAI21_X1  g164(.A(G472), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n238), .B1(new_n342), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G214), .B1(G237), .B2(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT81), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(G110), .B(G122), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(new_n358), .B2(G107), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G101), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(G101), .ZN(new_n367));
  INV_X1    g181(.A(G101), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n359), .A2(new_n362), .A3(new_n368), .A4(new_n363), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n297), .A2(new_n302), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n293), .A2(KEYINPUT5), .A3(new_n294), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(G113), .C1(KEYINPUT5), .C2(new_n294), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n361), .A2(KEYINPUT79), .A3(G104), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n361), .B2(G104), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n358), .A2(G107), .ZN(new_n377));
  OAI211_X1 g191(.A(G101), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n369), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n301), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n357), .B1(new_n371), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n382), .A2(KEYINPUT6), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n371), .A2(new_n381), .A3(new_n357), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT82), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n371), .A2(new_n386), .A3(new_n381), .A4(new_n357), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n382), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n250), .A2(new_n254), .A3(new_n187), .ZN(new_n391));
  OAI211_X1 g205(.A(KEYINPUT83), .B(new_n391), .C1(new_n280), .C2(new_n187), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(KEYINPUT83), .B2(new_n391), .ZN(new_n393));
  INV_X1    g207(.A(G953), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G224), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT84), .Z(new_n396));
  XNOR2_X1  g210(.A(new_n393), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(KEYINPUT7), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n392), .B(new_n399), .C1(KEYINPUT83), .C2(new_n391), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n187), .B1(new_n276), .B2(new_n279), .ZN(new_n401));
  INV_X1    g215(.A(new_n391), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n391), .A2(KEYINPUT83), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT7), .B(new_n395), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n373), .A2(new_n301), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n379), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n381), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n356), .B(KEYINPUT8), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n400), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n385), .A2(new_n387), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G210), .B1(G237), .B2(G902), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n398), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n398), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n355), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT85), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n398), .A2(new_n414), .ZN(new_n420));
  INV_X1    g234(.A(new_n415), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n398), .A2(new_n414), .A3(new_n415), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n355), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G143), .B1(new_n318), .B2(G214), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  AND2_X1   g243(.A1(KEYINPUT72), .A2(G953), .ZN(new_n430));
  NOR2_X1   g244(.A1(KEYINPUT72), .A2(G953), .ZN(new_n431));
  OAI211_X1 g245(.A(G214), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n243), .ZN(new_n433));
  OAI21_X1  g247(.A(G131), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n243), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n220), .A2(G143), .A3(G214), .A4(new_n429), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n260), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n435), .B(new_n260), .C1(new_n436), .C2(new_n437), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n196), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT17), .B(G131), .C1(new_n428), .C2(new_n433), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(KEYINPUT88), .A3(new_n194), .A4(new_n195), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n434), .A2(KEYINPUT89), .A3(new_n435), .A4(new_n438), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n441), .A2(new_n444), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(G113), .B(G122), .Z(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT87), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n358), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n190), .A2(G146), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n214), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n436), .B(new_n437), .C1(new_n455), .C2(new_n260), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n454), .B(new_n456), .C1(new_n455), .C2(new_n434), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n457), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n190), .B(KEYINPUT19), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n195), .B1(new_n460), .B2(G146), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n434), .B2(new_n438), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n451), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G475), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n227), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT90), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT91), .B1(new_n468), .B2(KEYINPUT20), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n464), .A2(new_n470), .A3(new_n471), .A4(new_n467), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n458), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n452), .B1(new_n448), .B2(new_n457), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n227), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G475), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n475), .A2(KEYINPUT92), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT92), .B1(new_n475), .B2(new_n479), .ZN(new_n481));
  XNOR2_X1  g295(.A(G128), .B(G143), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n257), .B1(new_n482), .B2(KEYINPUT13), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n243), .A2(G128), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(KEYINPUT13), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n257), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT94), .ZN(new_n487));
  XNOR2_X1  g301(.A(G116), .B(G122), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n488), .B(KEYINPUT93), .Z(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n361), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n489), .A2(new_n361), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n485), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n291), .A2(KEYINPUT14), .A3(G122), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(G107), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT95), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n482), .B(new_n257), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n490), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT9), .B(G234), .Z(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n503), .A2(new_n234), .A3(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n493), .A2(new_n500), .A3(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(KEYINPUT96), .A3(new_n507), .ZN(new_n508));
  OR3_X1    g322(.A1(new_n501), .A2(KEYINPUT96), .A3(new_n505), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n227), .ZN(new_n510));
  INV_X1    g324(.A(G478), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n510), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(G234), .A2(G237), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n515), .A2(G952), .A3(new_n394), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n227), .B(new_n220), .C1(G234), .C2(G237), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT21), .B(G898), .Z(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n480), .A2(new_n481), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G221), .B1(new_n503), .B2(G902), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n283), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n276), .A2(new_n370), .A3(new_n279), .A4(new_n366), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT10), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n251), .A2(new_n198), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n529), .A2(new_n253), .B1(new_n249), .B2(new_n251), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n530), .B2(new_n379), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n380), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n526), .A2(new_n527), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n220), .A2(G227), .ZN(new_n534));
  XNOR2_X1  g348(.A(G110), .B(G140), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT80), .B1(new_n255), .B2(new_n380), .ZN(new_n538));
  INV_X1    g352(.A(new_n254), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n249), .A2(new_n251), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n380), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT80), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n250), .A2(new_n379), .A3(new_n254), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n544), .A2(KEYINPUT12), .A3(new_n283), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT12), .B1(new_n544), .B2(new_n283), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n537), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n527), .A2(new_n531), .A3(new_n532), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n283), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n533), .ZN(new_n550));
  INV_X1    g364(.A(new_n536), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(G469), .B(G902), .C1(new_n547), .C2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(G469), .B2(G902), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n533), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n551), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n537), .A2(new_n549), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G469), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n525), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n427), .A2(new_n523), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n352), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G101), .ZN(G3));
  NAND2_X1  g378(.A1(new_n339), .A2(new_n227), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G472), .ZN(new_n566));
  INV_X1    g380(.A(new_n238), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n337), .A4(new_n560), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n508), .A2(new_n509), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n507), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n507), .A2(new_n572), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(KEYINPUT33), .A3(new_n506), .A4(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n571), .A2(new_n575), .A3(G478), .A4(new_n227), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n510), .A2(new_n511), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n475), .A2(new_n479), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n475), .A2(KEYINPUT92), .A3(new_n479), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n354), .B1(new_n422), .B2(new_n423), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n584), .A2(new_n585), .A3(new_n521), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n569), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT34), .B(G104), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  XNOR2_X1  g403(.A(new_n510), .B(new_n512), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n448), .A2(new_n457), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n451), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n593), .B2(new_n458), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n594), .B2(new_n465), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n478), .A2(KEYINPUT98), .A3(G475), .ZN(new_n596));
  INV_X1    g410(.A(new_n473), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n464), .A2(new_n467), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n595), .A2(new_n596), .B1(new_n474), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n521), .B(KEYINPUT99), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AND4_X1   g415(.A1(new_n585), .A2(new_n590), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n569), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NAND2_X1  g419(.A1(new_n315), .A2(new_n321), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT74), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n315), .A2(new_n240), .A3(new_n321), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n333), .A2(new_n335), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n337), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n561), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n217), .B(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(new_n227), .C1(new_n234), .C2(G234), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n236), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT37), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n197), .ZN(G12));
  NAND2_X1  g435(.A1(new_n474), .A2(new_n598), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n517), .B1(new_n519), .B2(G900), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n594), .A2(new_n591), .A3(new_n465), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT98), .B1(new_n478), .B2(G475), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n626), .B2(new_n514), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n599), .A2(new_n590), .A3(new_n628), .A4(new_n623), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n585), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n627), .A2(KEYINPUT101), .A3(new_n629), .A4(new_n585), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n339), .A2(new_n340), .A3(new_n239), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n340), .B1(new_n339), .B2(new_n239), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n351), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n634), .A2(new_n637), .A3(new_n560), .A4(new_n618), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  XOR2_X1   g453(.A(new_n424), .B(KEYINPUT38), .Z(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n354), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n321), .B1(new_n331), .B2(new_n308), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n343), .A2(new_n320), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n227), .B1(new_n644), .B2(KEYINPUT102), .ZN(new_n646));
  OAI21_X1  g460(.A(G472), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n635), .B2(new_n636), .ZN(new_n648));
  INV_X1    g462(.A(new_n618), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n480), .A2(new_n481), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n514), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n641), .A2(new_n648), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT103), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n623), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n560), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G143), .ZN(G45));
  OAI211_X1 g473(.A(new_n578), .B(new_n623), .C1(new_n480), .C2(new_n481), .ZN(new_n660));
  INV_X1    g474(.A(new_n560), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n660), .A2(new_n661), .A3(new_n418), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n637), .A2(new_n618), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  INV_X1    g478(.A(G469), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n547), .A2(new_n552), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(new_n227), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n553), .A3(new_n525), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n637), .A2(new_n567), .A3(new_n586), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  NAND4_X1  g485(.A1(new_n637), .A2(new_n567), .A3(new_n602), .A4(new_n668), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G116), .ZN(G18));
  INV_X1    g487(.A(new_n668), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n418), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n585), .A2(new_n676), .A3(new_n668), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n637), .A2(new_n523), .A3(new_n618), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G119), .ZN(G21));
  OAI21_X1  g494(.A(new_n321), .B1(new_n344), .B2(new_n345), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n333), .A2(new_n681), .A3(new_n335), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n565), .A2(G472), .B1(new_n239), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n585), .B(new_n590), .C1(new_n480), .C2(new_n481), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n674), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n685), .A3(new_n567), .A4(new_n601), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n239), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n618), .B(new_n688), .C1(new_n611), .C2(new_n612), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n584), .A2(new_n623), .A3(new_n675), .A4(new_n677), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n187), .ZN(G27));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n559), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n558), .A2(KEYINPUT105), .A3(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n554), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n524), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n660), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n424), .A2(new_n354), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT107), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n352), .A2(new_n698), .A3(new_n699), .A4(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n637), .A2(new_n567), .A3(new_n698), .A4(new_n699), .ZN(new_n704));
  INV_X1    g518(.A(new_n700), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n260), .ZN(G33));
  AND4_X1   g522(.A1(new_n524), .A2(new_n627), .A3(new_n629), .A4(new_n696), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n352), .A2(new_n699), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G134), .ZN(G36));
  NAND2_X1  g525(.A1(new_n650), .A2(new_n578), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT43), .Z(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n613), .A3(new_n618), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n558), .A2(KEYINPUT45), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n665), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n558), .A2(KEYINPUT45), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n558), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(G469), .A2(G902), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n728));
  INV_X1    g542(.A(new_n553), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n724), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n725), .A2(new_n731), .A3(new_n726), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n524), .A3(new_n654), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n613), .A4(new_n618), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n699), .B(KEYINPUT110), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n716), .A2(new_n734), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n739));
  INV_X1    g553(.A(new_n660), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n524), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT47), .B1(new_n733), .B2(new_n524), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n740), .B(new_n699), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n637), .A2(new_n567), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n739), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n743), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n660), .B1(new_n748), .B2(new_n741), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT111), .A3(new_n699), .A4(new_n745), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  INV_X1    g566(.A(new_n648), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n712), .A2(new_n238), .A3(new_n354), .A4(new_n525), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n667), .A2(new_n553), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT49), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n754), .A3(new_n640), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n699), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n674), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n753), .A2(new_n567), .A3(new_n516), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n582), .A2(new_n583), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n760), .A2(new_n761), .A3(new_n578), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n713), .A2(new_n516), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n683), .A2(new_n567), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n640), .A2(new_n354), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n668), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n762), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n759), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(new_n689), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n763), .A2(new_n764), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n736), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n755), .A2(new_n525), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n748), .A2(new_n741), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n777), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n770), .A2(new_n785), .A3(KEYINPUT51), .A4(new_n772), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n394), .A2(G952), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n776), .B2(new_n678), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n672), .A2(new_n679), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n669), .A2(new_n686), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n600), .B1(new_n419), .B2(new_n426), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n584), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n761), .A2(new_n514), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n792), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n584), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n569), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n352), .A2(new_n562), .B1(new_n614), .B2(new_n618), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n790), .A2(new_n791), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n703), .A2(new_n706), .A3(new_n710), .ZN(new_n803));
  INV_X1    g617(.A(new_n626), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n637), .A2(new_n560), .A3(new_n514), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n683), .A2(new_n698), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n649), .B(new_n758), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n802), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n684), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n696), .A2(new_n524), .A3(new_n623), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n648), .A2(new_n649), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n689), .A2(new_n690), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n638), .A2(new_n811), .A3(new_n812), .A4(new_n663), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n649), .B1(new_n342), .B2(new_n351), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n661), .B1(new_n632), .B2(new_n633), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n691), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT52), .A3(new_n663), .A4(new_n811), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n815), .A2(new_n819), .A3(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n808), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n808), .A2(new_n826), .A3(new_n820), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n760), .A2(new_n650), .A3(new_n579), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n808), .A2(new_n822), .A3(new_n826), .A4(new_n823), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n669), .A2(new_n672), .A3(new_n679), .A4(new_n686), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n584), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT112), .B1(new_n792), .B2(new_n584), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n568), .B1(new_n834), .B2(new_n797), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n703), .A2(new_n706), .A3(new_n710), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n805), .A2(new_n806), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n618), .A3(new_n699), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n836), .A2(new_n837), .A3(new_n801), .A4(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n815), .A2(new_n819), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT53), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT54), .B1(new_n830), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n789), .A2(new_n828), .A3(new_n829), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n352), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n771), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(KEYINPUT48), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n847), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n848), .B2(KEYINPUT48), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n781), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(G952), .A2(G953), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n757), .B1(new_n852), .B2(new_n853), .ZN(G75));
  XNOR2_X1  g668(.A(new_n390), .B(new_n397), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT55), .Z(new_n856));
  NAND4_X1  g670(.A1(new_n830), .A2(G210), .A3(new_n842), .A4(G902), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n856), .B1(new_n859), .B2(KEYINPUT117), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n861));
  INV_X1    g675(.A(new_n856), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n861), .A3(new_n858), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n220), .A2(G952), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n859), .B2(KEYINPUT117), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(G51));
  XOR2_X1   g685(.A(new_n724), .B(KEYINPUT57), .Z(new_n872));
  AND3_X1   g686(.A1(new_n830), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n843), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n666), .B(KEYINPUT119), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n830), .A2(new_n842), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n877), .A2(new_n227), .A3(new_n723), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n865), .B1(new_n876), .B2(new_n878), .ZN(G54));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n227), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(new_n464), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n865), .ZN(G60));
  NAND2_X1  g697(.A1(new_n571), .A2(new_n575), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(G478), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT59), .Z(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n885), .B(new_n888), .C1(new_n873), .C2(new_n843), .ZN(new_n889));
  INV_X1    g703(.A(new_n865), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n844), .B2(new_n828), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(new_n885), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(G63));
  NAND2_X1  g708(.A1(G217), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT60), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n830), .A2(new_n842), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n226), .A2(new_n228), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n830), .A2(new_n616), .A3(new_n842), .A4(new_n896), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(KEYINPUT61), .A3(new_n890), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n865), .B1(new_n897), .B2(new_n898), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT61), .A4(new_n900), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n900), .B(KEYINPUT121), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT61), .B1(new_n907), .B2(new_n903), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n900), .A2(new_n910), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n902), .A4(new_n905), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n909), .A2(new_n917), .ZN(G66));
  AOI21_X1  g732(.A(new_n394), .B1(new_n520), .B2(G224), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n802), .A2(new_n220), .B1(KEYINPUT124), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(KEYINPUT124), .B2(new_n919), .ZN(new_n921));
  INV_X1    g735(.A(new_n390), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(G898), .B2(new_n220), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n921), .B(new_n923), .ZN(G69));
  NAND3_X1  g738(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(new_n460), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n218), .A2(G900), .A3(new_n219), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n734), .A2(new_n352), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n803), .B1(new_n929), .B2(new_n809), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n818), .A2(new_n663), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n737), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n737), .B2(new_n933), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n751), .B(new_n930), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n934), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(KEYINPUT126), .A3(new_n751), .A4(new_n930), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n220), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n927), .B(new_n928), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n796), .A2(new_n584), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n846), .A2(new_n655), .A3(new_n758), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n747), .B2(new_n750), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT62), .B1(new_n658), .B2(new_n933), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n658), .A2(KEYINPUT62), .A3(new_n933), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n948), .B(new_n737), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n220), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n926), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n220), .B1(G227), .B2(G900), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n945), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n945), .B2(new_n953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n951), .B2(new_n802), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n642), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n349), .A2(new_n320), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n962), .A2(new_n642), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT127), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n825), .A2(new_n827), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n890), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n959), .B1(new_n943), .B2(new_n802), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n962), .B2(new_n968), .ZN(G57));
endmodule


