

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n591), .A2(n590), .ZN(n593) );
  OR2_X1 U556 ( .A1(n726), .A2(n719), .ZN(n521) );
  NOR2_X1 U557 ( .A1(n631), .A2(n726), .ZN(n522) );
  INV_X1 U558 ( .A(KEYINPUT93), .ZN(n653) );
  XNOR2_X1 U559 ( .A(n654), .B(n653), .ZN(n655) );
  INV_X1 U560 ( .A(n696), .ZN(n677) );
  INV_X1 U561 ( .A(KEYINPUT97), .ZN(n686) );
  INV_X1 U562 ( .A(KEYINPUT32), .ZN(n705) );
  XNOR2_X1 U563 ( .A(n706), .B(n705), .ZN(n714) );
  NAND2_X1 U564 ( .A1(n947), .A2(n521), .ZN(n720) );
  NAND2_X1 U565 ( .A1(n628), .A2(n627), .ZN(n696) );
  NAND2_X1 U566 ( .A1(G8), .A2(n696), .ZN(n726) );
  NOR2_X1 U567 ( .A1(G651), .A2(n545), .ZN(n789) );
  AND2_X1 U568 ( .A1(n593), .A2(n592), .ZN(G160) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n523), .Z(n872) );
  NAND2_X1 U571 ( .A1(n872), .A2(G138), .ZN(n526) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n876) );
  NAND2_X1 U573 ( .A1(G114), .A2(n876), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT83), .B(n524), .Z(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n531) );
  INV_X1 U576 ( .A(G2105), .ZN(n527) );
  AND2_X2 U577 ( .A1(n527), .A2(G2104), .ZN(n873) );
  NAND2_X1 U578 ( .A1(G102), .A2(n873), .ZN(n529) );
  NOR2_X2 U579 ( .A1(G2104), .A2(n527), .ZN(n877) );
  NAND2_X1 U580 ( .A1(G126), .A2(n877), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G164) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U584 ( .A1(G86), .A2(n783), .ZN(n534) );
  INV_X1 U585 ( .A(G651), .ZN(n535) );
  NOR2_X1 U586 ( .A1(G543), .A2(n535), .ZN(n532) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n532), .Z(n786) );
  NAND2_X1 U588 ( .A1(G61), .A2(n786), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n538) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n545) );
  NOR2_X1 U591 ( .A1(n545), .A2(n535), .ZN(n785) );
  NAND2_X1 U592 ( .A1(n785), .A2(G73), .ZN(n536) );
  XOR2_X1 U593 ( .A(KEYINPUT2), .B(n536), .Z(n537) );
  NOR2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U595 ( .A(n539), .B(KEYINPUT78), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G48), .A2(n789), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(G305) );
  NAND2_X1 U598 ( .A1(G49), .A2(n789), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G74), .A2(G651), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U601 ( .A1(n786), .A2(n544), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n545), .A2(G87), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(G288) );
  NAND2_X1 U604 ( .A1(G78), .A2(n785), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT66), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G91), .A2(n783), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G53), .A2(n789), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G65), .A2(n786), .ZN(n551) );
  XNOR2_X1 U610 ( .A(KEYINPUT67), .B(n551), .ZN(n552) );
  NOR2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G299) );
  NAND2_X1 U613 ( .A1(G52), .A2(n789), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G64), .A2(n786), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G90), .A2(n783), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G77), .A2(n785), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT65), .B(n560), .ZN(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT9), .B(n561), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U622 ( .A1(n783), .A2(G89), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G76), .A2(n785), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G51), .A2(n789), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G63), .A2(n786), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U632 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G88), .A2(n783), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G75), .A2(n785), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G50), .A2(n789), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G62), .A2(n786), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G166) );
  INV_X1 U641 ( .A(G166), .ZN(G303) );
  NAND2_X1 U642 ( .A1(G85), .A2(n783), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G72), .A2(n785), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G60), .A2(n786), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT64), .B(n582), .Z(n583) );
  NOR2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n789), .A2(G47), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(G290) );
  NAND2_X1 U650 ( .A1(G101), .A2(n873), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT23), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G113), .A2(n876), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G125), .A2(n877), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n872), .A2(G137), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G160), .A2(G40), .ZN(n626) );
  NOR2_X1 U657 ( .A1(G164), .A2(G1384), .ZN(n627) );
  NOR2_X1 U658 ( .A1(n626), .A2(n627), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n594), .B(KEYINPUT84), .ZN(n748) );
  XOR2_X1 U660 ( .A(KEYINPUT89), .B(n748), .Z(n613) );
  NAND2_X1 U661 ( .A1(G117), .A2(n876), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G129), .A2(n877), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G105), .A2(n873), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT87), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT38), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT88), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G141), .A2(n872), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n869) );
  NAND2_X1 U671 ( .A1(G1996), .A2(n869), .ZN(n612) );
  NAND2_X1 U672 ( .A1(G107), .A2(n876), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G119), .A2(n877), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U675 ( .A(KEYINPUT86), .B(n606), .Z(n610) );
  NAND2_X1 U676 ( .A1(G131), .A2(n872), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G95), .A2(n873), .ZN(n607) );
  AND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n883) );
  NAND2_X1 U680 ( .A1(G1991), .A2(n883), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n926) );
  NAND2_X1 U682 ( .A1(n613), .A2(n926), .ZN(n739) );
  XNOR2_X1 U683 ( .A(n739), .B(KEYINPUT90), .ZN(n625) );
  XNOR2_X1 U684 ( .A(KEYINPUT37), .B(G2067), .ZN(n746) );
  NAND2_X1 U685 ( .A1(G140), .A2(n872), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G104), .A2(n873), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U688 ( .A(KEYINPUT34), .B(n616), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G116), .A2(n876), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G128), .A2(n877), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U692 ( .A(KEYINPUT35), .B(n619), .ZN(n620) );
  XNOR2_X1 U693 ( .A(KEYINPUT85), .B(n620), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(KEYINPUT36), .B(n623), .ZN(n892) );
  NOR2_X1 U696 ( .A1(n746), .A2(n892), .ZN(n931) );
  NAND2_X1 U697 ( .A1(n748), .A2(n931), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n733) );
  XNOR2_X1 U699 ( .A(KEYINPUT91), .B(n626), .ZN(n628) );
  NOR2_X1 U700 ( .A1(G1981), .A2(G305), .ZN(n629) );
  XOR2_X1 U701 ( .A(n629), .B(KEYINPUT24), .Z(n630) );
  NOR2_X1 U702 ( .A1(n726), .A2(n630), .ZN(n731) );
  NAND2_X1 U703 ( .A1(G1976), .A2(G288), .ZN(n956) );
  INV_X1 U704 ( .A(n956), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G66), .A2(n786), .ZN(n638) );
  NAND2_X1 U706 ( .A1(G92), .A2(n783), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G54), .A2(n789), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n785), .A2(G79), .ZN(n634) );
  XOR2_X1 U710 ( .A(KEYINPUT70), .B(n634), .Z(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U713 ( .A(n639), .B(KEYINPUT15), .Z(n758) );
  INV_X1 U714 ( .A(n758), .ZN(n963) );
  NAND2_X1 U715 ( .A1(G56), .A2(n786), .ZN(n640) );
  XOR2_X1 U716 ( .A(KEYINPUT14), .B(n640), .Z(n647) );
  NAND2_X1 U717 ( .A1(n785), .A2(G68), .ZN(n641) );
  XNOR2_X1 U718 ( .A(KEYINPUT69), .B(n641), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n783), .A2(G81), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT12), .B(n642), .Z(n643) );
  NOR2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(KEYINPUT13), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n789), .A2(G43), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n769) );
  NAND2_X1 U726 ( .A1(G1996), .A2(n677), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n650), .B(KEYINPUT26), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G1341), .A2(n696), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n654) );
  NOR2_X1 U730 ( .A1(n769), .A2(n655), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n963), .A2(n662), .ZN(n661) );
  NAND2_X1 U732 ( .A1(G2067), .A2(n677), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(KEYINPUT94), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G1348), .A2(n696), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U736 ( .A(KEYINPUT95), .B(n659), .Z(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n664) );
  OR2_X1 U738 ( .A1(n963), .A2(n662), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n669) );
  INV_X1 U740 ( .A(G299), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n677), .A2(G2072), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(KEYINPUT27), .ZN(n667) );
  INV_X1 U743 ( .A(G1956), .ZN(n958) );
  NOR2_X1 U744 ( .A1(n958), .A2(n677), .ZN(n666) );
  NOR2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n674) );
  NOR2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U749 ( .A(n672), .B(KEYINPUT28), .Z(n673) );
  NAND2_X1 U750 ( .A1(n674), .A2(n673), .ZN(n676) );
  XOR2_X1 U751 ( .A(KEYINPUT29), .B(KEYINPUT96), .Z(n675) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(n682) );
  XOR2_X1 U753 ( .A(G2078), .B(KEYINPUT25), .Z(n1003) );
  NAND2_X1 U754 ( .A1(n677), .A2(n1003), .ZN(n679) );
  NAND2_X1 U755 ( .A1(G1961), .A2(n696), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U757 ( .A(KEYINPUT92), .B(n680), .Z(n688) );
  NAND2_X1 U758 ( .A1(n688), .A2(G171), .ZN(n681) );
  NAND2_X1 U759 ( .A1(n682), .A2(n681), .ZN(n695) );
  NOR2_X1 U760 ( .A1(G1966), .A2(n726), .ZN(n710) );
  NOR2_X1 U761 ( .A1(G2084), .A2(n696), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n710), .A2(n707), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G8), .A2(n683), .ZN(n684) );
  XNOR2_X1 U764 ( .A(KEYINPUT30), .B(n684), .ZN(n685) );
  NOR2_X1 U765 ( .A1(n685), .A2(G168), .ZN(n687) );
  XNOR2_X1 U766 ( .A(n687), .B(n686), .ZN(n691) );
  NOR2_X1 U767 ( .A1(G171), .A2(n688), .ZN(n689) );
  XNOR2_X1 U768 ( .A(KEYINPUT98), .B(n689), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U770 ( .A(n692), .B(KEYINPUT99), .ZN(n693) );
  XNOR2_X1 U771 ( .A(n693), .B(KEYINPUT31), .ZN(n694) );
  NAND2_X1 U772 ( .A1(n695), .A2(n694), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n708), .A2(G286), .ZN(n704) );
  INV_X1 U774 ( .A(G8), .ZN(n702) );
  NOR2_X1 U775 ( .A1(G2090), .A2(n696), .ZN(n697) );
  XNOR2_X1 U776 ( .A(n697), .B(KEYINPUT100), .ZN(n699) );
  NOR2_X1 U777 ( .A1(n726), .A2(G1971), .ZN(n698) );
  NOR2_X1 U778 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n700), .A2(G303), .ZN(n701) );
  OR2_X1 U780 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U781 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U782 ( .A1(G8), .A2(n707), .ZN(n712) );
  INV_X1 U783 ( .A(n708), .ZN(n709) );
  NOR2_X1 U784 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U785 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n724) );
  NOR2_X1 U787 ( .A1(G1976), .A2(G288), .ZN(n718) );
  NOR2_X1 U788 ( .A1(G1971), .A2(G303), .ZN(n715) );
  NOR2_X1 U789 ( .A1(n718), .A2(n715), .ZN(n953) );
  NAND2_X1 U790 ( .A1(n724), .A2(n953), .ZN(n716) );
  AND2_X1 U791 ( .A1(n522), .A2(n716), .ZN(n717) );
  NOR2_X1 U792 ( .A1(KEYINPUT33), .A2(n717), .ZN(n721) );
  XOR2_X1 U793 ( .A(G1981), .B(G305), .Z(n947) );
  NAND2_X1 U794 ( .A1(n718), .A2(KEYINPUT33), .ZN(n719) );
  OR2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n729) );
  NOR2_X1 U796 ( .A1(G2090), .A2(G303), .ZN(n722) );
  NAND2_X1 U797 ( .A1(G8), .A2(n722), .ZN(n723) );
  NAND2_X1 U798 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U799 ( .A(KEYINPUT101), .B(n725), .Z(n727) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U802 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U804 ( .A(n734), .B(KEYINPUT102), .ZN(n736) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n955) );
  NAND2_X1 U806 ( .A1(n955), .A2(n748), .ZN(n735) );
  NAND2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n751) );
  OR2_X1 U808 ( .A1(n883), .A2(G1991), .ZN(n928) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n737) );
  XOR2_X1 U810 ( .A(n737), .B(KEYINPUT104), .Z(n738) );
  NAND2_X1 U811 ( .A1(n928), .A2(n738), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n742) );
  NOR2_X1 U813 ( .A1(n869), .A2(G1996), .ZN(n741) );
  XNOR2_X1 U814 ( .A(n741), .B(KEYINPUT103), .ZN(n936) );
  NAND2_X1 U815 ( .A1(n742), .A2(n936), .ZN(n743) );
  XNOR2_X1 U816 ( .A(KEYINPUT39), .B(n743), .ZN(n744) );
  NOR2_X1 U817 ( .A1(n931), .A2(n744), .ZN(n745) );
  XNOR2_X1 U818 ( .A(n745), .B(KEYINPUT105), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n746), .A2(n892), .ZN(n923) );
  NAND2_X1 U820 ( .A1(n747), .A2(n923), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U823 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n752) );
  XNOR2_X1 U824 ( .A(n753), .B(n752), .ZN(G329) );
  AND2_X1 U825 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U826 ( .A(G171), .ZN(G301) );
  INV_X1 U827 ( .A(G57), .ZN(G237) );
  INV_X1 U828 ( .A(G132), .ZN(G219) );
  INV_X1 U829 ( .A(G82), .ZN(G220) );
  XOR2_X1 U830 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n757) );
  NAND2_X1 U831 ( .A1(G7), .A2(G661), .ZN(n755) );
  XOR2_X1 U832 ( .A(n755), .B(KEYINPUT10), .Z(n825) );
  NAND2_X1 U833 ( .A1(G567), .A2(n825), .ZN(n756) );
  XNOR2_X1 U834 ( .A(n757), .B(n756), .ZN(G234) );
  INV_X1 U835 ( .A(n769), .ZN(n946) );
  NAND2_X1 U836 ( .A1(n946), .A2(G860), .ZN(G153) );
  NAND2_X1 U837 ( .A1(G868), .A2(G301), .ZN(n760) );
  INV_X1 U838 ( .A(G868), .ZN(n808) );
  NAND2_X1 U839 ( .A1(n758), .A2(n808), .ZN(n759) );
  NAND2_X1 U840 ( .A1(n760), .A2(n759), .ZN(G284) );
  XOR2_X1 U841 ( .A(KEYINPUT71), .B(n808), .Z(n761) );
  NOR2_X1 U842 ( .A1(G286), .A2(n761), .ZN(n762) );
  XNOR2_X1 U843 ( .A(n762), .B(KEYINPUT72), .ZN(n764) );
  NOR2_X1 U844 ( .A1(G299), .A2(G868), .ZN(n763) );
  NOR2_X1 U845 ( .A1(n764), .A2(n763), .ZN(G297) );
  INV_X1 U846 ( .A(G559), .ZN(n765) );
  NOR2_X1 U847 ( .A1(G860), .A2(n765), .ZN(n766) );
  XNOR2_X1 U848 ( .A(KEYINPUT73), .B(n766), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n767), .A2(n963), .ZN(n768) );
  XNOR2_X1 U850 ( .A(n768), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U851 ( .A1(G868), .A2(n769), .ZN(n772) );
  NAND2_X1 U852 ( .A1(G868), .A2(n963), .ZN(n770) );
  NOR2_X1 U853 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U854 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U855 ( .A1(G99), .A2(n873), .ZN(n779) );
  NAND2_X1 U856 ( .A1(G111), .A2(n876), .ZN(n774) );
  NAND2_X1 U857 ( .A1(G135), .A2(n872), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n877), .A2(G123), .ZN(n775) );
  XOR2_X1 U860 ( .A(KEYINPUT18), .B(n775), .Z(n776) );
  NOR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U863 ( .A(n780), .B(KEYINPUT74), .ZN(n927) );
  XNOR2_X1 U864 ( .A(n927), .B(G2096), .ZN(n781) );
  XNOR2_X1 U865 ( .A(n781), .B(KEYINPUT75), .ZN(n782) );
  INV_X1 U866 ( .A(G2100), .ZN(n845) );
  NAND2_X1 U867 ( .A1(n782), .A2(n845), .ZN(G156) );
  NAND2_X1 U868 ( .A1(G93), .A2(n783), .ZN(n784) );
  XNOR2_X1 U869 ( .A(n784), .B(KEYINPUT76), .ZN(n794) );
  NAND2_X1 U870 ( .A1(G80), .A2(n785), .ZN(n788) );
  NAND2_X1 U871 ( .A1(G67), .A2(n786), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G55), .A2(n789), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT77), .B(n790), .ZN(n791) );
  NOR2_X1 U875 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n794), .A2(n793), .ZN(n807) );
  NAND2_X1 U877 ( .A1(n963), .A2(G559), .ZN(n805) );
  XOR2_X1 U878 ( .A(n946), .B(n805), .Z(n795) );
  NOR2_X1 U879 ( .A1(G860), .A2(n795), .ZN(n796) );
  XOR2_X1 U880 ( .A(n807), .B(n796), .Z(G145) );
  XNOR2_X1 U881 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n798) );
  XNOR2_X1 U882 ( .A(G288), .B(KEYINPUT79), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n798), .B(n797), .ZN(n801) );
  XOR2_X1 U884 ( .A(G299), .B(G305), .Z(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(n807), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n801), .B(n800), .ZN(n803) );
  XOR2_X1 U887 ( .A(G290), .B(G303), .Z(n802) );
  XNOR2_X1 U888 ( .A(n803), .B(n802), .ZN(n804) );
  XOR2_X1 U889 ( .A(n804), .B(n946), .Z(n895) );
  XNOR2_X1 U890 ( .A(n805), .B(n895), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n806), .A2(G868), .ZN(n810) );
  NAND2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n810), .A2(n809), .ZN(G295) );
  XOR2_X1 U894 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n814) );
  NAND2_X1 U895 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U897 ( .A1(n812), .A2(G2090), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U899 ( .A1(G2072), .A2(n815), .ZN(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U903 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U904 ( .A1(G96), .A2(n818), .ZN(n829) );
  NAND2_X1 U905 ( .A1(n829), .A2(G2106), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G69), .A2(G120), .ZN(n819) );
  NOR2_X1 U907 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G108), .A2(n820), .ZN(n830) );
  NAND2_X1 U909 ( .A1(n830), .A2(G567), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(n831) );
  NAND2_X1 U911 ( .A1(G661), .A2(G483), .ZN(n823) );
  XNOR2_X1 U912 ( .A(KEYINPUT82), .B(n823), .ZN(n824) );
  NOR2_X1 U913 ( .A1(n831), .A2(n824), .ZN(n828) );
  NAND2_X1 U914 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n825), .ZN(G217) );
  INV_X1 U916 ( .A(n825), .ZN(G223) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n831), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2474), .B(G1981), .Z(n833) );
  XNOR2_X1 U929 ( .A(G1996), .B(G1991), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U931 ( .A(n834), .B(KEYINPUT110), .Z(n836) );
  XNOR2_X1 U932 ( .A(G1971), .B(G1976), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n958), .B(G1961), .ZN(n838) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1966), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U937 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U938 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n848) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2678), .B(KEYINPUT109), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(G227) );
  NAND2_X1 U950 ( .A1(G124), .A2(n877), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n876), .A2(G112), .ZN(n854) );
  NAND2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U954 ( .A1(G136), .A2(n872), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G100), .A2(n873), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U957 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G118), .A2(n876), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G130), .A2(n877), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n873), .A2(G106), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT112), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G142), .A2(n872), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT45), .B(n865), .Z(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n871) );
  XOR2_X1 U967 ( .A(G160), .B(G162), .Z(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n885) );
  NAND2_X1 U970 ( .A1(G139), .A2(n872), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G103), .A2(n873), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U973 ( .A1(G115), .A2(n876), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G127), .A2(n877), .ZN(n878) );
  NAND2_X1 U975 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n919) );
  XOR2_X1 U978 ( .A(n883), .B(n919), .Z(n884) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U980 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U981 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U983 ( .A(n889), .B(n888), .Z(n891) );
  XNOR2_X1 U984 ( .A(G164), .B(n927), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n893) );
  XOR2_X1 U986 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U987 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U988 ( .A(KEYINPUT115), .B(n895), .Z(n897) );
  XOR2_X1 U989 ( .A(G301), .B(G286), .Z(n896) );
  XNOR2_X1 U990 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U991 ( .A(n898), .B(n963), .Z(n899) );
  NOR2_X1 U992 ( .A1(G37), .A2(n899), .ZN(G397) );
  XNOR2_X1 U993 ( .A(G2451), .B(G2427), .ZN(n909) );
  XOR2_X1 U994 ( .A(G2430), .B(G2443), .Z(n901) );
  XNOR2_X1 U995 ( .A(G2435), .B(KEYINPUT107), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U997 ( .A(G2438), .B(G2454), .Z(n903) );
  XNOR2_X1 U998 ( .A(G1341), .B(G1348), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G2446), .B(KEYINPUT108), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(n910), .A2(G14), .ZN(n918) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n918), .ZN(n915) );
  XNOR2_X1 U1006 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1016 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(n922), .B(KEYINPUT50), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n935) );
  XOR2_X1 U1021 ( .A(G160), .B(G2084), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n933) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(KEYINPUT118), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n940) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G162), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(n938), .B(KEYINPUT51), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(n941), .B(KEYINPUT52), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  XOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n1015) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n1015), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(n944), .A2(G29), .ZN(n1024) );
  INV_X1 U1037 ( .A(G16), .ZN(n995) );
  XOR2_X1 U1038 ( .A(n995), .B(KEYINPUT56), .Z(n972) );
  XOR2_X1 U1039 ( .A(G1341), .B(KEYINPUT126), .Z(n945) );
  XOR2_X1 U1040 ( .A(n946), .B(n945), .Z(n970) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G168), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(KEYINPUT123), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT57), .B(n950), .ZN(n968) );
  XOR2_X1 U1045 ( .A(G1961), .B(G301), .Z(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT124), .ZN(n962) );
  NAND2_X1 U1047 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1051 ( .A(n958), .B(G299), .Z(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1054 ( .A(G1348), .B(n963), .Z(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(KEYINPUT125), .B(n966), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1058 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1059 ( .A1(n972), .A2(n971), .ZN(n997) );
  XOR2_X1 U1060 ( .A(G20), .B(G1956), .Z(n976) );
  XNOR2_X1 U1061 ( .A(G1341), .B(G19), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G1981), .B(G6), .ZN(n973) );
  NOR2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n979) );
  XOR2_X1 U1065 ( .A(KEYINPUT59), .B(G1348), .Z(n977) );
  XNOR2_X1 U1066 ( .A(G4), .B(n977), .ZN(n978) );
  NOR2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(KEYINPUT60), .B(n980), .ZN(n984) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G21), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(G5), .B(G1961), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n992) );
  XNOR2_X1 U1073 ( .A(G1986), .B(G24), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G22), .B(G1971), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1976), .B(KEYINPUT127), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n987), .B(G23), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n990), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT61), .B(n993), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1022) );
  XNOR2_X1 U1084 ( .A(KEYINPUT121), .B(G2090), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n998), .B(G35), .ZN(n1014) );
  XNOR2_X1 U1086 ( .A(G2084), .B(G34), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n999), .B(KEYINPUT54), .ZN(n1012) );
  XOR2_X1 U1088 ( .A(G25), .B(G1991), .Z(n1000) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(G28), .ZN(n1009) );
  XNOR2_X1 U1090 ( .A(G2067), .B(G26), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G33), .B(G2072), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1996), .B(G32), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G27), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT53), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(n1016), .B(n1015), .ZN(n1018) );
  INV_X1 U1102 ( .A(G29), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT122), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1025), .ZN(G150) );
  INV_X1 U1109 ( .A(G150), .ZN(G311) );
endmodule

