//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT27), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT64), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n196), .B1(new_n201), .B2(new_n195), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n194), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n196), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n205), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n198), .A2(new_n200), .A3(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n195), .A2(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n203), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n207), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI211_X1 g034(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n217), .C2(G134), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT67), .B1(new_n217), .B2(G134), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n217), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G131), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n219), .B1(new_n229), .B2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n218), .A2(new_n216), .A3(new_n219), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n225), .A4(new_n226), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(G137), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n218), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n222), .A2(new_n227), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n212), .A2(new_n241), .A3(G128), .A4(new_n213), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n244), .B2(new_n202), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n215), .A2(new_n236), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  INV_X1    g062(.A(G119), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G116), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G119), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G119), .ZN(new_n255));
  AND4_X1   g069(.A1(KEYINPUT69), .A2(new_n253), .A3(new_n255), .A4(G116), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT2), .B(G113), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n252), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n253), .A2(new_n255), .A3(G116), .ZN(new_n260));
  INV_X1    g074(.A(new_n250), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n251), .A2(KEYINPUT69), .A3(G116), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n247), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n252), .B2(new_n256), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n263), .A3(new_n257), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n193), .B1(new_n246), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n228), .A2(KEYINPUT71), .A3(new_n235), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT71), .B1(new_n228), .B2(new_n235), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n215), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n238), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n245), .A2(new_n235), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n265), .A2(new_n268), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n228), .A2(new_n235), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n207), .A2(new_n211), .A3(new_n214), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n280), .A3(KEYINPUT72), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n270), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT28), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n283), .B1(new_n282), .B2(KEYINPUT28), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n192), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n273), .A2(KEYINPUT30), .A3(new_n275), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n277), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n192), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n276), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n276), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n286), .B1(new_n300), .B2(new_n285), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n192), .A2(KEYINPUT29), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G472), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n305), .A2(G472), .A3(G902), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT74), .B(new_n294), .C1(new_n287), .C2(new_n288), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n293), .A2(new_n192), .A3(new_n276), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT73), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n286), .A3(new_n284), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT74), .B1(new_n314), .B2(new_n294), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n306), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n294), .B1(new_n287), .B2(new_n288), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n310), .A3(new_n307), .ZN(new_n321));
  NOR2_X1   g135(.A1(G472), .A2(G902), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT32), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n187), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n251), .B2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n249), .A2(new_n243), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n251), .B2(new_n243), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n325), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  OAI22_X1  g144(.A1(new_n329), .A2(G110), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n209), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT77), .B(G125), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n338), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n338), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(G146), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n331), .A2(new_n336), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n329), .A2(G110), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT76), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n337), .A2(KEYINPUT77), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n337), .A2(KEYINPUT77), .ZN(new_n352));
  OAI21_X1  g166(.A(G140), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n353), .B2(new_n339), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n197), .B1(new_n354), .B2(new_n345), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n347), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n328), .A2(new_n330), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n348), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n348), .B(new_n363), .C1(new_n350), .C2(new_n358), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n297), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n365), .A2(KEYINPUT25), .A3(new_n297), .A4(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G234), .B2(new_n297), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n365), .A2(new_n366), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(G902), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n322), .B1(new_n311), .B2(new_n315), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n305), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n316), .A4(new_n304), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n324), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n245), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n340), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n279), .B1(new_n351), .B2(new_n352), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(KEYINPUT91), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n361), .A2(G224), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(KEYINPUT91), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(KEYINPUT7), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n390), .ZN(new_n392));
  OAI211_X1 g206(.A(G224), .B(new_n361), .C1(new_n392), .C2(new_n387), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n392), .B2(new_n387), .ZN(new_n395));
  XOR2_X1   g209(.A(G110), .B(G122), .Z(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT90), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(KEYINPUT8), .Z(new_n398));
  OR2_X1    g212(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(G113), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT5), .B1(new_n252), .B2(new_n256), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n264), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G101), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT82), .A2(G107), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(KEYINPUT82), .A2(G107), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G107), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G104), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n403), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(KEYINPUT3), .ZN(new_n412));
  AOI21_X1  g226(.A(G101), .B1(new_n404), .B2(G107), .ZN(new_n413));
  OR2_X1    g227(.A1(KEYINPUT82), .A2(G107), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n416), .A3(new_n405), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT3), .B1(new_n415), .B2(G104), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n412), .B(new_n413), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT83), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n406), .A2(new_n407), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n404), .B2(KEYINPUT81), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n423), .A3(new_n416), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n412), .A4(new_n413), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n411), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n402), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n402), .A2(new_n427), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n398), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n391), .A2(new_n393), .A3(new_n395), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n420), .A2(new_n426), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n404), .A2(G107), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n412), .B(new_n435), .C1(new_n417), .C2(new_n418), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n436), .B2(G101), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n436), .A2(new_n434), .A3(G101), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(new_n268), .A3(new_n265), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT88), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n439), .B1(new_n433), .B2(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n277), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n445), .A3(new_n428), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n397), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n297), .B1(new_n432), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n428), .B1(new_n441), .B2(KEYINPUT88), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n443), .B1(new_n277), .B2(new_n444), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT89), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n442), .A2(new_n445), .A3(new_n452), .A4(new_n428), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n453), .A3(new_n397), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT6), .B1(new_n446), .B2(new_n397), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n453), .A4(new_n397), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n393), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n448), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n462), .B(KEYINPUT92), .Z(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT93), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n467));
  INV_X1    g281(.A(new_n460), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n456), .B2(new_n457), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n463), .C1(new_n469), .C2(new_n448), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G214), .B1(G237), .B2(G902), .ZN(new_n472));
  AOI21_X1  g286(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT18), .A2(G131), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n341), .A2(new_n197), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n335), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n475), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n482), .B2(new_n473), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n474), .A2(new_n234), .A3(new_n475), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT19), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n332), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n209), .B(new_n487), .C1(new_n341), .C2(new_n486), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n347), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G104), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n481), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT17), .B(G131), .C1(new_n482), .C2(new_n473), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n483), .A2(new_n484), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n355), .A2(new_n347), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n496), .A2(new_n481), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n492), .B1(new_n497), .B2(new_n491), .ZN(new_n498));
  NOR2_X1   g312(.A1(G475), .A2(G902), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT94), .B(new_n492), .C1(new_n497), .C2(new_n491), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n504));
  INV_X1    g318(.A(new_n492), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n491), .B1(new_n496), .B2(new_n481), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n507), .A3(new_n499), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n502), .B1(new_n508), .B2(KEYINPUT20), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n491), .A2(KEYINPUT95), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n497), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n497), .B2(new_n510), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G475), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n361), .A2(G952), .ZN(new_n517));
  NAND2_X1  g331(.A1(G234), .A2(G237), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(G902), .A3(G953), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G116), .ZN(new_n526));
  INV_X1    g340(.A(G116), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G122), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n421), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n407), .B2(new_n406), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n195), .B2(G128), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n243), .A2(KEYINPUT97), .A3(G143), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n243), .A2(G143), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n229), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n538), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G134), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT98), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n542), .A2(new_n537), .B1(new_n534), .B2(new_n535), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n229), .B1(new_n548), .B2(new_n544), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n532), .A2(new_n539), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n536), .A2(new_n538), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G134), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n539), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(KEYINPUT99), .A3(new_n539), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n527), .A3(G122), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n409), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n528), .A2(KEYINPUT14), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n565), .A2(new_n561), .A3(KEYINPUT100), .A4(new_n526), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(new_n564), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n529), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n547), .A2(new_n552), .B1(new_n559), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT9), .B(G234), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n572), .A2(new_n372), .A3(G953), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OAI221_X1 g389(.A(new_n573), .B1(new_n559), .B2(new_n570), .C1(new_n547), .C2(new_n552), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G478), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(G902), .B(new_n579), .C1(new_n575), .C2(new_n576), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n516), .A2(new_n524), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G221), .B1(new_n572), .B2(G902), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n361), .A2(G227), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT80), .ZN(new_n589));
  XNOR2_X1  g403(.A(G110), .B(G140), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n271), .A2(new_n272), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n212), .A2(new_n213), .ZN(new_n595));
  OAI21_X1  g409(.A(G128), .B1(new_n196), .B2(new_n241), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n411), .B1(new_n597), .B2(new_n242), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n433), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n245), .B2(new_n427), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT12), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT85), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n603));
  INV_X1    g417(.A(new_n411), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n433), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n605), .A2(new_n384), .B1(new_n433), .B2(new_n598), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n606), .B2(new_n593), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT85), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n278), .A2(new_n603), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n602), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n384), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n444), .A2(new_n215), .B1(new_n614), .B2(new_n427), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT84), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n599), .B2(new_n613), .ZN(new_n617));
  AOI211_X1 g431(.A(KEYINPUT84), .B(KEYINPUT10), .C1(new_n433), .C2(new_n598), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n615), .B(new_n593), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n592), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n444), .A2(new_n215), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n614), .A2(new_n427), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n594), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(KEYINPUT86), .A3(new_n619), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT86), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n627), .B(new_n594), .C1(new_n621), .C2(new_n624), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n591), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G469), .B1(new_n630), .B2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n591), .A3(new_n628), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n611), .B1(new_n601), .B2(KEYINPUT85), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n607), .A2(new_n608), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n592), .B(new_n619), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n635), .A3(KEYINPUT87), .ZN(new_n636));
  INV_X1    g450(.A(G469), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT87), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n626), .A2(new_n638), .A3(new_n591), .A4(new_n628), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n636), .A2(new_n637), .A3(new_n297), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n587), .B1(new_n631), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n471), .A2(new_n472), .A3(new_n585), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n383), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  INV_X1    g459(.A(new_n462), .ZN(new_n646));
  OAI211_X1 g460(.A(KEYINPUT102), .B(new_n646), .C1(new_n469), .C2(new_n448), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n472), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n646), .B1(new_n469), .B2(new_n448), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n466), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n578), .A2(G902), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n575), .A2(new_n576), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n575), .B2(new_n576), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n577), .B2(G478), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n577), .A2(KEYINPUT103), .A3(G478), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n515), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n652), .A2(new_n524), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n297), .B1(new_n311), .B2(new_n315), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(new_n641), .A3(new_n379), .A4(new_n380), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT34), .B(G104), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  XNOR2_X1  g486(.A(new_n508), .B(KEYINPUT20), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n584), .A2(new_n673), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n652), .A2(new_n514), .A3(new_n524), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n669), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n359), .B(new_n679), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n371), .A2(new_n373), .B1(new_n377), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n667), .A2(new_n380), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n642), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n684), .B(new_n687), .ZN(G12));
  INV_X1    g502(.A(new_n641), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT106), .B(G900), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n522), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n519), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n513), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n674), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n652), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(new_n324), .A3(new_n382), .A4(new_n682), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XOR2_X1   g512(.A(new_n471), .B(KEYINPUT38), .Z(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n316), .ZN(new_n701));
  INV_X1    g515(.A(G472), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n703), .B1(new_n300), .B2(new_n192), .ZN(new_n704));
  OAI211_X1 g518(.A(KEYINPUT107), .B(new_n294), .C1(new_n298), .C2(new_n299), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n308), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n702), .B1(new_n706), .B2(new_n297), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n381), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n515), .A2(new_n583), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n472), .A2(new_n709), .A3(new_n681), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n692), .B(KEYINPUT39), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n641), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT40), .Z(new_n714));
  NAND3_X1  g528(.A1(new_n700), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  NAND2_X1  g530(.A1(new_n663), .A2(new_n692), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n652), .A2(new_n689), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n324), .A3(new_n382), .A4(new_n682), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND3_X1  g534(.A1(new_n636), .A2(new_n297), .A3(new_n639), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT108), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n636), .A2(new_n723), .A3(new_n297), .A4(new_n639), .ZN(new_n724));
  AND4_X1   g538(.A1(KEYINPUT109), .A2(new_n722), .A3(G469), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n640), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n637), .B1(new_n721), .B2(KEYINPUT108), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n724), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n586), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n383), .A2(new_n731), .A3(new_n665), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND3_X1  g548(.A1(new_n383), .A2(new_n731), .A3(new_n675), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AND2_X1   g550(.A1(new_n648), .A2(new_n651), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n586), .C1(new_n729), .C2(new_n725), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n324), .A2(new_n382), .A3(new_n585), .A4(new_n682), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n249), .ZN(G21));
  INV_X1    g556(.A(new_n524), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n648), .A2(new_n651), .A3(new_n743), .A4(new_n710), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n730), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n192), .B1(new_n301), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n746), .B2(new_n301), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n310), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n322), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n666), .A2(KEYINPUT111), .A3(G472), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT111), .B1(new_n666), .B2(G472), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n379), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(G122), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G24));
  INV_X1    g571(.A(new_n717), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n682), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n739), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n465), .A2(new_n472), .A3(new_n466), .A4(new_n470), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n619), .B1(new_n633), .B2(new_n634), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n591), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT113), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n626), .A2(new_n628), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n592), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n770), .A3(new_n591), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(G469), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(G469), .A2(G902), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n640), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n586), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n324), .A3(new_n379), .A4(new_n382), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n763), .B1(new_n777), .B2(new_n717), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n317), .A2(new_n323), .ZN(new_n779));
  INV_X1    g593(.A(new_n379), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n764), .A2(new_n775), .A3(new_n717), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT42), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT114), .B(G131), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G33));
  NAND3_X1  g600(.A1(new_n383), .A2(new_n694), .A3(new_n776), .ZN(new_n787));
  XOR2_X1   g601(.A(KEYINPUT115), .B(G134), .Z(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G36));
  OR2_X1    g603(.A1(new_n630), .A2(KEYINPUT45), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n767), .A2(KEYINPUT45), .A3(new_n769), .A4(new_n771), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(G469), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(new_n773), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT46), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n640), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n586), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n661), .B2(new_n515), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT43), .Z(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n682), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n380), .B2(new_n667), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT44), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n764), .B1(new_n802), .B2(KEYINPUT44), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n798), .A2(new_n803), .A3(new_n712), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  INV_X1    g620(.A(new_n764), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n780), .A3(new_n758), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n324), .B2(new_n382), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n796), .A2(KEYINPUT47), .A3(new_n586), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT47), .B1(new_n796), .B2(new_n586), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n739), .A2(new_n740), .B1(new_n745), .B2(new_n754), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n383), .B(new_n731), .C1(new_n665), .C2(new_n675), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n583), .A2(new_n509), .A3(new_n514), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n817), .A2(new_n818), .B1(new_n516), .B2(new_n661), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n516), .B2(new_n583), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n471), .A2(new_n821), .A3(new_n472), .A4(new_n743), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n668), .A2(new_n822), .B1(new_n642), .B2(new_n683), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n643), .B2(new_n383), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n784), .A2(new_n815), .A3(new_n816), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n673), .A2(new_n513), .A3(new_n583), .A4(new_n692), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n681), .ZN(new_n828));
  INV_X1    g642(.A(new_n640), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n769), .A2(new_n766), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n637), .B1(new_n830), .B2(new_n297), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n586), .B(new_n828), .C1(new_n829), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n764), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n324), .A3(new_n382), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n324), .A3(KEYINPUT118), .A4(new_n382), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n782), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n777), .A2(new_n695), .B1(new_n839), .B2(new_n759), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n826), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n837), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n760), .A2(new_n782), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(KEYINPUT119), .A3(new_n787), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n825), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n751), .A2(new_n752), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n682), .A3(new_n758), .A4(new_n750), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n697), .B1(new_n848), .B2(new_n738), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n648), .A2(new_n651), .A3(new_n710), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n381), .B2(new_n708), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n681), .A2(new_n692), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n774), .A2(new_n586), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n774), .A2(KEYINPUT120), .A3(new_n586), .A4(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n719), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n846), .B1(new_n849), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n324), .A2(new_n382), .A3(new_n682), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n861), .A2(new_n718), .B1(new_n851), .B2(new_n857), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n761), .A2(new_n862), .A3(KEYINPUT52), .A4(new_n697), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n845), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n841), .A2(new_n844), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n784), .A2(new_n815), .A3(new_n816), .A4(new_n824), .ZN(new_n867));
  AND4_X1   g681(.A1(KEYINPUT53), .A2(new_n866), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n814), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n864), .A3(new_n867), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n864), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT54), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NOR2_X1   g690(.A1(KEYINPUT121), .A2(KEYINPUT50), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n472), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n699), .A2(new_n731), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(KEYINPUT121), .B2(KEYINPUT50), .ZN(new_n880));
  INV_X1    g694(.A(new_n725), .ZN(new_n881));
  INV_X1    g695(.A(new_n729), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n586), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n810), .A2(new_n811), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(new_n807), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n754), .A2(new_n520), .A3(new_n800), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(KEYINPUT121), .B(KEYINPUT50), .C1(new_n879), .C2(new_n886), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n730), .A2(new_n519), .A3(new_n764), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n709), .A2(new_n780), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n515), .A3(new_n890), .A4(new_n662), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n760), .A3(new_n800), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n876), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n889), .A2(new_n781), .A3(new_n800), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT48), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n889), .A2(new_n663), .A3(new_n890), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n517), .C1(new_n738), .C2(new_n886), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n887), .A2(new_n876), .A3(new_n893), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n875), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT122), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT49), .B1(new_n881), .B2(new_n882), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n379), .A2(new_n472), .A3(new_n586), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n709), .A2(new_n516), .A3(new_n662), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT49), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n881), .A2(new_n882), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n907), .B(new_n699), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n902), .A2(new_n904), .B1(new_n905), .B2(new_n910), .ZN(G75));
  NOR2_X1   g725(.A1(new_n361), .A2(G952), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n458), .A2(new_n460), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n469), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n872), .A2(new_n873), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(G210), .A3(G902), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n916), .A2(G902), .A3(new_n463), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n915), .A2(new_n918), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n912), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(G51));
  XOR2_X1   g736(.A(new_n773), .B(KEYINPUT57), .Z(new_n923));
  NAND3_X1  g737(.A1(new_n869), .A2(new_n874), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n636), .A2(new_n639), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n297), .B(new_n792), .C1(new_n872), .C2(new_n873), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  INV_X1    g744(.A(new_n912), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n927), .B1(new_n924), .B2(new_n925), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT123), .B1(new_n933), .B2(new_n912), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(G54));
  NAND4_X1  g749(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n503), .A2(new_n507), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n912), .ZN(G60));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT59), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n869), .A2(new_n874), .A3(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n655), .A2(new_n656), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n931), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n945), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT124), .B1(new_n943), .B2(new_n945), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND3_X1  g766(.A1(new_n916), .A2(new_n680), .A3(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n916), .A2(new_n952), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n375), .B(KEYINPUT125), .Z(new_n955));
  OAI211_X1 g769(.A(new_n931), .B(new_n953), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n523), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n815), .A2(new_n824), .A3(new_n816), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n962), .B2(G953), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n456), .B(new_n457), .C1(G898), .C2(new_n361), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G69));
  NAND2_X1  g779(.A1(new_n290), .A2(new_n292), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n487), .B1(new_n341), .B2(new_n486), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT126), .Z(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n713), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n383), .A2(new_n970), .A3(new_n807), .A4(new_n821), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n805), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n761), .A2(new_n697), .A3(new_n719), .ZN(new_n973));
  INV_X1    g787(.A(new_n715), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT62), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n973), .B2(new_n974), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n972), .A2(new_n812), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n969), .B1(new_n977), .B2(new_n361), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n978), .A2(KEYINPUT127), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n805), .A2(new_n787), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n798), .A2(new_n712), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n779), .A2(new_n850), .A3(new_n780), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n973), .B1(new_n778), .B2(new_n783), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n361), .A3(new_n812), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(G900), .A2(G953), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n969), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n979), .A2(new_n980), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n361), .B1(G227), .B2(G900), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n979), .A2(new_n992), .A3(new_n980), .A4(new_n988), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n977), .B2(new_n961), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n293), .A2(new_n276), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n192), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n996), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n984), .A2(new_n812), .A3(new_n985), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n962), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n999), .B(new_n931), .C1(new_n1002), .C2(new_n295), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n295), .A2(new_n996), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n192), .B2(new_n998), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n916), .B2(new_n1005), .ZN(G57));
endmodule


