//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n204), .A2(KEYINPUT71), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n204), .A2(KEYINPUT71), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT69), .B(G113gat), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n208), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT70), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n205), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT26), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT27), .B(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G190gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n230), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT27), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n238));
  AND4_X1   g037(.A1(new_n230), .A2(new_n233), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n237), .B2(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n235), .A3(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT27), .ZN(new_n248));
  INV_X1    g047(.A(G190gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n232), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n229), .B1(new_n240), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n221), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n228), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT24), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n228), .A2(new_n259), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n257), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n228), .A2(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n237), .A2(new_n249), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n257), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n255), .A3(new_n254), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n256), .A2(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n218), .B1(new_n252), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n272), .A2(new_n273), .A3(new_n213), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n215), .B1(new_n274), .B2(new_n210), .ZN(new_n275));
  INV_X1    g074(.A(new_n202), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT71), .B(KEYINPUT1), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(new_n278), .A3(new_n217), .ZN(new_n279));
  INV_X1    g078(.A(new_n205), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n227), .A2(new_n228), .ZN(new_n282));
  AOI21_X1  g081(.A(G190gat), .B1(new_n241), .B2(new_n243), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT28), .B1(new_n283), .B2(new_n248), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n231), .A2(new_n230), .A3(new_n233), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n282), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n256), .A2(new_n264), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n269), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n281), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n271), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G227gat), .A2(G233gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT34), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n295), .B(KEYINPUT64), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT34), .ZN(new_n299));
  OAI22_X1  g098(.A1(new_n296), .A2(new_n297), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G43gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT73), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT74), .ZN(new_n304));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n303), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT33), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n271), .A2(new_n293), .A3(new_n298), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT32), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n313), .B2(KEYINPUT32), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(new_n314), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(KEYINPUT32), .B(new_n313), .C1(new_n311), .C2(new_n312), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n301), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n325), .B(new_n300), .C1(new_n319), .C2(new_n321), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT36), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n313), .A2(KEYINPUT32), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT32), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n320), .B1(new_n331), .B2(new_n314), .ZN(new_n332));
  INV_X1    g131(.A(new_n321), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n300), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT36), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n322), .A2(new_n323), .A3(new_n301), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G211gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT22), .B1(new_n346), .B2(G218gat), .ZN(new_n347));
  XOR2_X1   g146(.A(G197gat), .B(G204gat), .Z(new_n348));
  OAI21_X1  g147(.A(new_n341), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n348), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT76), .B(G211gat), .ZN(new_n351));
  INV_X1    g150(.A(G218gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(KEYINPUT77), .B(new_n350), .C1(new_n353), .C2(KEYINPUT22), .ZN(new_n354));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n347), .A2(new_n348), .ZN(new_n357));
  INV_X1    g156(.A(new_n355), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT78), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n289), .A2(new_n292), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n289), .A2(new_n292), .B1(new_n365), .B2(new_n362), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n360), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n360), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n365), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n252), .B2(new_n270), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n368), .A2(new_n370), .A3(new_n371), .A4(new_n363), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n370), .A3(new_n363), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377));
  XOR2_X1   g176(.A(G64gat), .B(G92gat), .Z(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n340), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n379), .A4(new_n375), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n379), .B(KEYINPUT80), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n279), .A2(KEYINPUT83), .A3(new_n280), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT83), .B1(new_n279), .B2(new_n280), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394));
  INV_X1    g193(.A(G155gat), .ZN(new_n395));
  INV_X1    g194(.A(G162gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n395), .B2(new_n396), .ZN(new_n398));
  INV_X1    g197(.A(G141gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n399), .B2(G148gat), .ZN(new_n401));
  INV_X1    g200(.A(G148gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(G141gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n399), .A2(G148gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n394), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G155gat), .B(G162gat), .Z(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n393), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n409), .A3(new_n393), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(KEYINPUT82), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n409), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n388), .B1(new_n392), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n281), .B2(new_n413), .ZN(new_n420));
  INV_X1    g219(.A(new_n413), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT85), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT85), .B1(new_n420), .B2(new_n422), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n417), .B(new_n418), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n281), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n413), .A3(new_n389), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n429), .A2(KEYINPUT84), .B1(new_n421), .B2(new_n218), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n392), .A2(new_n431), .A3(new_n413), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n387), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n434));
  INV_X1    g233(.A(new_n410), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n436), .A2(new_n428), .A3(new_n389), .A4(new_n414), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n437), .A2(new_n387), .A3(new_n420), .A4(new_n422), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT5), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n426), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G1gat), .B(G29gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT0), .ZN(new_n442));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n447));
  OAI211_X1 g246(.A(new_n426), .B(new_n444), .C1(new_n433), .C2(new_n439), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n447), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n440), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n386), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n356), .A2(new_n359), .A3(new_n365), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n421), .B1(new_n453), .B2(new_n393), .ZN(new_n454));
  OAI211_X1 g253(.A(G228gat), .B(G233gat), .C1(new_n454), .C2(KEYINPUT87), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n411), .A2(new_n365), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n360), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(G22gat), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n459), .A2(new_n454), .A3(G22gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT31), .B(G50gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n459), .A2(new_n454), .A3(G22gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n455), .A3(new_n460), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n463), .B2(new_n468), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n452), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n339), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n430), .A2(new_n387), .A3(new_n432), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n420), .A2(new_n422), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n477), .A2(new_n423), .B1(new_n392), .B2(new_n416), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n474), .B(KEYINPUT39), .C1(new_n478), .C2(new_n387), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n437), .B1(new_n424), .B2(new_n425), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n388), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n444), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n479), .A2(KEYINPUT40), .A3(new_n444), .A4(new_n482), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(new_n446), .A3(new_n386), .A4(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n376), .A2(new_n380), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n375), .A2(new_n489), .A3(new_n372), .A4(new_n367), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n367), .B2(new_n374), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n491), .A2(KEYINPUT38), .A3(new_n383), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n449), .A2(new_n493), .A3(new_n451), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n489), .B1(new_n373), .B2(new_n375), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n380), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT38), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT88), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(KEYINPUT38), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n487), .B(new_n471), .C1(new_n494), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n452), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n335), .A2(new_n471), .A3(new_n337), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n324), .A2(new_n326), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(new_n452), .A3(new_n507), .A4(new_n471), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n473), .A2(new_n502), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  INV_X1    g309(.A(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT14), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G29gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT90), .B1(new_n511), .B2(KEYINPUT14), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT15), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n512), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G43gat), .B(G50gat), .Z(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g320(.A(new_n514), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n517), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT91), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(G1gat), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n530), .A2(new_n531), .A3(G8gat), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n526), .A2(G1gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n529), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n523), .A3(KEYINPUT91), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n525), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n532), .A2(new_n535), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n515), .A2(new_n523), .A3(KEYINPUT91), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n524), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT13), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n540), .B2(new_n524), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n515), .A2(new_n523), .A3(KEYINPUT17), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n536), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n541), .A2(KEYINPUT18), .A3(new_n543), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT12), .Z(new_n558));
  OR2_X1    g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n549), .A2(new_n543), .A3(new_n541), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n545), .B(new_n566), .C1(new_n550), .C2(new_n551), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n567), .A3(new_n562), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n558), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT93), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n571), .A3(new_n558), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n564), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n509), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G57gat), .A2(G64gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G57gat), .A2(G64gat), .ZN(new_n576));
  AND2_X1   g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n539), .B1(KEYINPUT21), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT95), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n395), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(G127gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n596), .A2(new_n597), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n591), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n598), .A3(new_n590), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n525), .A2(new_n537), .ZN(new_n605));
  NAND2_X1  g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT7), .ZN(new_n607));
  XNOR2_X1  g406(.A(G99gat), .B(G106gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n607), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n605), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G190gat), .B(G218gat), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n615), .B(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n547), .A2(new_n620), .A3(new_n548), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n617), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OR3_X1    g426(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n622), .B2(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n604), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n585), .A2(new_n615), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n583), .B(new_n584), .C1(new_n614), .C2(new_n613), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n585), .A2(new_n615), .A3(KEYINPUT10), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G230gat), .ZN(new_n638));
  INV_X1    g437(.A(G233gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n632), .A2(new_n634), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n640), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT97), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  NOR2_X1   g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n642), .A2(new_n647), .A3(new_n651), .A4(new_n645), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n647), .A2(new_n645), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n656), .A2(KEYINPUT98), .A3(new_n651), .A4(new_n642), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n652), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n631), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n574), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n451), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n450), .B1(new_n440), .B2(new_n445), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n448), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(new_n386), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n527), .A2(G8gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n671));
  OAI221_X1 g470(.A(new_n669), .B1(KEYINPUT100), .B2(KEYINPUT42), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  NOR2_X1   g473(.A1(new_n669), .A2(new_n533), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT99), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(G1325gat));
  INV_X1    g476(.A(new_n339), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n661), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n506), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n661), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n661), .A2(new_n471), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  NOR3_X1   g484(.A1(new_n604), .A2(new_n630), .A3(new_n659), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n574), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n516), .A3(new_n665), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n509), .B2(new_n630), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n505), .A2(new_n508), .ZN(new_n693));
  INV_X1    g492(.A(new_n471), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n665), .B2(new_n386), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n502), .A2(new_n695), .A3(new_n327), .A4(new_n338), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n630), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n604), .B(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(new_n573), .A3(new_n659), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n692), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n692), .A2(KEYINPUT102), .A3(new_n699), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n449), .A2(new_n451), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n687), .A2(G36gat), .A3(new_n668), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n707), .B2(new_n668), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  XOR2_X1   g514(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n705), .A2(new_n339), .A3(new_n706), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n564), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n568), .A2(new_n571), .A3(new_n558), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n571), .B1(new_n568), .B2(new_n558), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n680), .A2(G43gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n722), .A3(new_n686), .A4(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n716), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n692), .A2(new_n339), .A3(new_n699), .A4(new_n702), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G43gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT105), .B(new_n729), .C1(new_n727), .C2(G43gat), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT106), .B1(new_n725), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n717), .A2(G43gat), .B1(new_n688), .B2(new_n723), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n735), .B(new_n736), .C1(new_n737), .C2(new_n716), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(G1330gat));
  NOR3_X1   g538(.A1(new_n687), .A2(G50gat), .A3(new_n471), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G50gat), .B1(new_n703), .B2(new_n471), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n705), .A2(new_n694), .A3(new_n706), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n740), .B1(new_n745), .B2(G50gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(G1331gat));
  NOR3_X1   g547(.A1(new_n631), .A2(new_n722), .A3(new_n658), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n697), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n665), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g552(.A(new_n668), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT108), .Z(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n751), .A2(G71gat), .A3(new_n339), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n506), .B(KEYINPUT109), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n750), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(G71gat), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n762), .B(new_n763), .Z(G1334gat));
  NAND2_X1  g563(.A1(new_n751), .A2(new_n694), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  INV_X1    g565(.A(new_n604), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n573), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT111), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n692), .A2(new_n659), .A3(new_n699), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n708), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n697), .A3(new_n698), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT51), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n665), .A2(new_n610), .A3(new_n659), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g575(.A(G92gat), .B1(new_n770), .B2(new_n668), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n659), .A2(new_n611), .A3(new_n386), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT52), .ZN(G1337gat));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n506), .A2(new_n659), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n770), .A2(new_n678), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n773), .A2(new_n782), .B1(new_n783), .B2(new_n781), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n770), .B2(new_n471), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n471), .A2(new_n658), .A3(G106gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT114), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n773), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g589(.A(new_n604), .B(KEYINPUT101), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n635), .A2(new_n640), .A3(new_n636), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n640), .B1(new_n635), .B2(new_n636), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n637), .A2(new_n794), .A3(new_n641), .ZN(new_n796));
  INV_X1    g595(.A(new_n651), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT115), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n657), .A2(new_n655), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(KEYINPUT55), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n635), .A2(new_n640), .A3(new_n636), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n651), .B1(new_n793), .B2(new_n794), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n655), .A2(new_n657), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n813), .A2(KEYINPUT116), .A3(new_n809), .A4(new_n800), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n722), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n549), .A2(new_n541), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n816), .A2(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n557), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n658), .A2(new_n564), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n698), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n812), .A2(new_n814), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n564), .A2(new_n818), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n698), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n791), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n660), .A2(new_n573), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n708), .B(new_n504), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n668), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n573), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(G113gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n212), .B2(new_n830), .ZN(G1340gat));
  NOR2_X1   g631(.A1(new_n829), .A2(new_n658), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(new_n213), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n829), .B2(new_n791), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n604), .A2(new_n595), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n829), .B2(new_n836), .ZN(G1342gat));
  NOR2_X1   g636(.A1(new_n630), .A2(new_n386), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n838), .B(KEYINPUT117), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n828), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(KEYINPUT56), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(KEYINPUT56), .B2(new_n843), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n678), .A2(new_n694), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n665), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n826), .A2(new_n827), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n668), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n399), .B1(new_n852), .B2(new_n573), .ZN(new_n853));
  INV_X1    g652(.A(new_n827), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n804), .B2(new_n805), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n801), .A2(new_n802), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n819), .B1(new_n722), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n630), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT119), .B(new_n819), .C1(new_n722), .C2(new_n860), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n863), .A2(new_n864), .B1(new_n822), .B2(new_n824), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n854), .B1(new_n865), .B2(new_n767), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n471), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n678), .A2(new_n665), .A3(new_n668), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n471), .B1(new_n826), .B2(new_n827), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n722), .A2(G141gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n853), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n853), .B(KEYINPUT58), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(new_n852), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n402), .A3(new_n659), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n868), .A2(new_n658), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  OR3_X1    g682(.A1(new_n810), .A2(new_n883), .A3(new_n630), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n810), .B2(new_n630), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n823), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n863), .B2(new_n864), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n854), .B1(new_n887), .B2(new_n767), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n471), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n886), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n858), .A2(new_n859), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n820), .B1(new_n573), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n698), .B1(new_n893), .B2(KEYINPUT119), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n861), .A2(new_n862), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n827), .B1(new_n896), .B2(new_n604), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n869), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n882), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n881), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n872), .A2(new_n658), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .A3(new_n402), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n880), .B1(new_n906), .B2(new_n908), .ZN(G1345gat));
  OAI21_X1  g708(.A(G155gat), .B1(new_n872), .B2(new_n791), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n604), .A2(new_n395), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n852), .B2(new_n911), .ZN(G1346gat));
  OAI21_X1  g711(.A(G162gat), .B1(new_n872), .B2(new_n630), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n851), .A2(new_n396), .A3(new_n842), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  NOR4_X1   g714(.A1(new_n760), .A2(new_n665), .A3(new_n694), .A4(new_n668), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n850), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(G169gat), .A3(new_n722), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n665), .B1(new_n826), .B2(new_n827), .ZN(new_n920));
  AND4_X1   g719(.A1(new_n471), .A2(new_n920), .A3(new_n386), .A4(new_n506), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n722), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n922), .B2(G169gat), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT124), .ZN(G1348gat));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n220), .A3(new_n659), .ZN(new_n925));
  OAI21_X1  g724(.A(G176gat), .B1(new_n917), .B2(new_n658), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  NAND3_X1  g726(.A1(new_n918), .A2(KEYINPUT125), .A3(new_n701), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n245), .A2(new_n247), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n917), .B2(new_n791), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n921), .A2(new_n231), .A3(new_n604), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n917), .B2(new_n630), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT61), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n249), .A3(new_n698), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1351gat));
  AND4_X1   g738(.A1(new_n694), .A2(new_n920), .A3(new_n386), .A4(new_n678), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n722), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(new_n899), .B2(new_n904), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n889), .B(new_n827), .C1(new_n896), .C2(new_n604), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n694), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n888), .A2(new_n889), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n870), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n869), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT121), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n942), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n665), .A2(new_n668), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n678), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G197gat), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n954), .A2(new_n955), .A3(new_n573), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n941), .B1(new_n952), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n958), .A3(new_n659), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n961), .B2(new_n959), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n678), .A2(new_n659), .A3(new_n953), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n965), .B1(new_n942), .B2(new_n951), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n966), .B2(new_n958), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n940), .A2(new_n351), .A3(new_n604), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n954), .A2(new_n767), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n946), .B2(new_n949), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT63), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(new_n342), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n899), .B2(new_n904), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n940), .B2(new_n698), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n954), .A2(new_n352), .A3(new_n630), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n952), .B2(new_n978), .ZN(G1355gat));
endmodule


