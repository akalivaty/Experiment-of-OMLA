

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U558 ( .A(n642), .B(KEYINPUT98), .ZN(n645) );
  XNOR2_X1 U559 ( .A(KEYINPUT28), .B(n644), .ZN(n524) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n613) );
  AND2_X1 U561 ( .A1(n645), .A2(n524), .ZN(n646) );
  NAND2_X1 U562 ( .A1(n662), .A2(n661), .ZN(n673) );
  XNOR2_X1 U563 ( .A(n671), .B(KEYINPUT32), .ZN(n679) );
  NOR2_X1 U564 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n525), .Z(n800) );
  AND2_X1 U566 ( .A1(n550), .A2(n549), .ZN(G160) );
  INV_X1 U567 ( .A(G651), .ZN(n531) );
  NOR2_X1 U568 ( .A1(G543), .A2(n531), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G63), .A2(n800), .ZN(n528) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n581) );
  NOR2_X1 U571 ( .A1(G651), .A2(n581), .ZN(n526) );
  XNOR2_X1 U572 ( .A(KEYINPUT64), .B(n526), .ZN(n805) );
  NAND2_X1 U573 ( .A1(G51), .A2(n805), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U575 ( .A(KEYINPUT6), .B(n529), .ZN(n537) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n801) );
  NAND2_X1 U577 ( .A1(n801), .A2(G89), .ZN(n530) );
  XNOR2_X1 U578 ( .A(KEYINPUT4), .B(n530), .ZN(n534) );
  NOR2_X1 U579 ( .A1(n581), .A2(n531), .ZN(n804) );
  NAND2_X1 U580 ( .A1(n804), .A2(G76), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT75), .B(n532), .Z(n533) );
  NAND2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U583 ( .A(n535), .B(KEYINPUT5), .Z(n536) );
  NOR2_X1 U584 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U585 ( .A(KEYINPUT7), .B(n538), .Z(n539) );
  XNOR2_X1 U586 ( .A(KEYINPUT76), .B(n539), .ZN(G168) );
  XOR2_X1 U587 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  XOR2_X2 U589 ( .A(KEYINPUT17), .B(n540), .Z(n889) );
  NAND2_X1 U590 ( .A1(n889), .A2(G137), .ZN(n543) );
  AND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U592 ( .A1(n894), .A2(G113), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT65), .B(n541), .Z(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n544), .B(KEYINPUT66), .ZN(n546) );
  INV_X1 U596 ( .A(G2105), .ZN(n547) );
  NOR2_X1 U597 ( .A1(G2104), .A2(n547), .ZN(n895) );
  AND2_X1 U598 ( .A1(n895), .A2(G125), .ZN(n545) );
  NOR2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n550) );
  AND2_X1 U600 ( .A1(n547), .A2(G2104), .ZN(n890) );
  NAND2_X1 U601 ( .A1(G101), .A2(n890), .ZN(n548) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n548), .Z(n549) );
  NAND2_X1 U603 ( .A1(n889), .A2(G138), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G114), .A2(n894), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT87), .B(n551), .Z(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G102), .A2(n890), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G126), .A2(n895), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U610 ( .A1(n557), .A2(n556), .ZN(G164) );
  NAND2_X1 U611 ( .A1(G65), .A2(n800), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G91), .A2(n801), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U614 ( .A1(n804), .A2(G78), .ZN(n561) );
  NAND2_X1 U615 ( .A1(G53), .A2(n805), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U617 ( .A1(n563), .A2(n562), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G90), .A2(n801), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G77), .A2(n804), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U621 ( .A(n566), .B(KEYINPUT9), .ZN(n571) );
  NAND2_X1 U622 ( .A1(G64), .A2(n800), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G52), .A2(n805), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U625 ( .A(KEYINPUT68), .B(n569), .Z(n570) );
  NAND2_X1 U626 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U627 ( .A(n572), .B(KEYINPUT69), .ZN(G171) );
  NAND2_X1 U628 ( .A1(n804), .A2(G75), .ZN(n574) );
  NAND2_X1 U629 ( .A1(G50), .A2(n805), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U631 ( .A1(G62), .A2(n800), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G88), .A2(n801), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U635 ( .A(n579), .B(KEYINPUT83), .ZN(G303) );
  NAND2_X1 U636 ( .A1(n805), .A2(G49), .ZN(n580) );
  XNOR2_X1 U637 ( .A(n580), .B(KEYINPUT82), .ZN(n586) );
  NAND2_X1 U638 ( .A1(G87), .A2(n581), .ZN(n583) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U641 ( .A1(n800), .A2(n584), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G61), .A2(n800), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G86), .A2(n801), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n804), .A2(G73), .ZN(n589) );
  XOR2_X1 U647 ( .A(KEYINPUT2), .B(n589), .Z(n590) );
  NOR2_X1 U648 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U649 ( .A1(G48), .A2(n805), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n593), .A2(n592), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G47), .A2(n805), .ZN(n595) );
  NAND2_X1 U652 ( .A1(n800), .A2(G60), .ZN(n594) );
  NAND2_X1 U653 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U654 ( .A(KEYINPUT67), .B(n596), .ZN(n600) );
  NAND2_X1 U655 ( .A1(G85), .A2(n801), .ZN(n598) );
  NAND2_X1 U656 ( .A1(G72), .A2(n804), .ZN(n597) );
  AND2_X1 U657 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U658 ( .A1(n600), .A2(n599), .ZN(G290) );
  INV_X1 U659 ( .A(G40), .ZN(n601) );
  OR2_X1 U660 ( .A1(n601), .A2(G1384), .ZN(n602) );
  NOR2_X1 U661 ( .A1(G164), .A2(n602), .ZN(n603) );
  NAND2_X1 U662 ( .A1(G160), .A2(n603), .ZN(n635) );
  NAND2_X1 U663 ( .A1(G8), .A2(n635), .ZN(n705) );
  NAND2_X1 U664 ( .A1(G56), .A2(n800), .ZN(n604) );
  XOR2_X1 U665 ( .A(KEYINPUT14), .B(n604), .Z(n610) );
  NAND2_X1 U666 ( .A1(n801), .A2(G81), .ZN(n605) );
  XNOR2_X1 U667 ( .A(n605), .B(KEYINPUT12), .ZN(n607) );
  NAND2_X1 U668 ( .A1(G68), .A2(n804), .ZN(n606) );
  NAND2_X1 U669 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U670 ( .A(KEYINPUT13), .B(n608), .Z(n609) );
  NOR2_X1 U671 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U672 ( .A1(G43), .A2(n805), .ZN(n611) );
  NAND2_X1 U673 ( .A1(n612), .A2(n611), .ZN(n948) );
  INV_X1 U674 ( .A(G1996), .ZN(n920) );
  NOR2_X1 U675 ( .A1(n635), .A2(n920), .ZN(n614) );
  XNOR2_X1 U676 ( .A(n614), .B(n613), .ZN(n616) );
  NAND2_X1 U677 ( .A1(n635), .A2(G1341), .ZN(n615) );
  NAND2_X1 U678 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U679 ( .A1(n948), .A2(n617), .ZN(n628) );
  NAND2_X1 U680 ( .A1(n805), .A2(G54), .ZN(n618) );
  XNOR2_X1 U681 ( .A(n618), .B(KEYINPUT74), .ZN(n625) );
  NAND2_X1 U682 ( .A1(G92), .A2(n801), .ZN(n620) );
  NAND2_X1 U683 ( .A1(G79), .A2(n804), .ZN(n619) );
  NAND2_X1 U684 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U685 ( .A1(G66), .A2(n800), .ZN(n621) );
  XNOR2_X1 U686 ( .A(KEYINPUT73), .B(n621), .ZN(n622) );
  NOR2_X1 U687 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U688 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X2 U689 ( .A(KEYINPUT15), .B(n626), .ZN(n949) );
  NOR2_X1 U690 ( .A1(n628), .A2(n949), .ZN(n627) );
  XNOR2_X1 U691 ( .A(n627), .B(KEYINPUT97), .ZN(n634) );
  NAND2_X1 U692 ( .A1(n628), .A2(n949), .ZN(n632) );
  INV_X1 U693 ( .A(n635), .ZN(n647) );
  NOR2_X1 U694 ( .A1(n647), .A2(G1348), .ZN(n630) );
  NOR2_X1 U695 ( .A1(G2067), .A2(n635), .ZN(n629) );
  NOR2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U698 ( .A1(n634), .A2(n633), .ZN(n641) );
  INV_X1 U699 ( .A(G2072), .ZN(n1000) );
  NOR2_X1 U700 ( .A1(n635), .A2(n1000), .ZN(n637) );
  XNOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n636) );
  XNOR2_X1 U702 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U703 ( .A(n647), .ZN(n663) );
  NAND2_X1 U704 ( .A1(n663), .A2(G1956), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n643) );
  OR2_X1 U706 ( .A1(G299), .A2(n643), .ZN(n640) );
  NAND2_X1 U707 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U708 ( .A1(G299), .A2(n643), .ZN(n644) );
  XNOR2_X1 U709 ( .A(n646), .B(KEYINPUT29), .ZN(n653) );
  NOR2_X1 U710 ( .A1(n647), .A2(G1961), .ZN(n648) );
  XOR2_X1 U711 ( .A(KEYINPUT94), .B(n648), .Z(n651) );
  XOR2_X1 U712 ( .A(G2078), .B(KEYINPUT25), .Z(n918) );
  NOR2_X1 U713 ( .A1(n918), .A2(n663), .ZN(n649) );
  XNOR2_X1 U714 ( .A(KEYINPUT95), .B(n649), .ZN(n650) );
  NAND2_X1 U715 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U716 ( .A1(G171), .A2(n657), .ZN(n652) );
  NAND2_X1 U717 ( .A1(n653), .A2(n652), .ZN(n662) );
  NOR2_X1 U718 ( .A1(G1966), .A2(n705), .ZN(n675) );
  NOR2_X1 U719 ( .A1(G2084), .A2(n663), .ZN(n672) );
  NOR2_X1 U720 ( .A1(n675), .A2(n672), .ZN(n654) );
  NAND2_X1 U721 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U723 ( .A1(G168), .A2(n656), .ZN(n659) );
  NOR2_X1 U724 ( .A1(G171), .A2(n657), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U726 ( .A(KEYINPUT31), .B(n660), .Z(n661) );
  NAND2_X1 U727 ( .A1(n673), .A2(G286), .ZN(n669) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n705), .ZN(n665) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U731 ( .A(KEYINPUT99), .B(n666), .Z(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(G303), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U734 ( .A1(n670), .A2(G8), .ZN(n671) );
  NAND2_X1 U735 ( .A1(G8), .A2(n672), .ZN(n677) );
  INV_X1 U736 ( .A(n673), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n702) );
  NOR2_X1 U740 ( .A1(G288), .A2(G1976), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT100), .ZN(n961) );
  NOR2_X1 U742 ( .A1(G1971), .A2(G303), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n961), .A2(n681), .ZN(n682) );
  AND2_X1 U744 ( .A1(n702), .A2(n682), .ZN(n683) );
  NOR2_X1 U745 ( .A1(n705), .A2(n683), .ZN(n690) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n955) );
  INV_X1 U747 ( .A(KEYINPUT33), .ZN(n692) );
  INV_X1 U748 ( .A(n961), .ZN(n684) );
  OR2_X1 U749 ( .A1(n705), .A2(n684), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n692), .A2(n685), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(KEYINPUT101), .ZN(n691) );
  AND2_X1 U752 ( .A1(n955), .A2(n691), .ZN(n688) );
  XNOR2_X1 U753 ( .A(G1981), .B(G305), .ZN(n945) );
  INV_X1 U754 ( .A(n945), .ZN(n687) );
  AND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n709) );
  INV_X1 U757 ( .A(n691), .ZN(n693) );
  OR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U759 ( .A1(n945), .A2(n694), .ZN(n699) );
  NOR2_X1 U760 ( .A1(G1981), .A2(G305), .ZN(n695) );
  XNOR2_X1 U761 ( .A(n695), .B(KEYINPUT93), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n696), .B(KEYINPUT24), .ZN(n697) );
  OR2_X1 U763 ( .A1(n697), .A2(n705), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n707) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n700) );
  XNOR2_X1 U766 ( .A(n700), .B(KEYINPUT102), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n701), .A2(G8), .ZN(n703) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U771 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n757) );
  XNOR2_X1 U775 ( .A(G1986), .B(KEYINPUT88), .ZN(n712) );
  XNOR2_X1 U776 ( .A(n712), .B(G290), .ZN(n957) );
  NAND2_X1 U777 ( .A1(n757), .A2(n957), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n744) );
  NAND2_X1 U779 ( .A1(n889), .A2(G140), .ZN(n715) );
  XOR2_X1 U780 ( .A(KEYINPUT89), .B(n715), .Z(n717) );
  NAND2_X1 U781 ( .A1(n890), .A2(G104), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n718), .ZN(n724) );
  NAND2_X1 U784 ( .A1(n895), .A2(G128), .ZN(n719) );
  XNOR2_X1 U785 ( .A(n719), .B(KEYINPUT90), .ZN(n721) );
  NAND2_X1 U786 ( .A1(G116), .A2(n894), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U788 ( .A(KEYINPUT35), .B(n722), .Z(n723) );
  NOR2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U790 ( .A(KEYINPUT36), .B(n725), .ZN(n881) );
  XNOR2_X1 U791 ( .A(KEYINPUT37), .B(G2067), .ZN(n755) );
  NOR2_X1 U792 ( .A1(n881), .A2(n755), .ZN(n1021) );
  NAND2_X1 U793 ( .A1(n757), .A2(n1021), .ZN(n753) );
  XOR2_X1 U794 ( .A(n757), .B(KEYINPUT91), .Z(n741) );
  NAND2_X1 U795 ( .A1(G131), .A2(n889), .ZN(n727) );
  NAND2_X1 U796 ( .A1(G119), .A2(n895), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U798 ( .A1(G107), .A2(n894), .ZN(n729) );
  NAND2_X1 U799 ( .A1(G95), .A2(n890), .ZN(n728) );
  NAND2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n886) );
  NAND2_X1 U802 ( .A1(G1991), .A2(n886), .ZN(n740) );
  NAND2_X1 U803 ( .A1(G141), .A2(n889), .ZN(n733) );
  NAND2_X1 U804 ( .A1(G129), .A2(n895), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n890), .A2(G105), .ZN(n734) );
  XOR2_X1 U807 ( .A(KEYINPUT38), .B(n734), .Z(n735) );
  NOR2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U809 ( .A1(n894), .A2(G117), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n903) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n903), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n1012) );
  NAND2_X1 U813 ( .A1(n741), .A2(n1012), .ZN(n746) );
  NAND2_X1 U814 ( .A1(n753), .A2(n746), .ZN(n742) );
  XNOR2_X1 U815 ( .A(KEYINPUT92), .B(n742), .ZN(n743) );
  XNOR2_X1 U816 ( .A(n745), .B(KEYINPUT103), .ZN(n760) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n903), .ZN(n1006) );
  INV_X1 U818 ( .A(n746), .ZN(n749) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n886), .ZN(n1013) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U821 ( .A1(n1013), .A2(n747), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n1006), .A2(n750), .ZN(n751) );
  XNOR2_X1 U824 ( .A(KEYINPUT104), .B(n751), .ZN(n752) );
  XNOR2_X1 U825 ( .A(n752), .B(KEYINPUT39), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n881), .A2(n755), .ZN(n1018) );
  NAND2_X1 U828 ( .A1(n756), .A2(n1018), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U831 ( .A(n761), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U832 ( .A(G2427), .B(G2435), .Z(n763) );
  XNOR2_X1 U833 ( .A(G2454), .B(G2443), .ZN(n762) );
  XNOR2_X1 U834 ( .A(n763), .B(n762), .ZN(n770) );
  XOR2_X1 U835 ( .A(G2451), .B(KEYINPUT105), .Z(n765) );
  XNOR2_X1 U836 ( .A(G2430), .B(G2438), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n765), .B(n764), .ZN(n766) );
  XOR2_X1 U838 ( .A(n766), .B(G2446), .Z(n768) );
  XNOR2_X1 U839 ( .A(G1348), .B(G1341), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n770), .B(n769), .ZN(n771) );
  AND2_X1 U842 ( .A1(n771), .A2(G14), .ZN(G401) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  INV_X1 U845 ( .A(G120), .ZN(G236) );
  INV_X1 U846 ( .A(G132), .ZN(G219) );
  INV_X1 U847 ( .A(G82), .ZN(G220) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U849 ( .A(n772), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n774) );
  INV_X1 U851 ( .A(G223), .ZN(n839) );
  NAND2_X1 U852 ( .A1(G567), .A2(n839), .ZN(n773) );
  XNOR2_X1 U853 ( .A(n774), .B(n773), .ZN(G234) );
  XNOR2_X1 U854 ( .A(G860), .B(KEYINPUT71), .ZN(n780) );
  OR2_X1 U855 ( .A1(n948), .A2(n780), .ZN(G153) );
  XOR2_X1 U856 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U857 ( .A1(G868), .A2(G301), .ZN(n776) );
  OR2_X1 U858 ( .A1(n949), .A2(G868), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(G284) );
  XNOR2_X1 U860 ( .A(KEYINPUT77), .B(G868), .ZN(n777) );
  NOR2_X1 U861 ( .A1(G286), .A2(n777), .ZN(n779) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n781), .A2(n949), .ZN(n782) );
  XNOR2_X1 U866 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U867 ( .A1(n949), .A2(G868), .ZN(n783) );
  NOR2_X1 U868 ( .A1(G559), .A2(n783), .ZN(n784) );
  XNOR2_X1 U869 ( .A(n784), .B(KEYINPUT78), .ZN(n786) );
  NOR2_X1 U870 ( .A1(n948), .A2(G868), .ZN(n785) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(G282) );
  XOR2_X1 U872 ( .A(KEYINPUT18), .B(KEYINPUT80), .Z(n788) );
  NAND2_X1 U873 ( .A1(G123), .A2(n895), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n788), .B(n787), .ZN(n789) );
  XNOR2_X1 U875 ( .A(n789), .B(KEYINPUT79), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n894), .A2(G111), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G135), .A2(n889), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G99), .A2(n890), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n1011) );
  XNOR2_X1 U882 ( .A(n1011), .B(G2096), .ZN(n797) );
  INV_X1 U883 ( .A(G2100), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(G156) );
  NAND2_X1 U885 ( .A1(G559), .A2(n949), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT81), .B(n798), .Z(n818) );
  XNOR2_X1 U887 ( .A(n948), .B(n818), .ZN(n799) );
  NOR2_X1 U888 ( .A1(n799), .A2(G860), .ZN(n810) );
  NAND2_X1 U889 ( .A1(G67), .A2(n800), .ZN(n803) );
  NAND2_X1 U890 ( .A1(G93), .A2(n801), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n809) );
  NAND2_X1 U892 ( .A1(n804), .A2(G80), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G55), .A2(n805), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U895 ( .A1(n809), .A2(n808), .ZN(n820) );
  XOR2_X1 U896 ( .A(n810), .B(n820), .Z(G145) );
  INV_X1 U897 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U898 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n812) );
  XNOR2_X1 U899 ( .A(G299), .B(G166), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n812), .B(n811), .ZN(n815) );
  XOR2_X1 U901 ( .A(G290), .B(n948), .Z(n813) );
  XNOR2_X1 U902 ( .A(G288), .B(n813), .ZN(n814) );
  XNOR2_X1 U903 ( .A(n815), .B(n814), .ZN(n817) );
  XOR2_X1 U904 ( .A(G305), .B(n820), .Z(n816) );
  XNOR2_X1 U905 ( .A(n817), .B(n816), .ZN(n907) );
  XNOR2_X1 U906 ( .A(n818), .B(n907), .ZN(n819) );
  NAND2_X1 U907 ( .A1(n819), .A2(G868), .ZN(n823) );
  INV_X1 U908 ( .A(G868), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2078), .A2(G2084), .ZN(n824) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U916 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U917 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U918 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U919 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U920 ( .A1(G96), .A2(n830), .ZN(n844) );
  AND2_X1 U921 ( .A1(G2106), .A2(n844), .ZN(n836) );
  NOR2_X1 U922 ( .A1(G236), .A2(G237), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G69), .A2(n831), .ZN(n832) );
  XNOR2_X1 U924 ( .A(KEYINPUT85), .B(n832), .ZN(n833) );
  NAND2_X1 U925 ( .A1(n833), .A2(G108), .ZN(n843) );
  NAND2_X1 U926 ( .A1(G567), .A2(n843), .ZN(n834) );
  XOR2_X1 U927 ( .A(KEYINPUT86), .B(n834), .Z(n835) );
  NOR2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G319) );
  INV_X1 U929 ( .A(G319), .ZN(n838) );
  NAND2_X1 U930 ( .A1(G483), .A2(G661), .ZN(n837) );
  NOR2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n842) );
  NAND2_X1 U932 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U935 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G188) );
  NOR2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G325) );
  XOR2_X1 U939 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U941 ( .A(G108), .ZN(G238) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2084), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n847), .B(G2100), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT107), .B(G2678), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U953 ( .A(G2474), .B(G1976), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1956), .B(G1971), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(n856), .B(KEYINPUT108), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(G1981), .B(G1961), .Z(n860) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1966), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G124), .A2(n895), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n894), .A2(G112), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G136), .A2(n889), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G100), .A2(n890), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U973 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(n885) );
  NAND2_X1 U976 ( .A1(G139), .A2(n889), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G103), .A2(n890), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G115), .A2(n894), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G127), .A2(n895), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n999) );
  XNOR2_X1 U984 ( .A(n881), .B(n999), .ZN(n883) );
  XNOR2_X1 U985 ( .A(G160), .B(G164), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n886), .B(n1011), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n905) );
  NAND2_X1 U990 ( .A1(G142), .A2(n889), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G106), .A2(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(KEYINPUT45), .ZN(n900) );
  NAND2_X1 U994 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U995 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(KEYINPUT110), .B(n898), .Z(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n901), .B(G162), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n903), .B(n902), .Z(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U1003 ( .A(n949), .B(n907), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G286), .B(n908), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(G171), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n911), .B(KEYINPUT49), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n912), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT113), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1016 ( .A(G2090), .B(G35), .Z(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT115), .B(n917), .ZN(n933) );
  XNOR2_X1 U1018 ( .A(G27), .B(n918), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(KEYINPUT117), .ZN(n928) );
  XOR2_X1 U1020 ( .A(G2067), .B(G26), .Z(n922) );
  XNOR2_X1 U1021 ( .A(n920), .B(G32), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n926) );
  XOR2_X1 U1023 ( .A(G1991), .B(G25), .Z(n923) );
  NAND2_X1 U1024 ( .A1(n923), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(KEYINPUT53), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(KEYINPUT118), .B(n934), .ZN(n937) );
  XOR2_X1 U1033 ( .A(G2084), .B(G34), .Z(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(n935), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(KEYINPUT119), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT55), .B(n939), .Z(n941) );
  XNOR2_X1 U1038 ( .A(G29), .B(KEYINPUT120), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n942), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n943), .A2(G11), .ZN(n997) );
  XNOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .ZN(n968) );
  XOR2_X1 U1043 ( .A(G168), .B(G1966), .Z(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n946), .Z(n966) );
  XNOR2_X1 U1046 ( .A(G171), .B(G1961), .ZN(n953) );
  XOR2_X1 U1047 ( .A(G1341), .B(KEYINPUT123), .Z(n947) );
  XNOR2_X1 U1048 ( .A(n948), .B(n947), .ZN(n951) );
  XOR2_X1 U1049 ( .A(G1348), .B(n949), .Z(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(G166), .B(G1971), .ZN(n959) );
  XOR2_X1 U1053 ( .A(G1956), .B(G299), .Z(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT122), .B(n962), .Z(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n995) );
  INV_X1 U1062 ( .A(G16), .ZN(n993) );
  XOR2_X1 U1063 ( .A(G1986), .B(G24), .Z(n970) );
  XOR2_X1 U1064 ( .A(G1971), .B(G22), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G23), .B(G1976), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1068 ( .A(KEYINPUT58), .B(n973), .Z(n989) );
  XOR2_X1 U1069 ( .A(G1961), .B(G5), .Z(n984) );
  XOR2_X1 U1070 ( .A(G1981), .B(G6), .Z(n977) );
  XNOR2_X1 U1071 ( .A(G1956), .B(G20), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(G19), .B(G1341), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(n978), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT59), .B(G1348), .Z(n979) );
  XNOR2_X1 U1077 ( .A(G4), .B(n979), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(KEYINPUT60), .B(n982), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(G21), .B(G1966), .ZN(n985) );
  NOR2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(KEYINPUT125), .B(n987), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(n990), .B(KEYINPUT61), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(n991), .B(KEYINPUT126), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(n998), .B(KEYINPUT127), .ZN(n1027) );
  INV_X1 U1091 ( .A(G29), .ZN(n1025) );
  XNOR2_X1 U1092 ( .A(n999), .B(KEYINPUT114), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(n1000), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1004), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1007), .Z(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(G2084), .B(G160), .Z(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1022), .Z(n1023) );
  NOR2_X1 U1109 ( .A1(KEYINPUT55), .A2(n1023), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

