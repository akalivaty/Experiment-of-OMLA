//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  AOI21_X1  g003(.A(G8gat), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n206), .A2(new_n207), .A3(G1gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n202), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n203), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n210), .B(new_n203), .C1(new_n204), .C2(G8gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  OR3_X1    g014(.A1(new_n215), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT88), .B(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G43gat), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G43gat), .A2(G50gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT15), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n221), .B2(new_n222), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT89), .B(G43gat), .Z(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n222), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n225), .B1(new_n230), .B2(new_n220), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT17), .B1(new_n226), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n214), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(new_n231), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n214), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n235), .A2(new_n238), .A3(KEYINPUT18), .A4(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(KEYINPUT13), .Z(new_n241));
  INV_X1    g040(.A(new_n214), .ZN(new_n242));
  INV_X1    g041(.A(new_n236), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(new_n244), .B2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n232), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n237), .B1(new_n249), .B2(new_n214), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT18), .B1(new_n250), .B2(new_n239), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n240), .A2(new_n245), .A3(KEYINPUT92), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT11), .B(G169gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT12), .Z(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n253), .B(new_n258), .C1(new_n246), .C2(new_n251), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n260), .A2(KEYINPUT93), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT93), .B1(new_n260), .B2(new_n261), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT0), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT78), .B(G141gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G148gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n274));
  INV_X1    g073(.A(G141gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(G148gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277));
  OR2_X1    g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(KEYINPUT2), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n276), .B(new_n279), .C1(new_n274), .C2(new_n273), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(KEYINPUT76), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n281), .A2(new_n277), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n275), .A2(G148gat), .ZN(new_n283));
  INV_X1    g082(.A(G148gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G141gat), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n283), .A2(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n282), .B(new_n288), .C1(KEYINPUT76), .C2(new_n278), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(KEYINPUT69), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(KEYINPUT69), .B2(new_n293), .ZN(new_n295));
  XOR2_X1   g094(.A(G127gat), .B(G134gat), .Z(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT68), .B(G120gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G113gat), .A2(G120gat), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT1), .B1(new_n291), .B2(new_n292), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n296), .A2(KEYINPUT67), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(KEYINPUT67), .B2(new_n296), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n280), .A2(new_n300), .A3(new_n289), .A4(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n271), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n313));
  INV_X1    g112(.A(new_n290), .ZN(new_n314));
  INV_X1    g113(.A(new_n305), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT80), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT80), .B1(new_n307), .B2(KEYINPUT4), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n280), .A2(new_n323), .A3(new_n289), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n305), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n309), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n313), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT81), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n312), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n307), .B(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n332), .A3(new_n271), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n270), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n321), .A2(new_n313), .A3(new_n326), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT81), .B1(new_n328), .B2(new_n329), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n311), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n269), .A3(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(KEYINPUT6), .B(new_n270), .C1(new_n331), .C2(new_n334), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT23), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT65), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT23), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n349), .A2(KEYINPUT65), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT64), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n360));
  INV_X1    g159(.A(G183gat), .ZN(new_n361));
  INV_X1    g160(.A(G190gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(KEYINPUT64), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT25), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n349), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n358), .B2(new_n363), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT26), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n351), .A2(KEYINPUT66), .A3(KEYINPUT26), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n348), .B2(new_n370), .ZN(new_n373));
  OAI221_X1 g172(.A(new_n352), .B1(new_n370), .B2(new_n348), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n362), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n376), .A2(KEYINPUT28), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n376), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n368), .ZN(new_n382));
  INV_X1    g181(.A(new_n379), .ZN(new_n383));
  INV_X1    g182(.A(new_n380), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n382), .A2(new_n383), .B1(KEYINPUT29), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g186(.A1(G211gat), .A2(G218gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT22), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(G197gat), .A2(G204gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(G197gat), .A2(G204gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n387), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G211gat), .B(G218gat), .Z(new_n396));
  OAI21_X1  g195(.A(KEYINPUT72), .B1(new_n396), .B2(KEYINPUT73), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n395), .A2(new_n396), .B1(new_n397), .B2(new_n393), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n385), .A3(new_n398), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(KEYINPUT74), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n403), .A3(new_n399), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n347), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OR3_X1    g204(.A1(new_n405), .A2(KEYINPUT75), .A3(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n404), .A3(new_n347), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT30), .B1(new_n405), .B2(KEYINPUT75), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n398), .B1(new_n324), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT3), .B1(new_n398), .B2(new_n410), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n413), .C1(new_n314), .C2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n396), .B1(new_n393), .B2(KEYINPUT82), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(KEYINPUT82), .B2(new_n393), .ZN(new_n417));
  INV_X1    g216(.A(new_n396), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT82), .A3(new_n393), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n410), .ZN(new_n420));
  OR3_X1    g219(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT83), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT83), .B1(new_n417), .B2(new_n420), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n323), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n411), .B1(new_n423), .B2(new_n290), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n415), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G22gat), .ZN(new_n426));
  INV_X1    g225(.A(G22gat), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n415), .B(new_n427), .C1(new_n413), .C2(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n425), .B2(G22gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT31), .B(G50gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n426), .A2(new_n430), .A3(new_n428), .A4(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G227gat), .ZN(new_n440));
  INV_X1    g239(.A(G233gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n369), .A2(new_n305), .A3(new_n379), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n315), .B1(new_n382), .B2(new_n383), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT34), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n445), .A2(KEYINPUT71), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n445), .B2(KEYINPUT71), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT70), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n443), .A2(new_n442), .A3(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT32), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G15gat), .B(G43gat), .Z(new_n455));
  XNOR2_X1  g254(.A(G71gat), .B(G99gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n457), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n451), .B(KEYINPUT32), .C1(new_n453), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n450), .B(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n343), .A2(new_n409), .A3(new_n439), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n461), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n447), .A2(new_n458), .A3(new_n460), .A4(new_n448), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n438), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n343), .A3(new_n409), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT87), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n469), .A2(new_n343), .A3(new_n409), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n407), .B1(new_n475), .B2(new_n346), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n400), .A2(new_n477), .A3(new_n401), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n398), .B1(new_n381), .B2(new_n385), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n479), .B2(KEYINPUT85), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT38), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(KEYINPUT86), .A3(new_n481), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n402), .A2(new_n404), .A3(KEYINPUT37), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n405), .B1(new_n488), .B2(KEYINPUT38), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n486), .A2(new_n342), .A3(new_n341), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n309), .B1(new_n332), .B2(new_n325), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT39), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n270), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT39), .B1(new_n308), .B2(new_n310), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n493), .B(KEYINPUT40), .C1(new_n491), .C2(new_n494), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n335), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n406), .A2(new_n408), .A3(new_n407), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n438), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n343), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n438), .B1(new_n503), .B2(new_n500), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT36), .B1(new_n465), .B2(new_n467), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n462), .B2(KEYINPUT36), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n265), .B1(new_n474), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G71gat), .A2(G78gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G71gat), .ZN(new_n513));
  INV_X1    g312(.A(G78gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G57gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G64gat), .ZN(new_n519));
  INV_X1    g318(.A(G64gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G57gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT9), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n510), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n517), .A2(KEYINPUT95), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n512), .A2(new_n515), .A3(new_n526), .A4(new_n516), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n510), .B1(new_n515), .B2(new_n523), .ZN(new_n528));
  OR3_X1    g327(.A1(new_n520), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(KEYINPUT96), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n521), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n525), .A2(new_n527), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  INV_X1    g334(.A(G127gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n242), .B1(KEYINPUT21), .B2(new_n532), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT97), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G155gat), .ZN(new_n542));
  XOR2_X1   g341(.A(G183gat), .B(G211gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n539), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(G85gat), .A3(G92gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G99gat), .ZN(new_n560));
  INV_X1    g359(.A(G106gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT8), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n553), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G99gat), .B(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n553), .A2(new_n559), .A3(new_n564), .A4(new_n562), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(KEYINPUT99), .A3(new_n565), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT100), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT100), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(G99gat), .B2(G106gat), .ZN(new_n574));
  AND2_X1   g373(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n577), .B2(new_n557), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n564), .B1(new_n578), .B2(new_n553), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n568), .A2(new_n567), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n570), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n249), .A2(new_n571), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n569), .A2(KEYINPUT100), .A3(new_n570), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT100), .B1(new_n569), .B2(new_n570), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n243), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n584), .A2(new_n586), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n585), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n591), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n593), .A2(new_n596), .B1(new_n599), .B2(new_n591), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n548), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n525), .A2(new_n527), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n531), .A2(new_n528), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n581), .B2(new_n582), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n568), .B1(new_n566), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT102), .B1(new_n563), .B2(new_n565), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n532), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT10), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n532), .A2(KEYINPUT10), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n583), .B2(new_n571), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n605), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n605), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n609), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  OR2_X1    g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n617), .A2(new_n625), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n509), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n503), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n474), .A2(new_n508), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(new_n500), .A3(new_n264), .A4(new_n629), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT16), .B(G8gat), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT42), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n637), .A2(KEYINPUT104), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT104), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT105), .B1(new_n635), .B2(G8gat), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n635), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n643));
  OAI22_X1  g442(.A1(new_n642), .A2(new_n643), .B1(new_n637), .B2(new_n638), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n633), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n646), .B(KEYINPUT106), .C1(new_n640), .C2(new_n639), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(G1325gat));
  AND2_X1   g447(.A1(new_n465), .A2(new_n467), .ZN(new_n649));
  AOI21_X1  g448(.A(G15gat), .B1(new_n630), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT107), .Z(new_n651));
  AND2_X1   g450(.A1(new_n506), .A2(G15gat), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n630), .B2(new_n652), .ZN(G1326gat));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n438), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  NOR2_X1   g455(.A1(new_n548), .A2(new_n628), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n603), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n509), .A2(new_n503), .A3(new_n218), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT45), .ZN(new_n661));
  INV_X1    g460(.A(new_n603), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n634), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  AOI211_X1 g463(.A(new_n664), .B(new_n603), .C1(new_n474), .C2(new_n508), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n260), .A2(new_n261), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n658), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n343), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n661), .B1(new_n671), .B2(new_n218), .ZN(G1328gat));
  NAND2_X1  g471(.A1(new_n509), .A2(new_n659), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(G36gat), .A3(new_n409), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT46), .ZN(new_n675));
  OAI21_X1  g474(.A(G36gat), .B1(new_n670), .B2(new_n409), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1329gat));
  INV_X1    g476(.A(new_n649), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n229), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n507), .A2(new_n229), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n670), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n509), .B2(new_n659), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n634), .A2(new_n683), .A3(new_n264), .A4(new_n659), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n439), .A2(G50gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI22_X1  g488(.A1(KEYINPUT35), .A2(new_n463), .B1(new_n470), .B2(KEYINPUT87), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n506), .B1(new_n490), .B2(new_n501), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n690), .A2(new_n473), .B1(new_n691), .B2(new_n504), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n664), .B1(new_n692), .B2(new_n603), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n634), .A2(KEYINPUT44), .A3(new_n662), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n438), .A3(new_n694), .A4(new_n669), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n685), .A2(new_n689), .B1(new_n695), .B2(G50gat), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT48), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n222), .B1(new_n695), .B2(KEYINPUT109), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n666), .A2(new_n700), .A3(new_n438), .A4(new_n669), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT48), .B1(new_n688), .B2(new_n684), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n698), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g504(.A(KEYINPUT110), .B(new_n703), .C1(new_n699), .C2(new_n701), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n697), .B1(new_n705), .B2(new_n706), .ZN(G1331gat));
  INV_X1    g506(.A(new_n628), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n604), .A2(new_n667), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n634), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n343), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n518), .ZN(G1332gat));
  AOI211_X1 g511(.A(new_n409), .B(new_n710), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n710), .B2(new_n507), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n649), .A2(new_n513), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g518(.A1(new_n710), .A2(new_n439), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n514), .ZN(G1335gat));
  NOR3_X1   g520(.A1(new_n548), .A2(new_n667), .A3(new_n708), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n666), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723), .B2(new_n343), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n548), .A2(new_n667), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n634), .A2(new_n662), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n343), .A2(G85gat), .A3(new_n708), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT111), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n731), .ZN(G1336gat));
  NAND4_X1  g531(.A1(new_n693), .A2(new_n500), .A3(new_n694), .A4(new_n722), .ZN(new_n733));
  INV_X1    g532(.A(new_n577), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT113), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(KEYINPUT52), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n500), .A2(new_n555), .A3(new_n628), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT112), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n728), .A2(new_n738), .B1(new_n733), .B2(new_n734), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n736), .B(new_n739), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n723), .B2(new_n507), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n728), .A2(new_n560), .A3(new_n649), .A4(new_n628), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1338gat));
  OAI21_X1  g542(.A(G106gat), .B1(new_n723), .B2(new_n439), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n561), .A3(new_n438), .A4(new_n628), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n748), .A3(KEYINPUT53), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n744), .B(new_n745), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1339gat));
  AND2_X1   g551(.A1(new_n546), .A2(new_n547), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT10), .ZN(new_n754));
  INV_X1    g553(.A(new_n568), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n579), .B2(KEYINPUT102), .ZN(new_n756));
  INV_X1    g555(.A(new_n612), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n608), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n532), .B1(new_n569), .B2(new_n570), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n615), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n587), .B2(new_n588), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n618), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n623), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n760), .A2(new_n762), .A3(new_n618), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n617), .A2(KEYINPUT54), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n765), .A2(new_n767), .A3(KEYINPUT55), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n627), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n768), .A2(new_n774), .A3(new_n769), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n771), .A2(new_n773), .A3(new_n667), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n246), .A2(new_n251), .A3(new_n258), .ZN(new_n777));
  INV_X1    g576(.A(new_n257), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n250), .A2(new_n239), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n244), .A2(new_n237), .A3(new_n241), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n628), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n662), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n771), .A2(new_n773), .A3(new_n775), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n601), .B2(new_n602), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n753), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n548), .A2(new_n668), .A3(new_n603), .A4(new_n708), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n343), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND4_X1   g589(.A1(new_n439), .A2(new_n790), .A3(new_n409), .A4(new_n462), .ZN(new_n791));
  AOI21_X1  g590(.A(G113gat), .B1(new_n791), .B2(new_n667), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n789), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n439), .ZN(new_n795));
  AOI211_X1 g594(.A(KEYINPUT116), .B(new_n438), .C1(new_n788), .C2(new_n789), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n503), .A2(new_n797), .A3(new_n409), .A4(new_n649), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n265), .A2(new_n291), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n792), .B1(new_n798), .B2(new_n799), .ZN(G1340gat));
  NAND3_X1  g599(.A1(new_n791), .A2(new_n299), .A3(new_n628), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n628), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n803), .B2(new_n292), .ZN(G1341gat));
  NAND3_X1  g603(.A1(new_n791), .A2(new_n536), .A3(new_n548), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n548), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n807), .B2(new_n536), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n809), .A3(new_n662), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT56), .Z(new_n811));
  NAND2_X1  g610(.A1(new_n798), .A2(new_n662), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n809), .ZN(G1343gat));
  XNOR2_X1  g613(.A(new_n783), .B(KEYINPUT117), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n768), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n768), .A2(new_n816), .ZN(new_n818));
  XOR2_X1   g617(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n264), .B(new_n773), .C1(new_n817), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n662), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n753), .B1(new_n822), .B2(new_n787), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n789), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT57), .B1(new_n824), .B2(new_n439), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n439), .B1(new_n788), .B2(new_n789), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n506), .A2(new_n343), .A3(new_n500), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n825), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n272), .B1(new_n830), .B2(new_n667), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n438), .A2(new_n790), .A3(new_n409), .A4(new_n507), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n832), .A2(new_n275), .A3(new_n264), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT58), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n272), .B1(new_n830), .B2(new_n264), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n833), .A2(KEYINPUT58), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(G1344gat));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n284), .A3(new_n628), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n629), .A2(new_n265), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n439), .B1(new_n823), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT57), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n826), .A2(KEYINPUT57), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n841), .B2(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n829), .A2(new_n847), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n846), .A2(new_n628), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n839), .B1(new_n850), .B2(G148gat), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT59), .B(new_n284), .C1(new_n830), .C2(new_n628), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n838), .B1(new_n851), .B2(new_n852), .ZN(G1345gat));
  INV_X1    g652(.A(G155gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n832), .A2(new_n854), .A3(new_n548), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n830), .A2(new_n548), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n854), .ZN(G1346gat));
  AOI21_X1  g656(.A(G162gat), .B1(new_n832), .B2(new_n662), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n662), .A2(G162gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n830), .B2(new_n859), .ZN(G1347gat));
  AOI21_X1  g659(.A(new_n503), .B1(new_n788), .B2(new_n789), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n439), .A2(new_n462), .A3(new_n500), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(G169gat), .B1(new_n867), .B2(new_n667), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n343), .A2(new_n500), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n678), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n795), .B2(new_n796), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT123), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(new_n870), .C1(new_n795), .C2(new_n796), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(G169gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(new_n265), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n868), .A2(new_n877), .ZN(G1348gat));
  OAI21_X1  g677(.A(G176gat), .B1(new_n875), .B2(new_n708), .ZN(new_n879));
  INV_X1    g678(.A(G176gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n867), .A2(new_n880), .A3(new_n628), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1349gat));
  OAI21_X1  g681(.A(G183gat), .B1(new_n875), .B2(new_n753), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n375), .A3(new_n548), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n872), .A2(new_n662), .A3(new_n874), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G190gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT61), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT125), .B1(new_n888), .B2(KEYINPUT61), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n887), .A2(new_n894), .A3(new_n895), .A4(G190gat), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n867), .A2(new_n362), .A3(new_n662), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1351gat));
  NAND3_X1  g698(.A1(new_n507), .A2(new_n438), .A3(new_n500), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n865), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT126), .Z(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n667), .ZN(new_n903));
  INV_X1    g702(.A(G197gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n869), .A2(new_n506), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n846), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n265), .A2(new_n904), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n903), .A2(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n628), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G204gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911));
  AOI21_X1  g710(.A(G204gat), .B1(new_n911), .B2(KEYINPUT62), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n901), .A2(new_n628), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(KEYINPUT62), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n915), .ZN(G1353gat));
  INV_X1    g715(.A(G211gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n917), .A3(new_n548), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n846), .A2(new_n548), .A3(new_n905), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n923), .A3(new_n662), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n906), .A2(new_n662), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n923), .ZN(G1355gat));
endmodule


