//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT68), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  AND2_X1   g049(.A1(new_n465), .A2(G136), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT70), .Z(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n475), .B(new_n479), .C1(G124), .C2(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT71), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n484), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AND4_X1   g065(.A1(G126), .A2(new_n461), .A3(new_n463), .A4(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n477), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n480), .A2(new_n495), .A3(G138), .A4(new_n477), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT6), .B1(new_n506), .B2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n506), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n512), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND2_X1  g091(.A1(new_n511), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n507), .A2(new_n510), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(G543), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n511), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n525), .B1(new_n504), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n522), .A2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n521), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n501), .A2(new_n503), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n511), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(G90), .A2(new_n534), .B1(new_n537), .B2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(new_n521), .A2(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n533), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(G81), .A2(new_n534), .B1(new_n544), .B2(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND4_X1  g128(.A1(new_n517), .A2(G53), .A3(G543), .A4(new_n519), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n500), .B1(new_n511), .B2(KEYINPUT73), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n557), .A2(new_n558), .A3(G53), .A4(new_n519), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n556), .B1(new_n555), .B2(new_n559), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n534), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n533), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n562), .A2(new_n569), .ZN(G299));
  AND3_X1   g145(.A1(new_n532), .A2(KEYINPUT77), .A3(new_n538), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT77), .B1(new_n532), .B2(new_n538), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G301));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n506), .B1(new_n533), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n534), .B2(G87), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n557), .A2(G49), .A3(new_n519), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n533), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n507), .A2(new_n510), .ZN(new_n583));
  AND2_X1   g158(.A1(G48), .A2(G543), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n582), .A2(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n534), .A2(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n521), .A2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n533), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(G85), .A2(new_n534), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n534), .A2(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n533), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n595), .B1(G651), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n521), .A2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n573), .B2(new_n602), .ZN(G284));
  XNOR2_X1  g179(.A(G284), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  XOR2_X1   g181(.A(G299), .B(KEYINPUT79), .Z(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(new_n601), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n601), .A2(G559), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n613), .A2(KEYINPUT80), .A3(new_n602), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT80), .B1(new_n613), .B2(new_n602), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n547), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n482), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n465), .A2(G135), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  INV_X1    g195(.A(G111), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n620), .A2(KEYINPUT82), .B1(new_n621), .B2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(KEYINPUT82), .B2(new_n620), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT83), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n480), .A2(new_n466), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT81), .B(G2100), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G14), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n642), .B2(new_n645), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n653), .B(KEYINPUT17), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n652), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n652), .A2(new_n653), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n662), .B(new_n655), .C1(new_n659), .C2(new_n652), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n672), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  OAI221_X1 g251(.A(new_n673), .B1(new_n668), .B2(new_n671), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n675), .ZN(new_n678));
  INV_X1    g253(.A(G1991), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(G1996), .ZN(new_n685));
  INV_X1    g260(.A(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  AND3_X1   g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n684), .B2(new_n687), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(G229));
  OR2_X1    g266(.A1(G16), .A2(G22), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(G303), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT91), .B(G1971), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n693), .A2(G6), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G305), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NOR4_X1   g278(.A1(new_n697), .A2(new_n698), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  NOR2_X1   g280(.A1(G288), .A2(KEYINPUT90), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n577), .B2(new_n578), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n705), .B1(new_n709), .B2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n704), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT34), .Z(new_n715));
  NOR2_X1   g290(.A1(G25), .A2(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n465), .A2(G131), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n477), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n482), .B2(G119), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT88), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(G29), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n723), .B(new_n725), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n693), .A2(G24), .ZN(new_n727));
  INV_X1    g302(.A(G290), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n693), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G1986), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n729), .A2(G1986), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n715), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(KEYINPUT92), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G20), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  MUX2_X1   g314(.A(new_n738), .B(new_n739), .S(KEYINPUT23), .Z(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT99), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT98), .B(G1956), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n693), .A2(G4), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n610), .B2(new_n693), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT93), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G1348), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G33), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n465), .A2(G139), .ZN(new_n752));
  INV_X1    g327(.A(new_n466), .ZN(new_n753));
  INV_X1    g328(.A(G103), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT25), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n753), .A2(KEYINPUT25), .A3(new_n754), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  INV_X1    g333(.A(G127), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n464), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(G2105), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n751), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G2072), .ZN(new_n764));
  INV_X1    g339(.A(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n765), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT29), .B(G2090), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n763), .A2(G2072), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n765), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n765), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2078), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n764), .A2(new_n769), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G32), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n465), .A2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n466), .A2(G105), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n482), .B2(G129), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT30), .B(G28), .ZN(new_n785));
  OR2_X1    g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  NAND2_X1  g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n785), .A2(new_n765), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n784), .B(new_n788), .C1(new_n765), .C2(new_n625), .ZN(new_n789));
  AND2_X1   g364(.A1(KEYINPUT24), .A2(G34), .ZN(new_n790));
  NOR2_X1   g365(.A1(KEYINPUT24), .A2(G34), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n765), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G160), .B2(G29), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n789), .B1(G2084), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n693), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n693), .ZN(new_n801));
  INV_X1    g376(.A(G1961), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n749), .A2(new_n774), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n765), .A2(G26), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n465), .A2(G140), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n477), .A2(G116), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n482), .B2(G128), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n805), .B1(new_n810), .B2(new_n765), .ZN(new_n811));
  MUX2_X1   g386(.A(new_n805), .B(new_n811), .S(KEYINPUT28), .Z(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(G2067), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(G2067), .ZN(new_n814));
  INV_X1    g389(.A(G2084), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n797), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n693), .A2(G19), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n546), .B2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1341), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n693), .A2(G21), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G168), .B2(new_n693), .ZN(new_n822));
  INV_X1    g397(.A(G1966), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n816), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n748), .A2(G1348), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n804), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AND4_X1   g402(.A1(new_n736), .A2(new_n744), .A3(new_n745), .A4(new_n827), .ZN(G311));
  NAND4_X1  g403(.A1(new_n736), .A2(new_n744), .A3(new_n745), .A4(new_n827), .ZN(G150));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n533), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(G93), .A2(new_n534), .B1(new_n832), .B2(G651), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n520), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NOR2_X1   g414(.A1(new_n601), .A2(new_n611), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n546), .B(new_n837), .Z(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n842), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n839), .B1(new_n844), .B2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n810), .B(new_n781), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n494), .A2(new_n496), .ZN(new_n850));
  INV_X1    g425(.A(G126), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n477), .B1(new_n486), .B2(new_n488), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n481), .A2(new_n851), .B1(new_n852), .B2(new_n484), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n492), .A2(new_n497), .A3(KEYINPUT100), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n848), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n761), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n465), .A2(G142), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n477), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G130), .B2(new_n482), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n721), .B(new_n865), .Z(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT101), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n628), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(KEYINPUT101), .ZN(new_n869));
  INV_X1    g444(.A(new_n628), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n860), .B1(new_n872), .B2(KEYINPUT102), .ZN(new_n873));
  XNOR2_X1  g448(.A(G160), .B(G162), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(new_n625), .Z(new_n875));
  NAND3_X1  g450(.A1(new_n859), .A2(new_n868), .A3(new_n871), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(KEYINPUT102), .ZN(new_n877));
  INV_X1    g452(.A(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n859), .B1(new_n868), .B2(new_n871), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n837), .A2(new_n602), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n706), .A2(new_n708), .ZN(new_n886));
  XNOR2_X1  g461(.A(G290), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G303), .B(G305), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n887), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT104), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n546), .B(new_n837), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n613), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n610), .A2(G299), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n601), .A2(new_n569), .A3(new_n562), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n896), .A2(KEYINPUT103), .A3(new_n897), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n903), .B2(new_n895), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n893), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n885), .B1(new_n905), .B2(new_n602), .ZN(G295));
  OAI21_X1  g481(.A(new_n885), .B1(new_n905), .B2(new_n602), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n896), .A2(new_n897), .ZN(new_n909));
  OAI21_X1  g484(.A(G168), .B1(new_n571), .B2(new_n572), .ZN(new_n910));
  NAND2_X1  g485(.A1(G171), .A2(G286), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n843), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(new_n894), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n909), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n894), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n912), .B(new_n917), .C1(new_n899), .C2(new_n898), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n890), .A2(new_n891), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n882), .ZN(new_n921));
  INV_X1    g496(.A(new_n891), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n887), .A2(new_n889), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n890), .B2(new_n891), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n916), .B2(new_n918), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n908), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  OAI22_X1  g504(.A1(new_n913), .A2(new_n915), .B1(new_n902), .B2(new_n901), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n918), .ZN(new_n931));
  INV_X1    g506(.A(new_n927), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n882), .A4(new_n920), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT44), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n921), .B2(new_n928), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n933), .A2(new_n908), .A3(new_n882), .A4(new_n920), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(G397));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n856), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT106), .B(G40), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n467), .A2(new_n471), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n721), .B(new_n725), .Z(new_n950));
  XNOR2_X1  g525(.A(new_n810), .B(G2067), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n781), .B(G1996), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1986), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n728), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G303), .A2(G8), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT55), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n492), .A2(KEYINPUT100), .A3(new_n497), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT100), .B1(new_n492), .B2(new_n497), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT45), .B(new_n943), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT107), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n856), .A2(new_n966), .A3(KEYINPUT45), .A4(new_n943), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n467), .A2(new_n471), .A3(new_n946), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n498), .A2(new_n943), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(new_n945), .ZN(new_n971));
  AOI21_X1  g546(.A(G1971), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n492), .B2(new_n497), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n969), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT109), .B(G2090), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(G8), .B(new_n961), .C1(new_n972), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n947), .B1(KEYINPUT45), .B2(new_n973), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n965), .B2(new_n967), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n989), .B2(G1971), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(KEYINPUT110), .A3(G8), .A4(new_n961), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n970), .A2(new_n969), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(G1976), .B1(new_n706), .B2(new_n708), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(G288), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(G305), .B2(G1981), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n585), .A2(KEYINPUT111), .A3(new_n1005), .A4(new_n586), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT112), .B(G86), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n534), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n585), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(KEYINPUT113), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1004), .A2(new_n1006), .B1(G1981), .B2(new_n1010), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n947), .A2(new_n973), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1016), .B2(KEYINPUT49), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1002), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n947), .B1(new_n974), .B2(new_n973), .ZN(new_n1023));
  INV_X1    g598(.A(new_n975), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n981), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n972), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1022), .B1(new_n960), .B2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n992), .A2(KEYINPUT124), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT124), .B1(new_n992), .B2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2078), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n968), .A2(new_n1031), .A3(new_n971), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1961), .B1(new_n979), .B2(new_n980), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT53), .B(new_n1031), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1038), .B2(new_n1037), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n854), .B2(new_n855), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n968), .B(new_n1040), .C1(KEYINPUT45), .C2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1036), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT125), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1046), .A3(G171), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n970), .A2(new_n945), .ZN(new_n1049));
  NOR4_X1   g624(.A1(new_n988), .A2(new_n1049), .A3(new_n1033), .A4(G2078), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1050), .B(new_n1035), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1051), .B2(G301), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1034), .A2(G301), .A3(new_n1036), .A4(new_n1042), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1051), .B2(G301), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n823), .B1(new_n988), .B2(new_n1049), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n973), .A2(new_n977), .A3(new_n974), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n977), .B1(new_n973), .B2(new_n974), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n980), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1059), .B2(G2084), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(KEYINPUT122), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n979), .A2(new_n815), .A3(new_n980), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1056), .ZN(new_n1067));
  AOI21_X1  g642(.A(G286), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1062), .A2(new_n995), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1063), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1060), .A2(KEYINPUT122), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1066), .B1(new_n1065), .B2(new_n1056), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G286), .A2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1055), .A2(new_n1048), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n966), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n964), .A2(KEYINPUT107), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n971), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT116), .B(G1956), .Z(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT57), .B(new_n569), .C1(new_n560), .C2(new_n561), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n555), .A2(new_n559), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n569), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n568), .B1(new_n555), .B2(new_n559), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1093), .A2(new_n1094), .A3(KEYINPUT57), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1088), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1083), .A2(new_n1087), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1079), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1083), .A2(new_n1087), .A3(new_n1096), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1088), .B(KEYINPUT118), .C1(new_n1092), .C2(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1086), .B1(new_n989), .B2(new_n1080), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT61), .B(new_n1100), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1018), .A2(G2067), .ZN(new_n1108));
  INV_X1    g683(.A(G1348), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1059), .B2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT60), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n601), .B1(new_n1110), .B2(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT121), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT120), .B(G1996), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n989), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT58), .B(G1341), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n994), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n547), .B(new_n1116), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n989), .B2(new_n1117), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1122), .A2(new_n546), .B1(KEYINPUT121), .B2(new_n1115), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1114), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1107), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1348), .B1(new_n979), .B2(new_n980), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n610), .B1(new_n1128), .B2(new_n1108), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1105), .B2(new_n1096), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1110), .A2(new_n601), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1100), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(KEYINPUT119), .C1(new_n1105), .C2(new_n1104), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1053), .B(new_n1078), .C1(new_n1125), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1071), .A2(new_n1139), .A3(new_n1077), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1051), .A2(G301), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1030), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1002), .A2(KEYINPUT114), .A3(new_n1021), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n1021), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1060), .A2(G8), .A3(G168), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT115), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n990), .A2(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n960), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(new_n992), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n992), .A2(new_n1027), .A3(new_n1149), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(KEYINPUT63), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n992), .A2(new_n1145), .A3(new_n1144), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1021), .A2(new_n1000), .A3(new_n578), .A4(new_n577), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1019), .B1(new_n1156), .B2(new_n1007), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n958), .B1(new_n1143), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n949), .A2(new_n681), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT46), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(KEYINPUT126), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1161), .B(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n948), .B1(new_n781), .B2(new_n951), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(KEYINPUT126), .B2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT47), .Z(new_n1168));
  NOR2_X1   g743(.A1(new_n955), .A2(new_n948), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT127), .Z(new_n1170));
  INV_X1    g745(.A(KEYINPUT48), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1170), .A2(new_n1171), .B1(new_n948), .B2(new_n953), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n951), .A2(new_n952), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n722), .A2(new_n725), .ZN(new_n1176));
  INV_X1    g751(.A(new_n810), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1175), .A2(new_n1176), .B1(G2067), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1168), .B(new_n1174), .C1(new_n949), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1160), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(G319), .ZN(new_n1182));
  OR3_X1    g756(.A1(G401), .A2(new_n1182), .A3(G227), .ZN(new_n1183));
  NOR3_X1   g757(.A1(new_n689), .A2(new_n690), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n939), .A2(new_n1184), .A3(new_n883), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


