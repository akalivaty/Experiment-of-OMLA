//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n227), .B1(new_n202), .B2(new_n228), .C1(new_n203), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n214), .A2(new_n220), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n228), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  INV_X1    g0046(.A(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT65), .ZN(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n248), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n216), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n257), .A3(new_n216), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n207), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n264), .A2(new_n266), .B1(G50), .B2(new_n263), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT69), .B1(new_n202), .B2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(G58), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT8), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(new_n273), .A3(KEYINPUT8), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n215), .A2(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n269), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n267), .B1(new_n279), .B2(new_n259), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT71), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT9), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G222), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G223), .A2(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n289), .B(new_n292), .C1(G77), .C2(new_n285), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n291), .A3(G274), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n293), .B(new_n297), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n282), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n308), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n282), .A2(new_n310), .A3(new_n305), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n301), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(G179), .B2(new_n301), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n280), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n275), .A2(new_n276), .A3(new_n265), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n275), .A2(new_n276), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n264), .A2(new_n319), .B1(new_n320), .B2(new_n263), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(G223), .A2(G1698), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n298), .A2(G1698), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G87), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n292), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n291), .A2(G232), .A3(new_n299), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n297), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(G200), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n291), .B1(new_n327), .B2(new_n328), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n297), .A2(new_n331), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n334), .A2(new_n335), .A3(G190), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT75), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n325), .A2(new_n326), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n215), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n283), .A2(new_n208), .A3(new_n284), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT7), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n344), .A3(G68), .ZN(new_n345));
  AND2_X1   g0145(.A1(G58), .A2(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G58), .A2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n268), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AND4_X1   g0151(.A1(new_n339), .A2(new_n345), .A3(KEYINPUT16), .A4(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n203), .B1(new_n343), .B2(KEYINPUT7), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n353), .B2(new_n342), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n339), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT64), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT7), .B1(new_n285), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n340), .A2(new_n341), .A3(new_n208), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(G68), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n351), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n255), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n322), .B(new_n338), .C1(new_n356), .C2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT17), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n322), .B1(new_n356), .B2(new_n367), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n330), .A2(new_n332), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT76), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n330), .A2(new_n332), .A3(new_n375), .A4(new_n372), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n313), .B1(new_n334), .B2(new_n335), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n351), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n354), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n255), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n364), .B2(new_n365), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n321), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT18), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n379), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n379), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n369), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n228), .A2(G1698), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n229), .A2(new_n286), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n285), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n244), .B2(new_n285), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n291), .B1(new_n396), .B2(KEYINPUT70), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(KEYINPUT70), .B2(new_n396), .ZN(new_n398));
  INV_X1    g0198(.A(new_n300), .ZN(new_n399));
  INV_X1    g0199(.A(G274), .ZN(new_n400));
  AND2_X1   g0200(.A1(G1), .A2(G13), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n290), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n399), .A2(G244), .B1(new_n402), .B2(new_n296), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n372), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT15), .B(G87), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n278), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT8), .B(G58), .ZN(new_n408));
  INV_X1    g0208(.A(new_n268), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n222), .A2(new_n215), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n255), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n261), .A2(new_n208), .A3(G1), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n222), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n384), .A2(new_n265), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n411), .B(new_n413), .C1(new_n222), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n404), .A2(G169), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n203), .A2(G20), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n420), .B1(new_n201), .B2(new_n409), .C1(new_n278), .C2(new_n222), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n421), .A2(new_n259), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(KEYINPUT11), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(KEYINPUT11), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n262), .A2(KEYINPUT12), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n420), .B1(new_n412), .B2(KEYINPUT12), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n414), .A2(KEYINPUT12), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(G68), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n298), .A2(new_n286), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n228), .A2(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n325), .C2(new_n326), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n436), .B2(new_n292), .ZN(new_n437));
  AOI211_X1 g0237(.A(KEYINPUT73), .B(new_n291), .C1(new_n434), .C2(new_n435), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n291), .A2(G238), .A3(new_n299), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT74), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n297), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n297), .B2(new_n439), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n437), .A2(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT13), .ZN(new_n446));
  NOR2_X1   g0246(.A1(G226), .A2(G1698), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n228), .B2(G1698), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(new_n285), .B1(G33), .B2(G97), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT73), .B1(new_n449), .B2(new_n291), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n436), .A2(new_n431), .A3(new_n292), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n443), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n441), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n446), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n430), .B(G169), .C1(new_n445), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n454), .A3(new_n446), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(G179), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n458), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n430), .B1(new_n461), .B2(G169), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n429), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n429), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(G200), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n303), .C2(new_n461), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n404), .A2(G190), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n398), .A2(new_n403), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n415), .B1(new_n468), .B2(G200), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n419), .A2(new_n463), .A3(new_n466), .A4(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n318), .A2(new_n392), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n285), .A2(new_n215), .A3(G87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n285), .A2(new_n215), .A3(new_n475), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n215), .A2(KEYINPUT23), .A3(G107), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G116), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(G20), .B2(new_n244), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT24), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n477), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n255), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n262), .A2(G20), .A3(new_n244), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT25), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n207), .A2(G33), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n256), .A2(new_n263), .A3(new_n258), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(G107), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(G257), .A2(G1698), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n325), .B2(new_n326), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT83), .ZN(new_n497));
  OAI211_X1 g0297(.A(G250), .B(new_n286), .C1(new_n325), .C2(new_n326), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT84), .B(G294), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G33), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT83), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n495), .C1(new_n325), .C2(new_n326), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n497), .A2(new_n498), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n292), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n207), .B(G45), .C1(new_n294), .C2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G41), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(new_n291), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n507), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n295), .A2(G1), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(G41), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n402), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n509), .A2(G190), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT85), .B1(new_n504), .B2(new_n508), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  INV_X1    g0317(.A(new_n508), .ZN(new_n518));
  AOI211_X1 g0318(.A(new_n517), .B(new_n518), .C1(new_n503), .C2(new_n292), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n513), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G200), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n515), .B1(new_n522), .B2(KEYINPUT86), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n494), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G179), .B(new_n513), .C1(new_n516), .C2(new_n519), .ZN(new_n527));
  OAI21_X1  g0327(.A(G169), .B1(new_n509), .B2(new_n514), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n527), .A2(new_n528), .B1(new_n487), .B2(new_n493), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT87), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n494), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n520), .A2(new_n524), .A3(new_n521), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n524), .B1(new_n520), .B2(new_n521), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n534), .A2(new_n535), .A3(new_n515), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n531), .B(new_n533), .C1(new_n536), .C2(new_n494), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G1698), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n540), .B(G244), .C1(new_n326), .C2(new_n325), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n223), .B1(new_n283), .B2(new_n284), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(KEYINPUT4), .ZN(new_n544));
  OAI21_X1  g0344(.A(G250), .B1(new_n325), .B2(new_n326), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n286), .B1(new_n545), .B2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n292), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(new_n291), .C1(new_n505), .C2(new_n507), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n513), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(KEYINPUT78), .B(new_n292), .C1(new_n544), .C2(new_n546), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n263), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G97), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n491), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n361), .A2(G107), .A3(new_n362), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT6), .ZN(new_n560));
  AND2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n244), .A2(KEYINPUT6), .A3(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(new_n360), .B1(G77), .B2(new_n268), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n558), .B1(new_n567), .B2(new_n255), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n547), .A2(G190), .A3(new_n551), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n554), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n229), .A2(new_n286), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n223), .A2(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n325), .C2(new_n326), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n291), .B1(new_n574), .B2(new_n479), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n225), .B1(new_n295), .B2(G1), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n207), .A2(new_n400), .A3(G45), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n291), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n575), .A2(G179), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n357), .A2(new_n359), .A3(G33), .A4(G97), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n224), .A2(new_n557), .A3(new_n244), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n435), .A2(new_n582), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n360), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n285), .A2(new_n215), .A3(G68), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n255), .B1(new_n412), .B2(new_n406), .ZN(new_n589));
  INV_X1    g0389(.A(new_n406), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n492), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n580), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n313), .B1(new_n575), .B2(new_n579), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n255), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n492), .A2(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n406), .A2(new_n412), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n574), .A2(new_n479), .ZN(new_n599));
  OAI211_X1 g0399(.A(G190), .B(new_n578), .C1(new_n599), .C2(new_n291), .ZN(new_n600));
  OAI21_X1  g0400(.A(G200), .B1(new_n575), .B2(new_n579), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n592), .A2(new_n593), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n549), .A2(new_n372), .A3(new_n551), .A4(new_n552), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n567), .A2(new_n255), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT79), .ZN(new_n606));
  INV_X1    g0406(.A(new_n558), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n547), .A2(new_n551), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n313), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n384), .B1(new_n559), .B2(new_n566), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT79), .B1(new_n611), .B2(new_n558), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n604), .A2(new_n608), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n571), .A2(new_n603), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT81), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n286), .A2(G257), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G264), .A2(G1698), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n325), .C2(new_n326), .ZN(new_n618));
  INV_X1    g0418(.A(G303), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n283), .A2(new_n619), .A3(new_n284), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n292), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(G270), .B(new_n291), .C1(new_n505), .C2(new_n507), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n513), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n490), .A2(G116), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n412), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n384), .B1(new_n247), .B2(new_n412), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n254), .A2(new_n216), .B1(G20), .B2(new_n247), .ZN(new_n628));
  INV_X1    g0428(.A(G33), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G97), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n542), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n360), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT20), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n215), .A2(new_n542), .A3(new_n630), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT20), .B1(new_n635), .B2(new_n628), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n627), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n615), .B1(new_n624), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n263), .A2(G116), .A3(new_n490), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n639), .A2(new_n255), .B1(G116), .B2(new_n263), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n633), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(KEYINPUT20), .A3(new_n628), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n623), .A2(G200), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(KEYINPUT81), .A3(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n623), .A2(new_n303), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n638), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n637), .A2(G169), .A3(new_n623), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT80), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n623), .A2(KEYINPUT21), .A3(G169), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n621), .A2(new_n513), .A3(G179), .A4(new_n622), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n654), .B2(new_n637), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n641), .A2(new_n642), .ZN(new_n656));
  AOI221_X4 g0456(.A(KEYINPUT80), .B1(new_n656), .B2(new_n627), .C1(new_n652), .C2(new_n653), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n647), .B(new_n650), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT82), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n637), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT80), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n654), .A2(new_n651), .A3(new_n637), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT82), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n647), .A4(new_n650), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n614), .B1(new_n659), .B2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n472), .A2(new_n538), .A3(new_n666), .ZN(G372));
  NAND2_X1  g0467(.A1(new_n604), .A2(new_n610), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n568), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n575), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n521), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT89), .B1(new_n597), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n672), .B(new_n675), .C1(new_n599), .C2(new_n291), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G200), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n589), .A4(new_n595), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(new_n679), .A3(new_n600), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n313), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n592), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n669), .A2(new_n680), .A3(new_n681), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n592), .A2(new_n593), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n598), .A2(new_n602), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n687), .B2(new_n613), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n684), .A2(new_n688), .A3(new_n683), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n571), .A2(new_n680), .A3(new_n613), .A4(new_n683), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n536), .B2(new_n494), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n650), .A2(new_n660), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n529), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n689), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n472), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n379), .A2(new_n388), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n460), .A2(new_n462), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n702), .A2(new_n429), .B1(new_n418), .B2(new_n466), .ZN(new_n703));
  AOI211_X1 g0503(.A(new_n321), .B(new_n337), .C1(new_n383), .C2(new_n385), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT17), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n701), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n316), .B1(new_n312), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n707), .ZN(G369));
  INV_X1    g0508(.A(new_n494), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n215), .A2(new_n262), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT91), .Z(new_n711));
  INV_X1    g0511(.A(KEYINPUT27), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(G213), .ZN(new_n715));
  INV_X1    g0515(.A(G343), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n538), .B1(new_n709), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n529), .A2(new_n717), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n659), .A2(new_n665), .B1(new_n637), .B2(new_n717), .ZN(new_n722));
  INV_X1    g0522(.A(new_n693), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n718), .A2(new_n723), .A3(new_n643), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n694), .A2(new_n696), .A3(new_n718), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n650), .B1(new_n657), .B2(new_n655), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n530), .A2(new_n537), .A3(new_n730), .A4(new_n718), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n211), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n584), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n218), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n717), .B(new_n614), .C1(new_n659), .C2(new_n665), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n530), .A3(new_n537), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n609), .A2(new_n653), .A3(new_n575), .A4(new_n579), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n516), .A2(new_n519), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT30), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n676), .A2(new_n372), .A3(new_n623), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n520), .A2(new_n553), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n717), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n750), .B2(new_n717), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n741), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G330), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT92), .ZN(new_n756));
  INV_X1    g0556(.A(G330), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n741), .B2(new_n753), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT92), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n763));
  INV_X1    g0563(.A(new_n515), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n525), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n690), .B1(new_n765), .B2(new_n709), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n532), .A2(new_n695), .A3(new_n494), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n695), .B1(new_n532), .B2(new_n494), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n723), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n717), .B1(new_n770), .B2(new_n689), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n680), .A2(new_n683), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n681), .B1(new_n775), .B2(new_n669), .ZN(new_n776));
  INV_X1    g0576(.A(new_n683), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n687), .A2(new_n613), .A3(KEYINPUT26), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n661), .A2(new_n662), .B1(new_n649), .B2(new_n648), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n533), .A2(new_n780), .A3(KEYINPUT94), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT94), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n529), .B2(new_n730), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n766), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(KEYINPUT29), .A3(new_n718), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n774), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n762), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n739), .B1(new_n790), .B2(G1), .ZN(G364));
  NOR2_X1   g0591(.A1(new_n360), .A2(new_n261), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G45), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n734), .A2(new_n794), .A3(new_n207), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n727), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G330), .B2(new_n725), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n208), .B1(KEYINPUT96), .B2(new_n313), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n313), .A2(KEYINPUT96), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n216), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G179), .A2(G200), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n360), .A2(new_n303), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G329), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n521), .A2(G179), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n360), .A2(new_n303), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n215), .A2(new_n372), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G190), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n804), .B1(new_n805), .B2(new_n807), .C1(new_n808), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n303), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G326), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n303), .A2(G200), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G322), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n801), .A2(G190), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n360), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n499), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n806), .A2(G20), .A3(G190), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n285), .B1(new_n824), .B2(G303), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n815), .A2(new_n819), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n813), .A2(G190), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT33), .B(G317), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n812), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n814), .ZN(new_n830));
  INV_X1    g0630(.A(new_n827), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n201), .A2(new_n830), .B1(new_n831), .B2(new_n203), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n340), .B1(new_n824), .B2(G87), .ZN(new_n833));
  INV_X1    g0633(.A(new_n821), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n244), .B2(new_n807), .C1(new_n557), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G159), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n802), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n202), .A2(new_n817), .B1(new_n811), .B2(new_n222), .ZN(new_n840));
  NOR4_X1   g0640(.A1(new_n832), .A2(new_n835), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n800), .B1(new_n829), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n795), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n211), .A2(new_n285), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(KEYINPUT95), .B2(G355), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(KEYINPUT95), .B2(G355), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n252), .A2(new_n295), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n733), .A2(new_n285), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(G45), .B2(new_n218), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n846), .B1(G116), .B2(new_n211), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(G13), .A2(G33), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(G20), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n800), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n843), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n853), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n842), .B(new_n855), .C1(new_n725), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n797), .A2(new_n857), .ZN(G396));
  NOR3_X1   g0658(.A1(new_n416), .A2(new_n417), .A3(new_n717), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n415), .A2(new_n717), .B1(new_n467), .B2(new_n469), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n418), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n772), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n418), .A2(new_n861), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n859), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n698), .A2(new_n865), .A3(new_n718), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n795), .B1(new_n762), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n762), .B2(new_n867), .ZN(new_n869));
  INV_X1    g0669(.A(new_n800), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n818), .A2(G294), .B1(G311), .B2(new_n803), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n224), .B2(new_n807), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n340), .B1(new_n823), .B2(new_n244), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G97), .B2(new_n821), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n874), .B1(new_n247), .B2(new_n811), .C1(new_n830), .C2(new_n619), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n872), .B(new_n875), .C1(G283), .C2(new_n827), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT98), .Z(new_n877));
  INV_X1    g0677(.A(new_n811), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n818), .B1(new_n878), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G150), .ZN(new_n880));
  INV_X1    g0680(.A(G137), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n831), .B2(new_n880), .C1(new_n881), .C2(new_n830), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT34), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n807), .A2(new_n203), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n285), .B1(new_n201), .B2(new_n823), .C1(new_n834), .C2(new_n202), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n886), .B(new_n887), .C1(G132), .C2(new_n803), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n877), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n870), .B1(new_n890), .B2(KEYINPUT99), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(KEYINPUT99), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n800), .A2(new_n851), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n843), .B1(new_n222), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n892), .B(new_n894), .C1(new_n852), .C2(new_n865), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n869), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(G384));
  NOR2_X1   g0697(.A1(new_n792), .A2(new_n207), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n472), .A2(new_n787), .A3(new_n774), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n707), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n345), .A2(new_n351), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n260), .B1(new_n902), .B2(new_n365), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n352), .B2(new_n355), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n715), .B1(new_n904), .B2(new_n322), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n392), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n386), .A2(new_n387), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n713), .A2(new_n714), .A3(G213), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT104), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n370), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT104), .B1(new_n386), .B2(new_n715), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n368), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n259), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n381), .B2(new_n382), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n378), .B1(new_n917), .B2(new_n321), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n368), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n905), .B1(new_n919), .B2(KEYINPUT102), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT102), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n368), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n915), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n914), .B1(new_n923), .B2(KEYINPUT103), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n387), .B1(new_n904), .B2(new_n322), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT102), .B1(new_n704), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n905), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(new_n922), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n906), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(KEYINPUT38), .B(new_n906), .C1(new_n924), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n717), .A2(new_n429), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n463), .A2(new_n466), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT101), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT101), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n463), .A2(new_n466), .A3(new_n939), .A4(new_n936), .ZN(new_n940));
  INV_X1    g0740(.A(new_n936), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n938), .A2(new_n940), .B1(new_n702), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n866), .B2(new_n860), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n935), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n701), .B2(new_n908), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n702), .A2(new_n429), .A3(new_n718), .ZN(new_n946));
  INV_X1    g0746(.A(new_n934), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT103), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n929), .A3(new_n914), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT38), .B1(new_n951), .B2(new_n906), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT39), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n910), .A2(new_n911), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n705), .B2(new_n700), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n912), .A2(new_n368), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n913), .B1(new_n912), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n955), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n913), .ZN(new_n960));
  AND4_X1   g0760(.A1(KEYINPUT106), .A2(new_n912), .A3(new_n368), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n932), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n963));
  NAND3_X1  g0763(.A1(new_n934), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n946), .B1(new_n953), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n945), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n901), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n934), .A2(new_n962), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n938), .A2(new_n940), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n702), .A2(new_n941), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n862), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(KEYINPUT40), .A3(new_n754), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n969), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n973), .A2(KEYINPUT40), .A3(new_n754), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n934), .A2(new_n962), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n754), .B(new_n973), .C1(new_n947), .C2(new_n952), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT40), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n975), .A2(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n981), .A2(new_n472), .A3(new_n754), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n472), .B2(new_n754), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n982), .A2(new_n983), .A3(new_n757), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n898), .B1(new_n968), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n968), .B2(new_n984), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n565), .A2(KEYINPUT35), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n565), .A2(KEYINPUT35), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n987), .A2(G116), .A3(new_n217), .A4(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n218), .A2(new_n346), .A3(new_n222), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n203), .A2(G50), .ZN(new_n993));
  OAI211_X1 g0793(.A(G1), .B(new_n261), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n986), .A2(new_n991), .A3(new_n994), .ZN(G367));
  OAI211_X1 g0795(.A(new_n613), .B(new_n571), .C1(new_n718), .C2(new_n568), .ZN(new_n996));
  INV_X1    g0796(.A(new_n669), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n718), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n731), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT42), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n613), .B1(new_n999), .B2(new_n533), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n718), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n775), .B1(new_n598), .B2(new_n718), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n717), .A2(new_n597), .A3(new_n777), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(KEYINPUT43), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1001), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n728), .A2(new_n999), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n734), .B(KEYINPUT41), .Z(new_n1017));
  OAI211_X1 g0817(.A(new_n719), .B(new_n720), .C1(new_n780), .C2(new_n717), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n1018), .A2(new_n726), .A3(new_n731), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n726), .B1(new_n1018), .B2(new_n731), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n789), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n731), .A2(new_n729), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n999), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n999), .ZN(new_n1026));
  XOR2_X1   g0826(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n728), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n727), .A3(new_n721), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1022), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1017), .B1(new_n1032), .B2(new_n790), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n794), .A2(new_n207), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1016), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n854), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n733), .B2(new_n590), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n848), .A2(new_n241), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n843), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n823), .A2(new_n247), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT46), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n803), .A2(G317), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n817), .A2(new_n619), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n811), .A2(new_n805), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n827), .A2(new_n499), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n807), .A2(new_n557), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n340), .B1(new_n834), .B2(new_n244), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G311), .C2(new_n814), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n807), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(G77), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n285), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n834), .A2(new_n203), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G58), .B2(new_n824), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n880), .B2(new_n817), .ZN(new_n1059));
  INV_X1    g0859(.A(G143), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n830), .B1(new_n831), .B2(new_n836), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n811), .A2(new_n201), .B1(new_n881), .B2(new_n802), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1052), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT47), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1040), .B1(new_n856), .B2(new_n1010), .C1(new_n1065), .C2(new_n870), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1036), .A2(new_n1066), .ZN(G387));
  INV_X1    g0867(.A(new_n1022), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1021), .A2(new_n789), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n734), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1021), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n719), .A2(new_n720), .A3(new_n853), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n844), .A2(new_n736), .B1(G107), .B2(new_n211), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n238), .A2(G45), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n736), .ZN(new_n1075));
  AOI211_X1 g0875(.A(G45), .B(new_n1075), .C1(G68), .C2(G77), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n408), .A2(G50), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n733), .B(new_n285), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1073), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n795), .B1(new_n1080), .B2(new_n1037), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n823), .A2(new_n222), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n803), .B2(G150), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT114), .Z(new_n1084));
  OAI22_X1  g0884(.A1(new_n201), .A2(new_n817), .B1(new_n811), .B2(new_n203), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n834), .A2(new_n406), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n1085), .A2(new_n340), .A3(new_n1048), .A4(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n320), .A2(new_n827), .B1(new_n814), .B2(G159), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n285), .B1(new_n803), .B2(G326), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G303), .A2(new_n878), .B1(new_n818), .B2(G317), .ZN(new_n1091));
  INV_X1    g0891(.A(G322), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1091), .B1(new_n831), .B2(new_n808), .C1(new_n1092), .C2(new_n830), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT48), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n499), .A2(new_n824), .B1(new_n821), .B2(G283), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1090), .B1(new_n247), .B2(new_n807), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1089), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1081), .B1(new_n1103), .B2(new_n800), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1071), .A2(new_n1035), .B1(new_n1072), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1070), .A2(new_n1105), .ZN(G393));
  NAND2_X1  g0906(.A1(new_n1032), .A2(new_n734), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1031), .A2(new_n1029), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1068), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n814), .A2(G317), .B1(new_n818), .B2(G311), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT52), .Z(new_n1111));
  NOR2_X1   g0911(.A1(new_n802), .A2(new_n1092), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n285), .B1(new_n824), .B2(G283), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n244), .B2(new_n807), .C1(new_n247), .C2(new_n834), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G294), .C2(new_n878), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1111), .B(new_n1115), .C1(new_n619), .C2(new_n831), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n814), .A2(G150), .B1(new_n818), .B2(G159), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT51), .Z(new_n1118));
  OAI22_X1  g0918(.A1(new_n811), .A2(new_n408), .B1(new_n1060), .B2(new_n802), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n834), .A2(new_n222), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n807), .A2(new_n224), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n285), .B1(new_n823), .B2(new_n203), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n1123), .C1(new_n201), .C2(new_n831), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n870), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n248), .A2(new_n848), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1037), .B1(G97), .B2(new_n733), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n843), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n856), .C2(new_n998), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1108), .B2(new_n1034), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1109), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G390));
  NAND2_X1  g0936(.A1(new_n758), .A2(new_n973), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT118), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n946), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n943), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n859), .B1(new_n771), .B2(new_n865), .ZN(new_n1141));
  OAI211_X1 g0941(.A(KEYINPUT118), .B(new_n946), .C1(new_n1141), .C2(new_n942), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1140), .A2(new_n953), .A3(new_n964), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT117), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n717), .B(new_n864), .C1(new_n779), .C2(new_n785), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n859), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n786), .A2(new_n718), .ZN(new_n1147));
  OAI211_X1 g0947(.A(KEYINPUT117), .B(new_n860), .C1(new_n1147), .C2(new_n864), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n942), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1139), .B1(new_n934), .B2(new_n962), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1137), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n761), .A2(KEYINPUT119), .A3(new_n865), .A4(new_n1149), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n759), .B1(new_n754), .B2(G330), .ZN(new_n1155));
  AOI211_X1 g0955(.A(KEYINPUT92), .B(new_n757), .C1(new_n741), .C2(new_n753), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n865), .B(new_n1149), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT119), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1143), .A2(new_n1152), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n953), .A2(new_n851), .A3(new_n964), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n893), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n795), .B1(new_n320), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n803), .A2(G294), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n557), .B2(new_n811), .C1(new_n247), .C2(new_n817), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n285), .B(new_n1120), .C1(G87), .C2(new_n824), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n203), .B2(new_n807), .C1(new_n244), .C2(new_n831), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G283), .C2(new_n814), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n814), .A2(G128), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n823), .A2(new_n880), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n340), .B1(new_n821), .B2(G159), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n818), .A2(G132), .B1(G125), .B2(new_n803), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1177), .B1(new_n201), .B2(new_n807), .C1(new_n811), .C2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G137), .C2(new_n827), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1170), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1165), .B1(new_n1181), .B2(new_n800), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1162), .A2(new_n1035), .B1(new_n1163), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1149), .B1(new_n758), .B2(new_n865), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1141), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n865), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT120), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(new_n942), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1149), .B1(new_n761), .B2(new_n865), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1137), .A2(KEYINPUT120), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1189), .B(new_n1192), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1188), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n472), .A2(new_n758), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n899), .A2(new_n707), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1161), .A2(new_n1160), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1153), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1198), .B1(new_n1188), .B2(new_n1195), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n735), .B1(new_n1205), .B2(new_n1162), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1206), .B2(KEYINPUT121), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(new_n735), .C1(new_n1205), .C2(new_n1162), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1183), .B1(new_n1207), .B2(new_n1209), .ZN(G378));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n979), .A2(new_n980), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n970), .A2(new_n969), .A3(new_n974), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT109), .B1(new_n976), .B2(new_n977), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1212), .B(G330), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n312), .B2(new_n317), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n312), .A2(new_n317), .A3(new_n1217), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n281), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1218), .A2(new_n1220), .B1(new_n1221), .B2(new_n715), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1218), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1221), .A2(new_n715), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n1219), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n981), .A2(G330), .A3(new_n1228), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1227), .A2(new_n1229), .A3(new_n966), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n966), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1198), .B1(new_n1162), .B2(new_n1196), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1211), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n967), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1227), .A2(new_n1229), .A3(new_n966), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1190), .A2(new_n942), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1194), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1141), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1192), .A2(new_n1241), .B1(new_n1160), .B2(new_n1185), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1199), .B1(new_n1203), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1243), .A3(KEYINPUT57), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1234), .A2(new_n734), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1226), .A2(new_n851), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n795), .B1(new_n1164), .B2(G50), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n244), .A2(new_n817), .B1(new_n811), .B2(new_n406), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1057), .A2(new_n1082), .A3(G41), .A4(new_n285), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1053), .A2(G58), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n557), .B2(new_n831), .C1(new_n247), .C2(new_n830), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1248), .B(new_n1252), .C1(G283), .C2(new_n803), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(KEYINPUT58), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n818), .A2(G128), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n821), .A2(G150), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1178), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n824), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n827), .A2(G132), .ZN(new_n1260));
  INV_X1    g1060(.A(G125), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n830), .B2(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1259), .B(new_n1262), .C1(G137), .C2(new_n878), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1264), .A2(KEYINPUT59), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(KEYINPUT59), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n629), .B(new_n294), .C1(new_n807), .C2(new_n836), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G124), .B2(new_n803), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1253), .A2(KEYINPUT58), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n201), .B1(new_n325), .B2(G41), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1254), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1247), .B1(new_n1272), .B2(new_n800), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1238), .A2(new_n1035), .B1(new_n1246), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1245), .A2(new_n1274), .ZN(G375));
  AOI22_X1  g1075(.A1(G107), .A2(new_n878), .B1(new_n818), .B2(G283), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n619), .B2(new_n802), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n285), .B(new_n1086), .C1(G97), .C2(new_n824), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n1054), .C1(new_n247), .C2(new_n831), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1277), .B(new_n1279), .C1(G294), .C2(new_n814), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n814), .A2(G132), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT124), .Z(new_n1282));
  NAND2_X1  g1082(.A1(new_n827), .A2(new_n1257), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n821), .A2(G50), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n340), .B1(new_n824), .B2(G159), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1283), .A2(new_n1250), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n878), .A2(G150), .B1(G128), .B2(new_n803), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n881), .B2(new_n817), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1282), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n800), .B1(new_n1280), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n843), .B1(new_n203), .B2(new_n893), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1290), .B(new_n1291), .C1(new_n1149), .C2(new_n852), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1242), .B2(new_n1034), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1188), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT123), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1188), .A2(new_n1195), .A3(KEYINPUT123), .A4(new_n1198), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1017), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1200), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1294), .B1(new_n1299), .B2(new_n1301), .ZN(G381));
  NOR2_X1   g1102(.A1(G375), .A2(G378), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OR4_X1    g1104(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1305));
  OR4_X1    g1105(.A1(G387), .A2(new_n1304), .A3(new_n1305), .A4(G381), .ZN(G407));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(G343), .C2(new_n1304), .ZN(G409));
  NAND4_X1  g1107(.A1(new_n1188), .A2(new_n1195), .A3(KEYINPUT60), .A4(new_n1198), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1308), .A2(new_n734), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1205), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1299), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1294), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n896), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(G384), .A3(new_n1294), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(KEYINPUT126), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n716), .A2(G213), .A3(G2897), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G384), .B1(new_n1312), .B2(new_n1294), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT60), .B1(new_n1242), .B2(new_n1198), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n896), .B(new_n1293), .C1(new_n1323), .C2(new_n1309), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1320), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n716), .A2(G213), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1245), .A2(G378), .A3(new_n1274), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1238), .A2(new_n1243), .A3(new_n1300), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1274), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n734), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1208), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1204), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1333), .A3(new_n1183), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1327), .A2(new_n1334), .ZN(new_n1335));
  AOI22_X1  g1135(.A1(new_n1319), .A2(new_n1325), .B1(new_n1326), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1320), .A3(new_n1318), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT61), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(G396), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(G393), .B(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(G387), .B2(KEYINPUT127), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(G387), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1135), .B1(new_n1342), .B2(new_n1344), .ZN(new_n1345));
  AND2_X1   g1145(.A1(G387), .A2(KEYINPUT127), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G390), .B(new_n1343), .C1(new_n1346), .C2(new_n1341), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1335), .A2(KEYINPUT63), .A3(new_n1326), .A4(new_n1349), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1335), .A2(new_n1326), .A3(new_n1349), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(KEYINPUT125), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT125), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1352), .A2(new_n1356), .A3(new_n1353), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1339), .A2(new_n1351), .A3(new_n1355), .A4(new_n1357), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1321), .A2(new_n1324), .A3(new_n1320), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1325), .B1(new_n1359), .B2(new_n1317), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1335), .A2(new_n1326), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1360), .A2(new_n1338), .A3(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT61), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1352), .A2(KEYINPUT62), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1335), .A2(new_n1365), .A3(new_n1326), .A4(new_n1349), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1362), .A2(new_n1363), .A3(new_n1364), .A4(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1348), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1358), .A2(new_n1369), .ZN(G405));
  NAND3_X1  g1170(.A1(G375), .A2(new_n1333), .A3(new_n1183), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(new_n1327), .ZN(new_n1372));
  XNOR2_X1  g1172(.A(new_n1372), .B(new_n1349), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1373), .B(new_n1368), .ZN(G402));
endmodule


