//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n212), .A2(new_n213), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  INV_X1    g0020(.A(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n228), .B1(new_n206), .B2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n230), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n220), .A2(new_n227), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n202), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n224), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n254), .B2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n257), .B1(new_n261), .B2(new_n202), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n225), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n262), .B1(new_n270), .B2(new_n259), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G222), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(G223), .A3(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G77), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(new_n275), .C1(new_n276), .C2(new_n272), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n281), .A2(new_n284), .A3(G274), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(G226), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n271), .A2(KEYINPUT9), .B1(new_n289), .B2(G200), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n290), .B1(KEYINPUT9), .B2(new_n271), .C1(new_n291), .C2(new_n289), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n268), .A2(G50), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n225), .B2(G68), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n265), .A2(new_n276), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n259), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT11), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  OR3_X1    g0100(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT70), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT70), .B1(new_n299), .B2(new_n300), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n256), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT12), .B1(new_n304), .B2(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(G68), .B2(new_n260), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n301), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n311));
  OR2_X1    g0111(.A1(G226), .A2(G1698), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G33), .ZN(new_n314));
  INV_X1    g0114(.A(G232), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G1698), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n311), .A2(new_n312), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n320), .A2(new_n321), .A3(new_n284), .ZN(new_n322));
  INV_X1    g0122(.A(G238), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n284), .A2(G274), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n286), .B1(new_n324), .B2(new_n280), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT13), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  INV_X1    g0127(.A(new_n325), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n321), .A2(new_n284), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n320), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n330), .A3(G179), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(new_n330), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n333), .A2(new_n332), .A3(new_n335), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n310), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n333), .A2(new_n291), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n310), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n271), .B1(new_n334), .B2(new_n289), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G179), .B2(new_n289), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n285), .B1(G244), .B2(new_n287), .ZN(new_n345));
  NOR2_X1   g0145(.A1(G232), .A2(G1698), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n273), .A2(G238), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n272), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n278), .C1(G107), .C2(new_n272), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G169), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n256), .A2(new_n276), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n261), .B2(new_n276), .ZN(new_n353));
  INV_X1    g0153(.A(new_n263), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n265), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n353), .B1(new_n357), .B2(new_n259), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n350), .A2(G190), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n358), .C1(new_n364), .C2(new_n350), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n344), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n293), .A2(new_n338), .A3(new_n342), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n264), .A2(new_n261), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n256), .B2(new_n264), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n272), .B2(G20), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n313), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT7), .B(new_n225), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT73), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n311), .A2(new_n314), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n225), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n378), .B2(new_n370), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G58), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n303), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n201), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n268), .A2(G159), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n272), .A2(new_n370), .A3(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n377), .B2(new_n225), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n259), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n369), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT74), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(new_n369), .C1(new_n387), .C2(new_n392), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n272), .A2(G226), .A3(G1698), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n272), .A2(G223), .A3(new_n273), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n402), .A2(KEYINPUT76), .A3(new_n278), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT76), .B1(new_n402), .B2(new_n278), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n286), .A2(new_n315), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n406), .A2(new_n285), .A3(G179), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n278), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n406), .A2(new_n285), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n405), .A2(new_n407), .B1(new_n334), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n394), .A2(new_n396), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  AOI21_X1  g0214(.A(G200), .B1(new_n408), .B2(new_n409), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n406), .A2(new_n285), .A3(G190), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n393), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n259), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n371), .A2(new_n374), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n385), .B1(new_n420), .B2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT73), .B1(new_n371), .B2(KEYINPUT7), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n385), .B1(new_n425), .B2(G68), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n422), .B1(new_n426), .B2(KEYINPUT16), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n408), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n402), .A2(KEYINPUT76), .A3(new_n278), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n416), .ZN(new_n431));
  INV_X1    g0231(.A(new_n415), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n427), .A2(new_n433), .A3(KEYINPUT17), .A4(new_n369), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n418), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n394), .A2(new_n436), .A3(new_n396), .A4(new_n411), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n413), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n256), .A2(new_n210), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n419), .B(new_n255), .C1(G1), .C2(new_n282), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n210), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n425), .A2(new_n442), .A3(G107), .ZN(new_n443));
  OAI21_X1  g0243(.A(G107), .B1(new_n375), .B2(new_n379), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  INV_X1    g0245(.A(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT6), .A3(G97), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n210), .A2(new_n446), .ZN(new_n448));
  NOR2_X1   g0248(.A1(G97), .A2(G107), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(KEYINPUT6), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n443), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n441), .B1(new_n453), .B2(new_n259), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G257), .A3(new_n284), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n455), .A2(new_n284), .A3(G274), .A4(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n311), .A2(new_n314), .A3(G244), .A4(new_n273), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n272), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n461), .B1(new_n278), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n364), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(G190), .B2(new_n469), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n454), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n278), .ZN(new_n473));
  INV_X1    g0273(.A(new_n461), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n473), .A2(new_n474), .A3(G179), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n334), .B1(new_n473), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n452), .B1(new_n444), .B2(KEYINPUT77), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n442), .B1(new_n425), .B2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n259), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n441), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n472), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n454), .A2(KEYINPUT78), .A3(new_n471), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n457), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n324), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n457), .A2(new_n209), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n284), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n311), .A2(new_n314), .A3(G238), .A4(new_n273), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n311), .A2(new_n314), .A3(G244), .A4(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT79), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n272), .A2(new_n496), .A3(G244), .A4(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n278), .B1(new_n498), .B2(KEYINPUT80), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n497), .ZN(new_n500));
  INV_X1    g0300(.A(new_n493), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT80), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G190), .B(new_n490), .C1(new_n499), .C2(new_n504), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n440), .A2(new_n208), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n356), .A2(new_n256), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n311), .A2(new_n314), .A3(new_n225), .A4(G68), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n265), .B2(new_n210), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n225), .B1(new_n319), .B2(new_n509), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n449), .A2(new_n208), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT81), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT81), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n506), .B(new_n507), .C1(new_n517), .C2(new_n419), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n490), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n284), .B1(new_n502), .B2(new_n503), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n498), .A2(KEYINPUT80), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n505), .B(new_n519), .C1(new_n523), .C2(new_n364), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n360), .B(new_n490), .C1(new_n499), .C2(new_n504), .ZN(new_n525));
  INV_X1    g0325(.A(new_n516), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n514), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n259), .B1(new_n527), .B2(new_n511), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n507), .C1(new_n356), .C2(new_n440), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n525), .B(new_n529), .C1(new_n523), .C2(G169), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n458), .A2(new_n284), .ZN(new_n532));
  INV_X1    g0332(.A(G270), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n460), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n377), .A2(new_n211), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n273), .B1(G303), .B2(new_n377), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n311), .A2(new_n314), .A3(G264), .A4(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT82), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n272), .A2(new_n539), .A3(G264), .A4(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n534), .B1(new_n542), .B2(new_n278), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G190), .ZN(new_n544));
  INV_X1    g0344(.A(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n256), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n440), .B2(new_n545), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(G33), .B2(G283), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n282), .A2(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n258), .A2(new_n224), .B1(G20), .B2(new_n545), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n550), .A2(new_n551), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT83), .B1(new_n548), .B2(new_n549), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT20), .B(new_n553), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n547), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n284), .B1(new_n536), .B2(new_n541), .ZN(new_n561));
  OAI21_X1  g0361(.A(G200), .B1(new_n561), .B2(new_n534), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n544), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  OAI21_X1  g0364(.A(G169), .B1(new_n561), .B2(new_n534), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n561), .A2(new_n360), .A3(new_n534), .ZN(new_n567));
  INV_X1    g0367(.A(new_n547), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT20), .B1(new_n552), .B2(new_n553), .ZN(new_n569));
  INV_X1    g0369(.A(new_n559), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n542), .A2(new_n278), .ZN(new_n573));
  INV_X1    g0373(.A(new_n534), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(new_n571), .A3(KEYINPUT21), .A4(G169), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n563), .A2(new_n566), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n311), .A2(new_n314), .A3(new_n225), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n272), .A2(new_n580), .A3(new_n225), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT84), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n225), .B2(G107), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT23), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n583), .B(new_n586), .C1(new_n225), .C2(G107), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n585), .A2(new_n587), .B1(G116), .B2(new_n266), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n582), .B2(new_n588), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n259), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT25), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n255), .B2(G107), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n255), .A2(new_n594), .A3(G107), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n440), .A2(new_n446), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n272), .A2(G257), .A3(G1698), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n272), .A2(G250), .A3(new_n273), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G33), .A2(G294), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n278), .B1(new_n457), .B2(new_n455), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n278), .B1(G264), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(G190), .A3(new_n460), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n278), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(G264), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n460), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n593), .A2(new_n599), .A3(new_n606), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n589), .B(KEYINPUT24), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n598), .B1(new_n612), .B2(new_n259), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n334), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n360), .A3(new_n460), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n611), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n531), .A2(new_n577), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NOR4_X1   g0419(.A1(new_n367), .A2(new_n438), .A3(new_n486), .A4(new_n619), .ZN(G372));
  INV_X1    g0420(.A(new_n344), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n293), .B(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n340), .A2(new_n341), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n338), .B1(new_n624), .B2(new_n362), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n435), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n393), .A2(new_n411), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(new_n436), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n621), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n367), .A2(new_n438), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n593), .A2(new_n599), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(new_n614), .A3(new_n615), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n566), .A3(new_n572), .A4(new_n576), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n490), .B1(new_n499), .B2(new_n504), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G200), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n518), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n528), .A2(KEYINPUT85), .A3(new_n507), .A4(new_n506), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n640), .A3(new_n505), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n530), .A3(new_n611), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n486), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n469), .A2(G179), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n644), .B(KEYINPUT86), .C1(new_n334), .C2(new_n469), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT86), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n475), .B2(new_n476), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n454), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n530), .A4(new_n641), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n480), .A2(new_n481), .ZN(new_n652));
  INV_X1    g0452(.A(new_n477), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT26), .B1(new_n531), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n655), .A3(new_n530), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n643), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n630), .A2(new_n658), .ZN(G369));
  NOR2_X1   g0459(.A1(new_n613), .A2(new_n616), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n230), .A2(G1), .A3(G20), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT27), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  INV_X1    g0464(.A(G213), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n661), .B2(new_n662), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G343), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n632), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n660), .B1(new_n671), .B2(new_n611), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n633), .A2(new_n670), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n566), .A2(new_n572), .A3(new_n576), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n668), .B(KEYINPUT89), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n673), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n676), .A2(new_n560), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n577), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n674), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n232), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  NOR4_X1   g0488(.A1(new_n688), .A2(new_n254), .A3(G116), .A4(new_n513), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n223), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  NAND4_X1  g0491(.A1(new_n618), .A2(new_n485), .A3(new_n484), .A4(new_n676), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n543), .A2(G179), .A3(new_n469), .A4(new_n605), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n635), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n605), .A2(new_n473), .A3(new_n474), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n523), .A2(KEYINPUT30), .A3(new_n697), .A4(new_n567), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n469), .A2(G179), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n635), .A2(new_n575), .A3(new_n699), .A4(new_n609), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(new_n670), .ZN(new_n702));
  XNOR2_X1  g0502(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(KEYINPUT31), .B2(new_n702), .ZN(new_n706));
  OAI21_X1  g0506(.A(G330), .B1(new_n693), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n657), .A2(new_n676), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n641), .A2(new_n530), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n652), .A2(new_n647), .A3(new_n645), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT26), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT91), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n530), .B(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n482), .A2(new_n650), .A3(new_n524), .A4(new_n530), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n676), .C1(new_n643), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n708), .B1(new_n711), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n691), .B1(new_n720), .B2(G1), .ZN(G364));
  NOR2_X1   g0521(.A1(new_n230), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n254), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n688), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n232), .A2(G355), .A3(new_n272), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G116), .B2(new_n232), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n272), .B(new_n687), .C1(new_n456), .C2(new_n223), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n252), .A2(G45), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n224), .B1(G20), .B2(new_n334), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n725), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n225), .B1(new_n738), .B2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n225), .A2(new_n291), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n360), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n225), .A2(G190), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI22_X1  g0548(.A1(G322), .A2(new_n745), .B1(new_n748), .B2(G311), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n364), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n377), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n291), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n741), .B(new_n753), .C1(G326), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n754), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n746), .A2(new_n738), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT95), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT95), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n742), .A2(new_n751), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT94), .Z(new_n769));
  AOI22_X1  g0569(.A1(new_n767), .A2(G329), .B1(G303), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n756), .A2(new_n761), .A3(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n744), .A2(new_n381), .B1(new_n747), .B2(new_n276), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT92), .ZN(new_n773));
  INV_X1    g0573(.A(new_n755), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n773), .B1(new_n202), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n773), .B2(new_n772), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT93), .Z(new_n777));
  NAND2_X1  g0577(.A1(new_n763), .A2(G159), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n272), .B1(new_n752), .B2(new_n446), .C1(new_n208), .C2(new_n768), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n739), .A2(new_n210), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n759), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n303), .ZN(new_n784));
  OR3_X1    g0584(.A1(new_n779), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n771), .B1(new_n777), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n737), .B1(new_n786), .B2(new_n734), .ZN(new_n787));
  INV_X1    g0587(.A(new_n733), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n682), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n725), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n683), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n682), .A2(G330), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(G396));
  OAI21_X1  g0593(.A(new_n365), .B1(new_n676), .B2(new_n358), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n362), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n676), .A2(new_n361), .A3(new_n359), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n709), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n797), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n676), .B(new_n799), .C1(new_n643), .C2(new_n656), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n725), .B1(new_n801), .B2(new_n707), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n798), .A2(new_n708), .A3(new_n800), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n734), .A2(new_n731), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n790), .B1(new_n276), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n799), .A2(new_n732), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT98), .B(G143), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n745), .A2(new_n809), .B1(new_n748), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n774), .B2(new_n811), .C1(new_n812), .C2(new_n783), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n752), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G68), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n272), .C1(new_n381), .C2(new_n739), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G50), .B2(new_n769), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n815), .B(new_n819), .C1(new_n820), .C2(new_n766), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n813), .A2(new_n814), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G303), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n782), .B1(new_n774), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n377), .B1(new_n744), .B2(new_n740), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n208), .A2(new_n752), .B1(new_n747), .B2(new_n545), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(new_n769), .C2(G107), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n766), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n825), .B(new_n830), .C1(G283), .C2(new_n759), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n823), .B1(new_n832), .B2(KEYINPUT97), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(KEYINPUT97), .B2(new_n832), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n807), .B(new_n808), .C1(new_n734), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n804), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  NOR2_X1   g0637(.A1(new_n722), .A2(new_n254), .ZN(new_n838));
  INV_X1    g0638(.A(G330), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n704), .B1(new_n701), .B2(new_n670), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n692), .A2(new_n842), .A3(KEYINPUT103), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT103), .B1(new_n692), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n670), .A2(new_n310), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n336), .A2(new_n337), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n342), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT100), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n338), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(KEYINPUT100), .B(new_n310), .C1(new_n336), .C2(new_n337), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n342), .A2(new_n846), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT101), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n853), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT101), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(new_n850), .A3(new_n856), .A4(new_n851), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n848), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n845), .A2(new_n858), .A3(new_n797), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n422), .B1(KEYINPUT16), .B2(new_n421), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n369), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n667), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n438), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n411), .ZN(new_n865));
  INV_X1    g0665(.A(new_n667), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(new_n866), .B1(new_n369), .B2(new_n860), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n393), .A2(new_n417), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n394), .A2(new_n396), .A3(new_n667), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n412), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n871), .ZN(new_n875));
  INV_X1    g0675(.A(new_n628), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n418), .A2(new_n434), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n627), .B1(new_n393), .B2(new_n417), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n872), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n859), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n864), .B2(new_n873), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT102), .B1(new_n874), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n877), .B1(KEYINPUT18), .B2(new_n412), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n862), .B1(new_n890), .B2(new_n437), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n869), .A2(new_n872), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  AOI211_X1 g0697(.A(KEYINPUT104), .B(KEYINPUT40), .C1(new_n859), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT104), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n843), .A2(new_n844), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n854), .A2(new_n857), .ZN(new_n901));
  INV_X1    g0701(.A(new_n848), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n797), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n874), .A2(new_n887), .A3(KEYINPUT102), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n900), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n899), .B1(new_n906), .B2(new_n884), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n886), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT105), .Z(new_n909));
  NOR3_X1   g0709(.A1(new_n845), .A2(new_n438), .A3(new_n367), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n839), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n796), .B(KEYINPUT99), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n902), .A2(new_n901), .B1(new_n800), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n897), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n874), .B2(new_n882), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n852), .A2(new_n676), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n893), .A2(new_n895), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n917), .B(new_n919), .C1(new_n920), .C2(new_n916), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n876), .A2(new_n866), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n711), .A2(new_n631), .A3(new_n719), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n630), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n838), .B1(new_n912), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n912), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(G116), .A3(new_n226), .A4(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n222), .A2(new_n276), .A3(new_n382), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n303), .A2(G50), .ZN(new_n934));
  OAI211_X1 g0734(.A(G1), .B(new_n230), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n928), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NOR2_X1   g0736(.A1(new_n676), .A2(new_n454), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n486), .A2(new_n937), .B1(new_n713), .B2(new_n676), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n678), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n660), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n670), .B1(new_n941), .B2(new_n654), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT43), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n676), .A2(new_n640), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n712), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n530), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n944), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n940), .C2(new_n942), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n684), .A2(new_n938), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n688), .B(KEYINPUT41), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n679), .A2(new_n938), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT107), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT107), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n679), .A2(new_n965), .A3(new_n938), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n679), .A2(new_n938), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n684), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n674), .B(new_n677), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(new_n683), .Z(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n720), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n969), .A2(new_n971), .A3(new_n685), .A4(new_n972), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n962), .B1(new_n979), .B2(new_n720), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n961), .B1(new_n980), .B2(new_n724), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT108), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n961), .B(new_n983), .C1(new_n724), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n950), .A2(new_n733), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n244), .A2(new_n232), .A3(new_n377), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n735), .B1(new_n232), .B2(new_n356), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n725), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n272), .B1(new_n768), .B2(new_n381), .ZN(new_n990));
  INV_X1    g0790(.A(new_n739), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(G68), .B2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n745), .A2(G150), .B1(new_n816), .B2(G77), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n748), .A2(G50), .B1(new_n763), .B2(G137), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n755), .A2(new_n809), .B1(new_n759), .B2(G159), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n769), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n752), .A2(new_n210), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n744), .A2(new_n824), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G317), .C2(new_n763), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n377), .B1(new_n747), .B2(new_n750), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G311), .B2(new_n755), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n991), .A2(G107), .B1(G294), .B2(new_n759), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n768), .A2(new_n545), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(KEYINPUT46), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n996), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n989), .B1(new_n1008), .B2(new_n734), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n986), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n985), .A2(new_n1010), .ZN(G387));
  AOI211_X1 g0811(.A(new_n377), .B(new_n998), .C1(G159), .C2(new_n755), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n739), .A2(new_n356), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n264), .A2(new_n759), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n768), .A2(new_n276), .B1(new_n747), .B2(new_n303), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n744), .A2(new_n202), .B1(new_n762), .B2(new_n812), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n272), .B1(new_n763), .B2(G326), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n768), .A2(new_n740), .B1(new_n739), .B2(new_n750), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G317), .A2(new_n745), .B1(new_n748), .B2(G303), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT110), .B(G322), .Z(new_n1022));
  OAI221_X1 g0822(.A(new_n1021), .B1(new_n774), .B2(new_n1022), .C1(new_n829), .C2(new_n783), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1019), .B1(new_n545), .B2(new_n752), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1018), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n734), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n241), .A2(G45), .A3(new_n377), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n263), .A2(G50), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n456), .B1(new_n303), .B2(new_n276), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n377), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1037), .A2(new_n208), .A3(new_n545), .A4(new_n449), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n687), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n735), .B1(new_n446), .B2(new_n232), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1031), .B(new_n725), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n674), .B2(new_n733), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n976), .B2(new_n724), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n977), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n688), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n976), .A2(new_n720), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  AND3_X1   g0847(.A1(new_n249), .A2(new_n232), .A3(new_n377), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n735), .B1(new_n210), .B2(new_n232), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n725), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(G159), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n774), .A2(new_n812), .B1(new_n744), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n739), .A2(new_n276), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n272), .B1(new_n752), .B2(new_n208), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G50), .C2(new_n759), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n768), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(G68), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n748), .A2(new_n354), .B1(new_n763), .B2(new_n809), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1053), .A2(new_n1056), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n377), .B1(new_n752), .B2(new_n446), .C1(new_n783), .C2(new_n824), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G116), .B2(new_n991), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1022), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n763), .A2(new_n1063), .B1(new_n748), .B2(G294), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(new_n750), .C2(new_n768), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n745), .A2(G311), .B1(G317), .B2(new_n755), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1060), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n734), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n938), .B2(new_n788), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n974), .A2(new_n978), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n723), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n979), .A2(new_n688), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1044), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  OAI211_X1 g0876(.A(new_n676), .B(new_n795), .C1(new_n643), .C2(new_n718), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n796), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT111), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n901), .A2(new_n902), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT111), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1081), .A3(new_n796), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n883), .A2(new_n919), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n882), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n895), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n920), .A2(new_n916), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1087), .A2(new_n1088), .B1(new_n914), .B2(new_n919), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1080), .A2(new_n799), .ZN(new_n1091));
  OAI21_X1  g0891(.A(G330), .B1(new_n843), .B2(new_n844), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n708), .A2(new_n1080), .A3(new_n799), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1085), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n858), .B1(new_n707), .B2(new_n797), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n800), .A2(new_n913), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n858), .B1(new_n1092), .B2(new_n797), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1095), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1092), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n631), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n924), .A2(new_n1107), .A3(new_n630), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1097), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1094), .A2(new_n1109), .A3(new_n1096), .A4(new_n1105), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n688), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT116), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n917), .B1(new_n916), .B2(new_n920), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1100), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n918), .B1(new_n1116), .B2(new_n858), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1115), .A2(new_n1117), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1093), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1096), .B(new_n724), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT112), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT112), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1094), .A2(new_n1122), .A3(new_n724), .A4(new_n1096), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n805), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n725), .B1(new_n264), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n767), .A2(G125), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n744), .A2(new_n820), .B1(new_n752), .B2(new_n202), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n377), .B(new_n1128), .C1(new_n748), .C2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n783), .A2(new_n811), .B1(new_n739), .B2(new_n1051), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G128), .B2(new_n755), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n768), .A2(new_n812), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1127), .A2(new_n1131), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n272), .B1(new_n769), .B2(G87), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT113), .Z(new_n1138));
  AOI21_X1  g0938(.A(new_n1054), .B1(G116), .B2(new_n745), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT114), .Z(new_n1140));
  OAI221_X1 g0940(.A(new_n817), .B1(new_n210), .B2(new_n747), .C1(new_n750), .C2(new_n774), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G107), .B2(new_n759), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n740), .C2(new_n766), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1126), .B1(new_n1144), .B2(new_n734), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT115), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1115), .B2(new_n731), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1114), .B1(new_n1124), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(KEYINPUT116), .B(new_n1148), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1113), .B1(new_n1150), .B2(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n745), .A2(G107), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1153), .A2(KEYINPUT117), .B1(new_n210), .B2(new_n783), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G116), .B2(new_n755), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n767), .A2(G283), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n377), .A2(new_n283), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n768), .A2(new_n276), .B1(new_n747), .B2(new_n356), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(G58), .C2(new_n816), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1153), .A2(KEYINPUT117), .B1(G68), .B2(new_n991), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1155), .A2(new_n1156), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT58), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1157), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT118), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1051), .B2(new_n752), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n783), .A2(new_n820), .B1(new_n747), .B2(new_n811), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT119), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n755), .A2(G125), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n991), .A2(G150), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G128), .A2(new_n745), .B1(new_n1057), .B2(new_n1130), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1168), .B1(new_n1174), .B2(KEYINPUT59), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(KEYINPUT59), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1162), .B2(new_n1161), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n734), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT120), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n790), .B(new_n1179), .C1(new_n202), .C2(new_n805), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n623), .A2(new_n344), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n271), .A2(new_n866), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT55), .Z(new_n1183));
  XNOR2_X1  g0983(.A(new_n1181), .B(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1185));
  XOR2_X1   g0985(.A(new_n1184), .B(new_n1185), .Z(new_n1186));
  OAI21_X1  g0986(.A(new_n1180), .B1(new_n1186), .B2(new_n732), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n839), .B1(new_n859), .B2(new_n885), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n898), .B2(new_n907), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n923), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n923), .B(new_n1189), .C1(new_n898), .C2(new_n907), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1186), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1186), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1188), .B1(new_n1196), .B2(new_n724), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1112), .A2(new_n1109), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1186), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1192), .A2(new_n1193), .A3(new_n1186), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1112), .B2(new_n1109), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n688), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1197), .B1(new_n1199), .B2(new_n1207), .ZN(G375));
  INV_X1    g1008(.A(new_n962), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1101), .A2(new_n1108), .A3(new_n1104), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1110), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1105), .A2(new_n724), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1125), .A2(G68), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1013), .B1(new_n774), .B2(new_n740), .C1(new_n545), .C2(new_n783), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n767), .A2(G303), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n769), .A2(G97), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n272), .B1(new_n816), .B2(G77), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G283), .A2(new_n745), .B1(new_n748), .B2(G107), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n767), .A2(G128), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n769), .A2(G159), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n377), .B1(new_n816), .B2(G58), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G137), .A2(new_n745), .B1(new_n748), .B2(G150), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1130), .A2(new_n759), .B1(G132), .B2(new_n755), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n202), .B2(new_n739), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1214), .A2(new_n1219), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n790), .B(new_n1213), .C1(new_n1227), .C2(new_n734), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1080), .B2(new_n732), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1211), .A2(new_n1212), .A3(new_n1229), .ZN(G381));
  NOR3_X1   g1030(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1075), .A2(new_n1231), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(G387), .A2(G378), .A3(G381), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G375), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT122), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1235), .B(new_n1236), .ZN(G407));
  INV_X1    g1037(.A(new_n1113), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT116), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1124), .A2(new_n1114), .A3(new_n1149), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1238), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n665), .A2(G343), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT123), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G375), .C2(new_n1245), .ZN(G409));
  NAND4_X1  g1046(.A1(new_n1101), .A2(new_n1108), .A3(KEYINPUT60), .A4(new_n1104), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n688), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1110), .A2(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1210), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1212), .A2(new_n1229), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n1250), .A2(new_n836), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n836), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1197), .C1(new_n1199), .C2(new_n1207), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1202), .A2(new_n1209), .A3(new_n1203), .A4(new_n1198), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1202), .A2(new_n724), .A3(new_n1203), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1187), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1242), .A2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1243), .B(new_n1254), .C1(new_n1255), .C2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT126), .B1(new_n1260), .B2(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1243), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1254), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1244), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1254), .A2(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT127), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(KEYINPUT127), .A3(new_n1270), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1261), .A2(new_n1268), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1244), .A2(G2897), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1254), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1252), .A2(G2897), .A3(new_n1243), .A4(new_n1253), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1269), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT61), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(new_n1075), .ZN(new_n1282));
  XOR2_X1   g1082(.A(G393), .B(G396), .Z(new_n1283));
  NAND3_X1  g1083(.A1(new_n985), .A2(G390), .A3(new_n1010), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1283), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G390), .B1(new_n985), .B2(new_n1010), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1010), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1288), .B(new_n1075), .C1(new_n982), .C2(new_n984), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1286), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1281), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1285), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1296));
  XOR2_X1   g1096(.A(new_n1296), .B(KEYINPUT124), .Z(new_n1297));
  AOI21_X1  g1097(.A(new_n1294), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1260), .A2(KEYINPUT63), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(KEYINPUT125), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1300), .A2(KEYINPUT125), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1298), .B(new_n1299), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1292), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1242), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1255), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1264), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1291), .ZN(G402));
endmodule


