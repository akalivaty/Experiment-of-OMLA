//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT65), .B(G77), .Z(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  OAI21_X1  g0024(.A(new_n212), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n206), .A2(new_n213), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n212), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  NAND4_X1  g0036(.A1(new_n227), .A2(new_n228), .A3(new_n233), .A4(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  OAI21_X1  g0053(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT70), .B1(new_n257), .B2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n231), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n256), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n230), .B1(new_n212), .B2(new_n257), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(new_n231), .A3(G1), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n265), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n213), .B1(new_n270), .B2(G20), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n269), .A2(new_n271), .B1(new_n213), .B2(new_n268), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(KEYINPUT72), .A3(new_n272), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(KEYINPUT9), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT73), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n221), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n284), .A2(G223), .B1(new_n285), .B2(new_n282), .ZN(new_n286));
  INV_X1    g0086(.A(G222), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT69), .B(G1698), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n286), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(G1), .A2(G13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n292), .B2(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n295), .A2(new_n301), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(G226), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n296), .A2(G190), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n296), .A2(new_n305), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n275), .A2(new_n276), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT74), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n278), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n278), .B2(new_n312), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n273), .B1(new_n307), .B2(G169), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n307), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G20), .B1(G159), .B2(new_n262), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT76), .B1(new_n257), .B2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n279), .A3(G33), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n326), .A3(new_n281), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n231), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G68), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n327), .B2(new_n231), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT16), .B(new_n323), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT16), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n322), .A2(G20), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n262), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n328), .B1(new_n289), .B2(G20), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n202), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n333), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n332), .A2(new_n340), .A3(new_n265), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n255), .B1(new_n270), .B2(G20), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n269), .B1(new_n268), .B2(new_n255), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT77), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(KEYINPUT77), .A3(new_n343), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n303), .B1(G232), .B2(new_n304), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G87), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n288), .A2(G223), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n327), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n324), .A2(new_n326), .A3(new_n281), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n214), .A2(new_n283), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(KEYINPUT78), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G226), .A2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n327), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n352), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(G179), .B(new_n348), .C1(new_n359), .C2(new_n294), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n295), .A2(new_n301), .ZN(new_n361));
  INV_X1    g0161(.A(G232), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n302), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n358), .ZN(new_n364));
  INV_X1    g0164(.A(new_n352), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n366), .B2(new_n295), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n360), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n346), .A2(new_n347), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n346), .A2(new_n372), .A3(new_n347), .A4(new_n369), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n348), .B1(new_n359), .B2(new_n294), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G200), .ZN(new_n376));
  OAI211_X1 g0176(.A(G190), .B(new_n348), .C1(new_n359), .C2(new_n294), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n341), .A3(new_n343), .A4(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n374), .B1(new_n378), .B2(KEYINPUT80), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n367), .B2(new_n308), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT80), .ZN(new_n382));
  INV_X1    g0182(.A(new_n344), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT17), .A4(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n371), .A2(new_n373), .A3(new_n379), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n268), .ZN(new_n387));
  OR3_X1    g0187(.A1(new_n387), .A2(KEYINPUT12), .A3(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT12), .B1(new_n387), .B2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n202), .B1(new_n270), .B2(G20), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n388), .A2(new_n389), .B1(new_n269), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G77), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n258), .B2(new_n260), .ZN(new_n393));
  INV_X1    g0193(.A(new_n262), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n394), .A2(new_n213), .B1(new_n231), .B2(G68), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n265), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT11), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n280), .A2(new_n281), .A3(G232), .A4(G1698), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n289), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n290), .A2(new_n214), .B1(new_n257), .B2(new_n215), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n295), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n303), .B1(G238), .B2(new_n304), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n257), .A2(new_n215), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT69), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G1698), .ZN(new_n416));
  AND4_X1   g0216(.A1(new_n280), .A2(new_n281), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(G226), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n406), .A2(new_n407), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n294), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G238), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n302), .B1(new_n361), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT13), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n402), .B(G169), .C1(new_n412), .C2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n410), .A2(new_n403), .A3(new_n411), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT13), .B1(new_n420), .B2(new_n422), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(G179), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n402), .B1(new_n429), .B2(G169), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n401), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G200), .B1(new_n412), .B2(new_n423), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n425), .A2(new_n426), .A3(G190), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n400), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n221), .A2(new_n231), .B1(new_n255), .B2(new_n394), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n258), .B2(new_n260), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n265), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n392), .B1(new_n270), .B2(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n269), .A2(new_n440), .B1(new_n221), .B2(new_n268), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n302), .B1(new_n361), .B2(new_n220), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n284), .A2(G238), .B1(G107), .B2(new_n282), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n362), .B2(new_n290), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n444), .B2(new_n295), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n439), .B(new_n441), .C1(new_n445), .C2(new_n308), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(KEYINPUT71), .B1(G190), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(KEYINPUT71), .B2(new_n446), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n445), .A2(new_n319), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(new_n441), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n445), .B2(G169), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n321), .A2(new_n386), .A3(new_n435), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT83), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n300), .A2(G1), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n299), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G264), .A3(new_n294), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n216), .A2(new_n283), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n324), .A2(new_n463), .A3(new_n326), .A4(new_n281), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G294), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n414), .A2(new_n416), .A3(G250), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n257), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n279), .A2(G33), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT87), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n324), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n414), .A2(new_n416), .A3(G250), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT87), .B1(new_n327), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n466), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT88), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n295), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(KEYINPUT88), .B(new_n466), .C1(new_n472), .C2(new_n474), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n462), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n298), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n479), .A2(G190), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(KEYINPUT89), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT89), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n462), .C1(new_n477), .C2(new_n478), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n480), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n486), .B2(new_n308), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n268), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT25), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n257), .A2(G1), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT81), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n269), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n494), .B2(new_n488), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT23), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n231), .B2(G107), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n488), .A2(KEYINPUT23), .A3(G20), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n257), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n497), .A2(new_n498), .B1(new_n500), .B2(new_n231), .ZN(new_n501));
  INV_X1    g0301(.A(G87), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n282), .A2(G20), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(KEYINPUT22), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT22), .A2(G87), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n327), .A2(G20), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g0307(.A(new_n507), .B(KEYINPUT24), .Z(new_n508));
  AOI21_X1  g0308(.A(new_n495), .B1(new_n508), .B2(new_n265), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n487), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G264), .A2(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n414), .A2(new_n416), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n216), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n514), .A2(new_n353), .ZN(new_n515));
  INV_X1    g0315(.A(G303), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n289), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(KEYINPUT86), .B(new_n295), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT86), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n514), .A2(new_n353), .B1(G303), .B2(new_n282), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n294), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n461), .A2(new_n294), .ZN(new_n523));
  INV_X1    g0323(.A(G270), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n480), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n480), .B(KEYINPUT85), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n387), .A2(G116), .ZN(new_n530));
  INV_X1    g0330(.A(new_n494), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n231), .C1(G33), .C2(new_n215), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n534), .B(new_n265), .C1(new_n231), .C2(G116), .ZN(new_n535));
  XOR2_X1   g0335(.A(new_n535), .B(KEYINPUT20), .Z(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n522), .A2(G179), .A3(new_n529), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n368), .B1(new_n532), .B2(new_n536), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n529), .A2(new_n518), .A3(new_n521), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT21), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n500), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n288), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n327), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT84), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G244), .A2(G1698), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n513), .B2(new_n421), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n353), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n545), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n294), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G250), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n459), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n294), .A2(new_n556), .B1(new_n298), .B2(new_n459), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(G200), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n552), .B1(new_n551), .B2(new_n545), .ZN(new_n560));
  AOI211_X1 g0360(.A(KEYINPUT84), .B(new_n500), .C1(new_n550), .C2(new_n353), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n295), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(G190), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n531), .A2(G87), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n215), .B1(new_n258), .B2(new_n260), .ZN(new_n565));
  AOI21_X1  g0365(.A(G20), .B1(new_n413), .B2(KEYINPUT19), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n210), .A2(G87), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n565), .A2(KEYINPUT19), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n327), .A2(G20), .A3(new_n202), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n265), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n437), .A2(new_n268), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n559), .A2(new_n563), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n368), .B1(new_n554), .B2(new_n558), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n562), .A2(new_n319), .A3(new_n557), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n570), .B(new_n571), .C1(new_n494), .C2(new_n437), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n537), .B1(new_n540), .B2(G200), .ZN(new_n580));
  INV_X1    g0380(.A(G190), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n540), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n268), .A2(new_n215), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n494), .B2(new_n215), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n488), .A2(KEYINPUT6), .A3(G97), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n215), .A2(new_n488), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n209), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n587), .B2(KEYINPUT6), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n337), .A2(new_n338), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G107), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n584), .B1(new_n592), .B2(new_n265), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n480), .B1(new_n523), .B2(new_n216), .ZN(new_n595));
  XOR2_X1   g0395(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n596));
  NAND3_X1  g0396(.A1(new_n414), .A2(new_n416), .A3(G244), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n327), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT4), .A4(G244), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n533), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n595), .B1(new_n601), .B2(new_n295), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n308), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(G190), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n602), .A2(G169), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n593), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n319), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n604), .A2(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n544), .A2(new_n579), .A3(new_n582), .A4(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n483), .A2(G179), .A3(new_n480), .A4(new_n485), .ZN(new_n611));
  OAI21_X1  g0411(.A(G169), .B1(new_n479), .B2(new_n481), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n509), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n511), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n455), .A2(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n369), .A2(new_n344), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT18), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n369), .A2(new_n372), .A3(new_n344), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n434), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n431), .B1(new_n621), .B2(new_n453), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n384), .A2(new_n379), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n316), .A2(new_n317), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n320), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n608), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n629), .A2(new_n606), .A3(new_n593), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n574), .A3(new_n578), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT26), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n572), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n564), .A2(new_n570), .A3(KEYINPUT90), .A4(new_n571), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n559), .A3(new_n563), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n630), .A4(new_n578), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n632), .A2(new_n578), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n637), .A2(new_n578), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n609), .B(new_n641), .C1(new_n487), .C2(new_n510), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n542), .A2(new_n543), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n613), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n640), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n628), .B1(new_n455), .B2(new_n646), .ZN(G369));
  NAND2_X1  g0447(.A1(new_n611), .A2(new_n612), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n510), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n270), .A2(new_n231), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n510), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n649), .B(new_n656), .C1(new_n510), .C2(new_n487), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n613), .A2(new_n655), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n655), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n532), .B2(new_n536), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n544), .A2(new_n582), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n486), .A2(new_n308), .ZN(new_n668));
  INV_X1    g0468(.A(new_n482), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n613), .B1(new_n670), .B2(new_n509), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n544), .A2(new_n655), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n613), .B2(new_n660), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  INV_X1    g0475(.A(new_n234), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(G41), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n234), .A2(KEYINPUT91), .A3(new_n299), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n567), .A2(new_n499), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n680), .A2(new_n270), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n229), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n562), .A2(new_n557), .A3(new_n602), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n529), .A2(G179), .A3(new_n518), .A4(new_n521), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n483), .A3(new_n485), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n562), .A2(new_n557), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n602), .A2(G179), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n692), .A2(new_n540), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n486), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(new_n483), .A3(KEYINPUT30), .A4(new_n485), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n698));
  AND3_X1   g0498(.A1(new_n697), .A2(new_n655), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n614), .B2(new_n660), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n691), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n695), .A2(KEYINPUT94), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT94), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n486), .A2(new_n704), .A3(new_n694), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n691), .B2(new_n696), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n655), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n685), .B1(new_n700), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n609), .A2(new_n578), .A3(new_n637), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n670), .B2(new_n509), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n649), .A2(KEYINPUT96), .A3(new_n544), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n613), .B2(new_n643), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n637), .A2(KEYINPUT26), .A3(new_n630), .A4(new_n578), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n578), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n631), .A2(new_n638), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n655), .B1(new_n717), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT97), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n727), .A3(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n645), .A2(new_n660), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n711), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n684), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n664), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n685), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n267), .A2(G20), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G45), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n270), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n680), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n736), .A2(new_n665), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n676), .A2(new_n282), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G355), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G116), .B2(new_n234), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n353), .A2(new_n676), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n300), .B2(new_n229), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n249), .A2(new_n300), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n230), .B1(G20), .B2(new_n368), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n743), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n231), .A2(G179), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  OR3_X1    g0564(.A1(new_n763), .A2(KEYINPUT32), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G87), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT32), .B1(new_n763), .B2(new_n764), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n765), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n761), .A2(new_n581), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n282), .B(new_n770), .C1(G107), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(G20), .A2(G179), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT99), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n581), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT100), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n775), .A2(new_n762), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT101), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n773), .B1(new_n201), .B2(new_n778), .C1(new_n782), .C2(new_n221), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n231), .B1(new_n776), .B2(new_n319), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT102), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT102), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n788), .A2(G97), .B1(new_n790), .B2(G68), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(new_n581), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(new_n213), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n788), .A2(G294), .B1(new_n792), .B2(G326), .ZN(new_n795));
  INV_X1    g0595(.A(new_n790), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT33), .B(G317), .Z(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n763), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n289), .B1(new_n799), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n800), .B1(new_n801), .B2(new_n771), .C1(new_n516), .C2(new_n766), .ZN(new_n802));
  INV_X1    g0602(.A(new_n777), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G322), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n782), .B2(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n783), .A2(new_n794), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n760), .B1(new_n807), .B2(new_n757), .ZN(new_n808));
  INV_X1    g0608(.A(new_n756), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n664), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n745), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  INV_X1    g0612(.A(new_n782), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G116), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G283), .A2(new_n790), .B1(new_n792), .B2(G303), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n282), .B1(new_n766), .B2(new_n488), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n799), .A2(G311), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n502), .B2(new_n771), .C1(new_n777), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G97), .B2(new_n788), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n814), .A2(new_n815), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n327), .B1(new_n799), .B2(G132), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n772), .A2(G68), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n213), .C2(new_n766), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G58), .B2(new_n788), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n792), .B1(new_n790), .B2(G150), .ZN(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n778), .C1(new_n782), .C2(new_n764), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n826), .B1(new_n831), .B2(KEYINPUT104), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT104), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n822), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n757), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n757), .A2(new_n754), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n744), .B1(new_n392), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n450), .A2(new_n655), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n452), .B1(new_n448), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n453), .A2(new_n655), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n836), .B(new_n838), .C1(new_n755), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n730), .B(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n711), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n743), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n737), .A2(new_n270), .ZN(new_n851));
  INV_X1    g0651(.A(new_n628), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n455), .B1(new_n731), .B2(new_n730), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n729), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n400), .A2(new_n660), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n431), .A2(new_n434), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT105), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT105), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n431), .A2(new_n859), .A3(new_n434), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n429), .A2(G169), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT14), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n434), .A2(new_n863), .A3(new_n427), .A4(new_n424), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n855), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT106), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT106), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n867), .A3(new_n855), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n841), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n645), .A2(new_n660), .A3(new_n842), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(new_n333), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n332), .A2(new_n265), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n343), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n653), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n385), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n346), .A2(new_n347), .A3(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n370), .A2(new_n883), .A3(new_n884), .A4(new_n378), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n878), .A2(new_n369), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n886), .A2(new_n880), .A3(new_n378), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n874), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n346), .A2(new_n347), .A3(new_n879), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n617), .A2(new_n378), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n885), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n623), .B2(new_n620), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n890), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n892), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n905));
  INV_X1    g0705(.A(new_n431), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n660), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n620), .A2(new_n653), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n894), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n854), .B(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  INV_X1    g0713(.A(new_n610), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n671), .A2(new_n914), .A3(new_n660), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n708), .A2(new_n915), .A3(new_n698), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n448), .A2(new_n839), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n453), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n872), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n861), .B2(new_n869), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n691), .A2(new_n696), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT93), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(new_n702), .A3(new_n703), .A4(new_n705), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n709), .A3(new_n655), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n916), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n893), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n913), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n913), .B1(new_n901), .B2(new_n892), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n928), .A2(new_n920), .A3(new_n924), .A4(new_n916), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n916), .A2(new_n924), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n455), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n685), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n851), .B1(new_n912), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n912), .B2(new_n934), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n588), .A2(KEYINPUT35), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n588), .A2(KEYINPUT35), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(G116), .A3(new_n232), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n229), .B(new_n285), .C1(new_n201), .C2(new_n202), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(G50), .B2(new_n202), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(G1), .A3(new_n267), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n940), .A3(new_n943), .ZN(G367));
  OAI21_X1  g0744(.A(new_n609), .B1(new_n593), .B2(new_n660), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n630), .A2(new_n655), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n667), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n649), .A2(new_n945), .ZN(new_n951));
  INV_X1    g0751(.A(new_n630), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT107), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n655), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n952), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT107), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n671), .A2(new_n672), .A3(new_n947), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n955), .A2(new_n957), .B1(KEYINPUT42), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(KEYINPUT42), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n641), .B1(new_n636), .B2(new_n660), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n578), .A2(new_n636), .A3(new_n660), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n965), .B1(new_n960), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n950), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n960), .A2(new_n966), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n964), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n949), .A3(new_n967), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n665), .ZN(new_n975));
  INV_X1    g0775(.A(new_n672), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n657), .A2(new_n658), .A3(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n649), .B(new_n672), .C1(new_n510), .C2(new_n487), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT108), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(KEYINPUT108), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT109), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n975), .A2(new_n978), .A3(new_n977), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT109), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n665), .A4(new_n982), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n673), .B2(new_n947), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n613), .A2(new_n660), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n978), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(KEYINPUT44), .A3(new_n948), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n993), .B2(new_n948), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n666), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n999), .A3(new_n667), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n733), .B1(new_n989), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n679), .B(KEYINPUT41), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT110), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n742), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1004), .A2(KEYINPUT110), .A3(new_n1006), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n974), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n758), .B1(new_n234), .B2(new_n437), .C1(new_n750), .C2(new_n245), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n743), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n327), .B1(new_n1014), .B2(new_n763), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n766), .A2(new_n499), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(G97), .C2(new_n772), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n782), .B2(new_n801), .C1(new_n516), .C2(new_n778), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n788), .A2(G107), .B1(new_n790), .B2(G294), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n805), .B2(new_n793), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n221), .A2(new_n771), .ZN(new_n1022));
  INV_X1    g0822(.A(G137), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n289), .B1(new_n763), .B2(new_n1023), .C1(new_n201), .C2(new_n766), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(G150), .C2(new_n803), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n782), .B2(new_n213), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n788), .A2(G68), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n796), .B2(new_n764), .C1(new_n828), .C2(new_n793), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1019), .A2(new_n1021), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT47), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1013), .B1(new_n1030), .B2(new_n757), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n961), .A2(new_n756), .A3(new_n962), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1011), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n813), .A2(G68), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n792), .A2(G159), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT111), .ZN(new_n1039));
  INV_X1    g0839(.A(G150), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n353), .B1(new_n1040), .B2(new_n763), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n285), .A2(new_n767), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n215), .B2(new_n771), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(G50), .C2(new_n803), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n787), .A2(new_n437), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n256), .B2(new_n790), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1037), .A2(new_n1039), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n353), .B1(G326), .B2(new_n799), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n787), .A2(new_n801), .B1(new_n819), .B2(new_n766), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G311), .A2(new_n790), .B1(new_n792), .B2(G322), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n1014), .B2(new_n778), .C1(new_n782), .C2(new_n516), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1048), .B1(new_n499), .B2(new_n771), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1047), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n757), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n659), .A2(new_n756), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n681), .A2(new_n746), .B1(new_n488), .B2(new_n676), .ZN(new_n1061));
  AOI211_X1 g0861(.A(G45), .B(new_n681), .C1(G68), .C2(G77), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT50), .B1(new_n256), .B2(new_n213), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n256), .A2(KEYINPUT50), .A3(new_n213), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n749), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n242), .A2(new_n300), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n744), .B1(new_n1068), .B2(new_n758), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1059), .A2(new_n1060), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n742), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n988), .A2(new_n985), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n987), .B1(new_n981), .B2(new_n982), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n733), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n680), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n733), .A2(new_n1074), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1070), .B1(new_n1071), .B2(new_n989), .C1(new_n1076), .C2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1003), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n995), .A2(new_n999), .A3(new_n667), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n667), .B1(new_n995), .B2(new_n999), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n733), .A2(new_n1074), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n680), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n948), .A2(new_n756), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n757), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n793), .A2(new_n1014), .B1(new_n777), .B2(new_n805), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n767), .A2(G283), .B1(new_n799), .B2(G322), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n282), .B1(new_n488), .B2(new_n771), .C1(new_n1089), .C2(KEYINPUT113), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n813), .B2(G294), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n788), .A2(G116), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n790), .A2(G303), .B1(KEYINPUT113), .B2(new_n1089), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n793), .A2(new_n1040), .B1(new_n777), .B2(new_n764), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n796), .A2(new_n213), .B1(new_n787), .B2(new_n392), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n813), .B2(new_n256), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n327), .B1(new_n799), .B2(G143), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n202), .B2(new_n766), .C1(new_n502), .C2(new_n771), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT112), .Z(new_n1101));
  NAND3_X1  g0901(.A1(new_n1096), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1086), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n252), .A2(new_n749), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n759), .B1(G97), .B2(new_n676), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n744), .B(new_n1103), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT114), .Z(new_n1107));
  AOI22_X1  g0907(.A1(new_n1082), .A2(new_n742), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1084), .A2(new_n1108), .ZN(G390));
  OR3_X1    g0909(.A1(new_n931), .A2(new_n685), .A3(new_n455), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n711), .A2(new_n842), .A3(new_n870), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n916), .A2(new_n924), .A3(G330), .A4(new_n842), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n871), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n841), .B1(new_n724), .B2(new_n918), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n873), .A2(new_n872), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT31), .B1(new_n923), .B2(new_n655), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n697), .A2(new_n655), .A3(new_n698), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n915), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n842), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n871), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n916), .A2(new_n920), .A3(new_n924), .A4(G330), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n854), .B(new_n1110), .C1(new_n1115), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n904), .A2(new_n905), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n874), .B2(new_n908), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n908), .B1(new_n901), .B2(new_n892), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1114), .B2(new_n871), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1128), .A3(new_n1111), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n907), .B1(new_n1116), .B2(new_n871), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n655), .B(new_n840), .C1(new_n717), .C2(new_n723), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n870), .B1(new_n1131), .B2(new_n841), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1130), .A2(new_n1125), .B1(new_n1132), .B2(new_n1127), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n1133), .B2(new_n1122), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n679), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1134), .B2(new_n1124), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n744), .B1(new_n255), .B2(new_n837), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n771), .A2(new_n213), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n282), .B(new_n1138), .C1(G125), .C2(new_n799), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n803), .A2(G132), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT53), .B1(new_n766), .B2(new_n1040), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n766), .A2(KEYINPUT53), .A3(new_n1040), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n788), .A2(G159), .B1(new_n790), .B2(G137), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n793), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1143), .B(new_n1146), .C1(new_n813), .C2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n813), .A2(G97), .B1(G107), .B2(new_n790), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(KEYINPUT115), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n803), .A2(G116), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n289), .B1(new_n799), .B2(G294), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n768), .A3(new_n824), .A4(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n793), .A2(new_n801), .B1(new_n787), .B2(new_n392), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1150), .A2(KEYINPUT115), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1149), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1137), .B1(new_n1158), .B2(new_n1086), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1125), .B2(new_n754), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1134), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n742), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1136), .A2(new_n1162), .ZN(G378));
  XOR2_X1   g0963(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n310), .A2(new_n879), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT55), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n321), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n321), .A2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1165), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n321), .A2(new_n1167), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n321), .A2(new_n1167), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1164), .A3(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n916), .A2(new_n920), .A3(new_n924), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT40), .B1(new_n1175), .B2(new_n893), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n929), .A2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n927), .A2(new_n1179), .A3(G330), .A4(new_n929), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1178), .A2(new_n911), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n911), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1179), .A2(new_n754), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1027), .B1(new_n499), .B2(new_n793), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n327), .A2(new_n299), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1042), .B1(new_n201), .B2(new_n771), .C1(new_n801), .C2(new_n763), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G107), .C2(new_n803), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n437), .B2(new_n782), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1185), .B(new_n1189), .C1(G97), .C2(new_n790), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT58), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT58), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1186), .B(new_n213), .C1(G33), .C2(G41), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n803), .A2(G128), .B1(new_n767), .B2(new_n1148), .ZN(new_n1195));
  INV_X1    g0995(.A(G132), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n796), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n813), .B2(G137), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n788), .A2(G150), .B1(new_n792), .B2(G125), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(KEYINPUT116), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1199), .A2(KEYINPUT116), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n764), .B2(new_n771), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1202), .B2(KEYINPUT59), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1194), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(new_n1086), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n744), .B(new_n1208), .C1(new_n213), .C2(new_n837), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1183), .A2(new_n742), .B1(new_n1184), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n729), .A2(new_n853), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n628), .A3(new_n1110), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1115), .A2(new_n1123), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1134), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1215), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n680), .B(new_n1216), .C1(new_n1217), .C2(KEYINPUT118), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT118), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1219), .B(KEYINPUT57), .C1(new_n1183), .C2(new_n1215), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1210), .B1(new_n1218), .B2(new_n1220), .ZN(G375));
  AOI21_X1  g1021(.A(new_n744), .B1(new_n202), .B2(new_n837), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT121), .Z(new_n1223));
  NOR2_X1   g1023(.A1(new_n777), .A2(new_n801), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n289), .B1(new_n799), .B2(G303), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n392), .B2(new_n771), .C1(new_n215), .C2(new_n766), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(new_n813), .C2(G107), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n793), .A2(new_n819), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1045), .B(new_n1228), .C1(G116), .C2(new_n790), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n793), .A2(new_n1196), .B1(new_n787), .B2(new_n213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n796), .A2(new_n1147), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n353), .B1(new_n1145), .B2(new_n763), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n201), .A2(new_n771), .B1(new_n766), .B2(new_n764), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n778), .A2(new_n1023), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n813), .B2(G150), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1227), .A2(new_n1229), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1223), .B1(new_n1086), .B2(new_n1237), .C1(new_n870), .C2(new_n755), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n742), .B(KEYINPUT119), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1116), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n870), .B1(new_n711), .B2(new_n842), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1122), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1239), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1238), .B1(new_n1245), .B2(KEYINPUT120), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT120), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1247), .B(new_n1239), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT122), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1214), .B2(new_n1239), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT122), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1245), .A2(KEYINPUT120), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1238), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1249), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1214), .A2(new_n1212), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1006), .A3(new_n1124), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(G381));
  NOR3_X1   g1057(.A1(G378), .A2(G396), .A3(G393), .ZN(new_n1258));
  INV_X1    g1058(.A(G384), .ZN(new_n1259));
  INV_X1    g1059(.A(G390), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G387), .A2(new_n1261), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n654), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G407), .B(G213), .C1(G375), .C2(new_n1264), .ZN(G409));
  OAI211_X1 g1065(.A(G378), .B(new_n1210), .C1(new_n1218), .C2(new_n1220), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1183), .A2(new_n1006), .A3(new_n1215), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1209), .A2(new_n1184), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1183), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1239), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1263), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n654), .A2(G213), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1255), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1214), .A2(KEYINPUT60), .A3(new_n1212), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n680), .A3(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1254), .A2(G384), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1254), .B2(new_n1278), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n654), .A2(G213), .A3(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1254), .A2(new_n1278), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1259), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1254), .A2(new_n1278), .A3(G384), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1281), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT124), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1272), .A2(new_n1273), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1291), .A2(KEYINPUT124), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1266), .A2(new_n1271), .B1(G213), .B2(new_n654), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1294), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(G396), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n724), .A2(new_n727), .A3(KEYINPUT29), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n727), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n732), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n846), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1008), .B1(new_n1305), .B2(new_n1005), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1071), .A3(new_n1010), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n970), .A2(new_n973), .ZN(new_n1308));
  AOI221_X4 g1108(.A(new_n1034), .B1(new_n1084), .B2(new_n1108), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1310), .B2(new_n1033), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1300), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1260), .B1(new_n1011), .B2(new_n1034), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(G393), .B(new_n811), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1310), .A2(new_n1033), .A3(G390), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1299), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT123), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1317), .B2(KEYINPUT61), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1312), .A2(new_n1316), .A3(KEYINPUT123), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1290), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n1274), .B2(new_n1288), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1290), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1274), .A2(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1323), .B(new_n1324), .C1(new_n1326), .C2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1318), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1263), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT125), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1290), .A2(new_n1266), .A3(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1290), .B1(new_n1332), .B2(new_n1266), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1331), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1317), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1266), .A2(new_n1332), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1327), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1331), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1290), .A2(new_n1266), .A3(new_n1332), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1335), .A2(new_n1337), .A3(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1312), .A2(new_n1316), .A3(KEYINPUT126), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1344), .B(new_n1347), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1348), .A2(new_n1335), .A3(new_n1337), .A4(new_n1342), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1346), .A2(new_n1349), .ZN(G402));
endmodule


