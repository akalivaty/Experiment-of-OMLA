//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n219), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G351));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n247), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n213), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT11), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT12), .B1(new_n260), .B2(G68), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n262));
  INV_X1    g0062(.A(new_n260), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n255), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n206), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n219), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n261), .A2(new_n262), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n258), .A2(new_n259), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT14), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G226), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G97), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(G232), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(new_n275), .C1(new_n276), .C2(new_n273), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(G238), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n279), .A2(new_n280), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n280), .B1(new_n279), .B2(new_n288), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n271), .B(G169), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n289), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n279), .A2(new_n288), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n289), .A2(new_n290), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n271), .B1(new_n298), .B2(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n270), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(G200), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n292), .B(G190), .C1(new_n293), .C2(new_n294), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n269), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT8), .B(G58), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n266), .ZN(new_n309));
  INV_X1    g0109(.A(G58), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n310), .A2(KEYINPUT8), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(KEYINPUT8), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT73), .B(new_n265), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n264), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(new_n263), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT74), .B1(new_n314), .B2(new_n315), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n272), .B2(G20), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n323));
  OAI211_X1 g0123(.A(KEYINPUT7), .B(new_n207), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT72), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n207), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n319), .ZN(new_n331));
  OAI21_X1  g0131(.A(G68), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n310), .A2(new_n219), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n333), .B2(new_n201), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n247), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT16), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n324), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n329), .B2(new_n207), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT16), .A3(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n255), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n318), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT75), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n318), .C1(new_n338), .C2(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n272), .A2(G226), .A3(G1698), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n272), .A2(G223), .A3(new_n273), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n278), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n286), .A2(G232), .A3(new_n282), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT76), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n286), .A2(new_n355), .A3(G232), .A4(new_n282), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n283), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G169), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n296), .B2(new_n358), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n345), .A2(new_n347), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT17), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n352), .A2(new_n357), .A3(G190), .ZN(new_n365));
  INV_X1    g0165(.A(new_n358), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n364), .B1(new_n344), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n255), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n320), .A2(new_n324), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n336), .B1(new_n371), .B2(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n326), .B1(new_n339), .B2(new_n340), .ZN(new_n374));
  INV_X1    g0174(.A(new_n331), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n336), .B1(new_n376), .B2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n373), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n367), .B1(new_n352), .B2(new_n357), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n366), .B2(G190), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n378), .A2(KEYINPUT17), .A3(new_n380), .A4(new_n318), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n369), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n362), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n345), .A2(new_n347), .A3(new_n360), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n363), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n306), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n272), .A2(G222), .A3(new_n273), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n272), .A2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G223), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n389), .B1(new_n252), .B2(new_n272), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n278), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n283), .B1(G226), .B2(new_n287), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT64), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT64), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G190), .ZN(new_n400));
  INV_X1    g0200(.A(new_n308), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(new_n250), .B1(G150), .B2(new_n247), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(KEYINPUT65), .B1(G20), .B2(new_n203), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(KEYINPUT65), .B2(new_n402), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n255), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n266), .A2(new_n202), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n264), .A2(new_n406), .B1(new_n202), .B2(new_n263), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n396), .A2(G200), .A3(new_n398), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(KEYINPUT9), .A3(new_n407), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n400), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT10), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n401), .A2(new_n247), .B1(G20), .B2(G77), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n250), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n370), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n264), .A2(G77), .A3(new_n265), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(G77), .B2(new_n260), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT67), .ZN(new_n422));
  OR3_X1    g0222(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n419), .B2(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G107), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n390), .A2(new_n220), .B1(new_n426), .B2(new_n272), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n276), .A2(G1698), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n278), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n283), .B1(G244), .B2(new_n287), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n296), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  INV_X1    g0232(.A(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n425), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(G190), .A3(new_n430), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n423), .A2(new_n436), .A3(new_n424), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(KEYINPUT68), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(KEYINPUT68), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n399), .A2(new_n296), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(KEYINPUT66), .B1(new_n405), .B2(new_n407), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT66), .B1(new_n399), .B2(G169), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n414), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT69), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n388), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G303), .B1(new_n322), .B2(new_n323), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n327), .A2(new_n328), .A3(G264), .A4(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n327), .A2(new_n328), .A3(G257), .A4(new_n273), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n278), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT80), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G41), .ZN(new_n462));
  INV_X1    g0262(.A(G41), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT81), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(new_n468), .A3(new_n464), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n206), .B(G45), .C1(new_n463), .C2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n466), .A2(new_n467), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G270), .B(new_n286), .C1(new_n465), .C2(new_n470), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n459), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n206), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n260), .A2(new_n475), .A3(new_n213), .A4(new_n254), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n263), .A2(new_n477), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n254), .A2(new_n213), .B1(G20), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  INV_X1    g0281(.A(G97), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n207), .C1(G33), .C2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n480), .A2(KEYINPUT20), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT20), .B1(new_n480), .B2(new_n483), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n478), .B(new_n479), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(G169), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n474), .A2(KEYINPUT21), .A3(new_n486), .A4(G169), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n469), .A2(new_n467), .A3(new_n471), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n468), .B1(new_n462), .B2(new_n464), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n473), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(new_n486), .A3(G179), .A4(new_n459), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n474), .A2(G200), .ZN(new_n497));
  INV_X1    g0297(.A(new_n486), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G190), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n474), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT86), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n489), .B(new_n496), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n207), .B2(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n426), .A2(KEYINPUT23), .A3(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n249), .A2(new_n477), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n207), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n327), .A2(new_n328), .A3(new_n207), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT22), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT22), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n272), .A2(new_n513), .A3(new_n207), .A4(G87), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n255), .B1(new_n515), .B2(KEYINPUT24), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n517), .B(new_n510), .C1(new_n512), .C2(new_n514), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n476), .A2(new_n426), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT88), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT87), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n522), .B(KEYINPUT25), .C1(new_n260), .C2(G107), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(KEYINPUT25), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT25), .ZN(new_n525));
  AOI21_X1  g0325(.A(G107), .B1(new_n525), .B2(KEYINPUT87), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n263), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n520), .A2(new_n521), .A3(new_n523), .A4(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n523), .C1(new_n426), .C2(new_n476), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT88), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n465), .A2(new_n470), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n278), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n272), .A2(G257), .A3(G1698), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n272), .A2(G250), .A3(new_n273), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G294), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n533), .A2(G264), .B1(new_n537), .B2(new_n278), .ZN(new_n538));
  AOI21_X1  g0338(.A(G200), .B1(new_n538), .B2(new_n472), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n278), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(new_n286), .C1(new_n465), .C2(new_n470), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n472), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n519), .B(new_n531), .C1(new_n539), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n329), .A2(G20), .ZN(new_n545));
  XNOR2_X1  g0345(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n250), .A2(G97), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(G68), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n207), .B1(new_n546), .B2(new_n275), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n221), .A2(new_n482), .A3(new_n426), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n370), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n416), .A2(new_n263), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n416), .B(KEYINPUT85), .Z(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n264), .A3(new_n475), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n206), .A2(new_n281), .A3(G45), .ZN(new_n559));
  INV_X1    g0359(.A(G45), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n222), .B1(new_n560), .B2(G1), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n286), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n327), .A2(new_n328), .A3(G238), .A4(new_n273), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT83), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT83), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n272), .A2(new_n566), .A3(G238), .A4(new_n273), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n327), .A2(new_n328), .A3(G244), .A4(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(new_n508), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n563), .B1(new_n573), .B2(new_n278), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n296), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n571), .B1(new_n567), .B2(new_n565), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n562), .B1(new_n576), .B2(new_n286), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n433), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n558), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n531), .B1(new_n516), .B2(new_n518), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n538), .A2(new_n296), .A3(new_n472), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n542), .A2(new_n433), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n574), .A2(G190), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n476), .A2(new_n221), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n552), .A2(new_n554), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n577), .A2(G200), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n544), .A2(new_n579), .A3(new_n583), .A4(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n503), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n263), .A2(new_n482), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n476), .B2(new_n482), .ZN(new_n592));
  OAI21_X1  g0392(.A(G107), .B1(new_n325), .B2(new_n331), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT78), .ZN(new_n594));
  INV_X1    g0394(.A(new_n247), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n596), .A2(new_n482), .A3(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(G97), .B(G107), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI221_X1 g0399(.A(new_n594), .B1(new_n252), .B2(new_n595), .C1(new_n599), .C2(new_n207), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n596), .ZN(new_n601));
  INV_X1    g0401(.A(new_n597), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n207), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n595), .A2(new_n252), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT78), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n593), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n592), .B1(new_n606), .B2(new_n255), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G257), .B(new_n286), .C1(new_n465), .C2(new_n470), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n491), .B2(new_n492), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n327), .A2(new_n328), .A3(G244), .A4(new_n273), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT4), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n272), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n481), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n278), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT79), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(KEYINPUT79), .A3(new_n278), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n610), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n296), .ZN(new_n622));
  INV_X1    g0422(.A(new_n610), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n617), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n433), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n608), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n616), .A2(KEYINPUT79), .A3(new_n278), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT79), .B1(new_n616), .B2(new_n278), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n610), .B1(new_n278), .B2(new_n616), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G190), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n607), .A3(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n626), .A2(KEYINPUT82), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT82), .B1(new_n626), .B2(new_n633), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n590), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n454), .A2(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n344), .A2(new_n360), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT18), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT18), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n344), .A2(new_n360), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n435), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n301), .B1(new_n642), .B2(new_n304), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n369), .A2(new_n381), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n639), .B(new_n641), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n645), .A2(new_n414), .B1(new_n447), .B2(new_n445), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n588), .A2(KEYINPUT26), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n626), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n588), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n583), .A2(new_n496), .A3(new_n489), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n633), .A3(new_n544), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n651), .B2(new_n626), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n648), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(new_n579), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n646), .B1(new_n454), .B2(new_n654), .ZN(G369));
  NAND2_X1  g0455(.A1(new_n496), .A2(new_n489), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI221_X1 g0464(.A(new_n657), .B1(new_n498), .B2(new_n664), .C1(new_n502), .C2(new_n501), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n656), .A2(new_n486), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n580), .A2(new_n663), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n544), .A2(new_n583), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n583), .B2(new_n664), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n657), .A2(new_n663), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n663), .B(KEYINPUT90), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n583), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT91), .Z(G399));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n550), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n217), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n663), .B1(new_n653), .B2(new_n579), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n680), .B1(new_n653), .B2(new_n579), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n693), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n590), .B(new_n679), .C1(new_n634), .C2(new_n635), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n542), .A2(new_n577), .A3(new_n296), .A4(new_n474), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n621), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n459), .A2(new_n472), .A3(G179), .A4(new_n473), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT92), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n540), .A2(new_n541), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n624), .A2(new_n577), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n494), .A2(new_n703), .A3(G179), .A4(new_n459), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n631), .A2(new_n574), .A3(new_n538), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT30), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n700), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n704), .A2(new_n701), .A3(new_n706), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT30), .B1(new_n710), .B2(new_n711), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n699), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n663), .B1(new_n717), .B2(KEYINPUT93), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  AOI211_X1 g0519(.A(new_n719), .B(new_n699), .C1(new_n715), .C2(new_n716), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n697), .B(new_n714), .C1(new_n721), .C2(KEYINPUT31), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n694), .B(new_n696), .C1(G330), .C2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  XNOR2_X1  g0524(.A(new_n670), .B(KEYINPUT94), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n207), .A2(G13), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n206), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n686), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n725), .B(new_n730), .C1(G330), .C2(new_n667), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT95), .Z(new_n732));
  AOI21_X1  g0532(.A(new_n213), .B1(G20), .B2(new_n433), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n207), .A2(new_n367), .A3(G179), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(new_n500), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G107), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n734), .A2(G190), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n272), .C1(new_n221), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT98), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G20), .A3(new_n500), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT32), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n207), .A2(new_n296), .A3(G190), .A4(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n207), .A2(new_n296), .A3(new_n367), .A4(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n749), .B1(new_n751), .B2(new_n252), .C1(new_n219), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(new_n296), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(new_n367), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n747), .A2(new_n748), .B1(new_n756), .B2(new_n310), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n207), .B1(new_n744), .B2(G190), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n202), .B1(new_n759), .B2(new_n482), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n743), .A2(new_n754), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n756), .ZN(new_n762));
  INV_X1    g0562(.A(new_n758), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G322), .A2(new_n762), .B1(new_n763), .B2(G326), .ZN(new_n764));
  INV_X1    g0564(.A(G294), .ZN(new_n765));
  INV_X1    g0565(.A(G303), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n764), .B1(new_n765), .B2(new_n759), .C1(new_n766), .C2(new_n741), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n738), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  OAI21_X1  g0570(.A(new_n329), .B1(new_n753), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  INV_X1    g0572(.A(G329), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n751), .A2(new_n772), .B1(new_n745), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n767), .A2(new_n769), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n733), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n685), .A2(new_n329), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n777), .A2(G355), .B1(new_n477), .B2(new_n685), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n210), .A2(new_n329), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT96), .Z(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n217), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n245), .A2(new_n560), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n733), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n730), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n786), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n776), .B(new_n788), .C1(new_n667), .C2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n732), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n642), .A2(new_n664), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n425), .A2(new_n663), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n438), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n435), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n695), .A2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n680), .B(new_n797), .C1(new_n653), .C2(new_n579), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n722), .A2(G330), .ZN(new_n801));
  OR3_X1    g0601(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n799), .B2(new_n800), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n802), .A2(new_n730), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n739), .A2(G87), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n772), .B2(new_n745), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT100), .Z(new_n807));
  OAI221_X1 g0607(.A(new_n329), .B1(new_n751), .B2(new_n477), .C1(new_n753), .C2(new_n768), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n741), .A2(new_n426), .B1(new_n482), .B2(new_n759), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n765), .A2(new_n756), .B1(new_n758), .B2(new_n766), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n739), .A2(G68), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n272), .B1(new_n745), .B2(new_n813), .C1(new_n310), .C2(new_n759), .ZN(new_n814));
  INV_X1    g0614(.A(new_n741), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G50), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n752), .A2(G150), .B1(new_n750), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n758), .C1(new_n819), .C2(new_n756), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT34), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n812), .B(new_n816), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n733), .B1(new_n811), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n733), .A2(new_n784), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT99), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n730), .B1(new_n827), .B2(new_n252), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n824), .B(new_n828), .C1(new_n798), .C2(new_n785), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n804), .A2(KEYINPUT102), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT102), .B1(new_n804), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G384));
  XNOR2_X1  g0634(.A(new_n599), .B(KEYINPUT103), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT35), .ZN(new_n836));
  OAI211_X1 g0636(.A(G116), .B(new_n214), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OR3_X1    g0640(.A1(new_n217), .A2(new_n252), .A3(new_n333), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n206), .B(G13), .C1(new_n841), .C2(new_n241), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n269), .A2(new_n664), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n305), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT105), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n300), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n270), .B(KEYINPUT105), .C1(new_n297), .C2(new_n299), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n297), .A2(new_n299), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n844), .B1(new_n850), .B2(new_n305), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n793), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n800), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n373), .B1(KEYINPUT16), .B2(new_n372), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(new_n318), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n661), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n386), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n661), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n345), .A2(new_n347), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n344), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT37), .B1(new_n861), .B2(new_n380), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n361), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n360), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n661), .B1(new_n855), .B2(new_n318), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n344), .A2(new_n368), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  INV_X1    g0670(.A(new_n857), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n644), .B1(new_n361), .B2(new_n362), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n385), .ZN(new_n873));
  INV_X1    g0673(.A(new_n868), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n854), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n639), .A2(new_n641), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n661), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  AOI211_X1 g0679(.A(KEYINPUT106), .B(new_n879), .C1(new_n875), .C2(new_n869), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n869), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(KEYINPUT39), .ZN(new_n883));
  INV_X1    g0683(.A(new_n860), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n877), .B2(new_n644), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n638), .B1(new_n344), .B2(new_n368), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n860), .ZN(new_n889));
  INV_X1    g0689(.A(new_n863), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n870), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n869), .A3(new_n879), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n880), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n663), .B1(new_n847), .B2(new_n848), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n878), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n453), .B1(new_n694), .B2(new_n696), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n646), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(KEYINPUT107), .A2(KEYINPUT31), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n718), .B2(new_n720), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n713), .A2(new_n719), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n717), .A2(KEYINPUT93), .ZN(new_n904));
  INV_X1    g0704(.A(new_n901), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n663), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n697), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n902), .A2(new_n697), .A3(new_n906), .A4(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n892), .A2(new_n869), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n852), .A2(new_n798), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n909), .B2(new_n910), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT40), .B1(new_n875), .B2(new_n869), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n915), .A2(KEYINPUT40), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n453), .A2(new_n911), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n669), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n900), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT109), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n924), .B1(new_n206), .B2(new_n726), .C1(new_n900), .C2(new_n922), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(KEYINPUT109), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n843), .B1(new_n925), .B2(new_n926), .ZN(G367));
  NOR2_X1   g0727(.A1(new_n626), .A2(new_n679), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT110), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n626), .B(new_n633), .C1(new_n607), .C2(new_n679), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n626), .B1(new_n932), .B2(new_n583), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n674), .A3(new_n677), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n933), .A2(new_n679), .B1(KEYINPUT42), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n586), .A2(new_n664), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n579), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n579), .A2(new_n938), .A3(new_n588), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT43), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n935), .A2(new_n943), .A3(new_n942), .A4(new_n936), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n675), .A2(new_n932), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n686), .B(KEYINPUT41), .Z(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT111), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n682), .A2(new_n932), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(KEYINPUT111), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n954), .B(new_n955), .Z(new_n956));
  NAND3_X1  g0756(.A1(new_n678), .A2(new_n681), .A3(new_n931), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT45), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(KEYINPUT112), .A3(new_n676), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n674), .B(new_n677), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n961), .A2(new_n669), .A3(new_n668), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n725), .B2(new_n961), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n676), .A2(KEYINPUT112), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n956), .A2(new_n964), .A3(new_n958), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n960), .A2(new_n723), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n951), .B1(new_n966), .B2(new_n723), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n950), .B1(new_n967), .B2(new_n728), .ZN(new_n968));
  INV_X1    g0768(.A(new_n780), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n787), .B1(new_n210), .B2(new_n416), .C1(new_n969), .C2(new_n236), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n729), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n739), .A2(G77), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n753), .A2(new_n746), .B1(new_n751), .B2(new_n202), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT113), .ZN(new_n974));
  INV_X1    g0774(.A(G150), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n272), .B1(new_n745), .B2(new_n818), .C1(new_n756), .C2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n973), .B2(KEYINPUT113), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n741), .A2(new_n310), .B1(new_n758), .B2(new_n819), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n759), .A2(new_n219), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n972), .A2(new_n974), .A3(new_n977), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n739), .A2(G97), .ZN(new_n982));
  INV_X1    g0782(.A(new_n759), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n762), .A2(G303), .B1(new_n983), .B2(G107), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n772), .C2(new_n758), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n741), .B2(new_n477), .ZN(new_n988));
  INV_X1    g0788(.A(new_n745), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n752), .A2(G294), .B1(new_n989), .B2(G317), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n272), .B1(new_n750), .B2(G283), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n986), .A2(new_n988), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n981), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n971), .B1(new_n994), .B2(new_n733), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n941), .B2(new_n789), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n968), .A2(new_n996), .ZN(G387));
  NAND2_X1  g0797(.A1(new_n963), .A2(new_n723), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(KEYINPUT116), .A3(new_n686), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n723), .B2(new_n963), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT116), .B1(new_n998), .B2(new_n686), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n688), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n777), .A2(new_n1003), .B1(new_n426), .B2(new_n685), .ZN(new_n1004));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n401), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT50), .B1(new_n401), .B2(new_n202), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n688), .B(new_n1005), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n780), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n233), .A2(new_n560), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1004), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n730), .B1(new_n1011), .B2(new_n787), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n674), .B2(new_n789), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n751), .A2(new_n219), .B1(new_n745), .B2(new_n975), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n329), .B(new_n1014), .C1(new_n401), .C2(new_n752), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n741), .A2(new_n252), .B1(new_n758), .B2(new_n746), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G50), .B2(new_n762), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n556), .A2(new_n983), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n982), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n272), .B1(new_n989), .B2(G326), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n815), .A2(G294), .B1(new_n983), .B2(G283), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n752), .A2(G311), .B1(new_n750), .B2(G303), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n763), .A2(G322), .ZN(new_n1023));
  INV_X1    g0823(.A(G317), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(new_n756), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT114), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1021), .B1(new_n1027), .B2(KEYINPUT48), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(KEYINPUT48), .B2(new_n1027), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT49), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1020), .B1(new_n477), .B2(new_n738), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1019), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1013), .B1(new_n1034), .B2(new_n733), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n728), .B2(new_n963), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1002), .A2(new_n1036), .ZN(G393));
  NAND2_X1  g0837(.A1(new_n959), .A2(new_n676), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n956), .A2(new_n675), .A3(new_n958), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(new_n727), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n932), .A2(new_n786), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n787), .B1(new_n482), .B2(new_n210), .C1(new_n969), .C2(new_n240), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n729), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n772), .A2(new_n756), .B1(new_n758), .B2(new_n1024), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n272), .B1(new_n989), .B2(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n751), .B2(new_n765), .C1(new_n766), .C2(new_n753), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n741), .A2(new_n768), .B1(new_n477), .B2(new_n759), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n740), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n753), .A2(new_n202), .B1(new_n751), .B2(new_n308), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n329), .B(new_n1052), .C1(G143), .C2(new_n989), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n815), .A2(G68), .B1(new_n983), .B2(G77), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n805), .A3(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n975), .A2(new_n758), .B1(new_n756), .B2(new_n746), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT51), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n1051), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT117), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n1044), .B1(new_n1059), .B2(new_n733), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1041), .B1(new_n1042), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1040), .A2(new_n998), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n686), .A3(new_n966), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(G390));
  AOI21_X1  g0864(.A(new_n669), .B1(new_n909), .B2(new_n910), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n453), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n898), .A2(new_n646), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n853), .B1(new_n692), .B2(new_n796), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n722), .A2(new_n852), .A3(G330), .A4(new_n798), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n669), .B(new_n797), .C1(new_n909), .C2(new_n910), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1072), .A2(KEYINPUT119), .A3(new_n852), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT119), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n911), .A2(G330), .A3(new_n798), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n852), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1071), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n800), .A2(new_n853), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1065), .A2(new_n914), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1076), .B1(new_n801), .B2(new_n797), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1067), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n895), .ZN(new_n1085));
  AOI221_X4 g0885(.A(new_n870), .B1(new_n863), .B2(new_n867), .C1(new_n386), .C2(new_n857), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT37), .B1(new_n884), .B2(new_n887), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n863), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT38), .B1(new_n1088), .B2(new_n885), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n692), .A2(new_n796), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n793), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1090), .B1(new_n1092), .B2(new_n852), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT38), .B1(new_n858), .B2(new_n868), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n882), .A2(new_n881), .A3(KEYINPUT39), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n854), .A2(new_n1085), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1093), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT118), .B1(new_n1100), .B2(new_n1080), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1069), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1080), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1096), .A2(new_n1097), .B1(new_n854), .B2(new_n1085), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1104), .C1(new_n1105), .C2(new_n1093), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1084), .A2(new_n1101), .A3(new_n1102), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1067), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT119), .B1(new_n1072), .B2(new_n852), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1075), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1070), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1111), .B2(new_n1082), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1093), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n854), .A2(new_n1085), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n894), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1103), .B1(new_n1116), .B2(new_n1104), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1112), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1107), .A2(new_n1118), .A3(new_n686), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1101), .A2(new_n728), .A3(new_n1102), .A4(new_n1106), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n729), .B1(new_n826), .B2(new_n401), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n741), .A2(new_n975), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n202), .B2(new_n738), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n272), .B1(new_n751), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n989), .A2(G125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n753), .B2(new_n818), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n763), .A2(G128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n813), .B2(new_n756), .C1(new_n746), .C2(new_n759), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT120), .Z(new_n1132));
  OAI21_X1  g0932(.A(new_n812), .B1(new_n765), .B2(new_n745), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT121), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n329), .B1(new_n751), .B2(new_n482), .C1(new_n753), .C2(new_n426), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n741), .A2(new_n221), .B1(new_n252), .B2(new_n759), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n477), .A2(new_n756), .B1(new_n758), .B2(new_n768), .ZN(new_n1137));
  OR3_X1    g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1132), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1121), .B1(new_n1139), .B2(new_n733), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n894), .B2(new_n785), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1120), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n1143), .ZN(G378));
  OAI21_X1  g0944(.A(KEYINPUT124), .B1(new_n918), .B2(new_n669), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT124), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n916), .A2(new_n917), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT40), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n916), .B2(new_n912), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1146), .B(G330), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n414), .A2(new_n448), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n408), .A2(new_n859), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1153), .B(new_n1154), .Z(new_n1155));
  NAND3_X1  g0955(.A1(new_n1145), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1157), .B(KEYINPUT124), .C1(new_n669), .C2(new_n918), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n897), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1156), .A2(new_n896), .A3(new_n878), .A4(new_n1158), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n728), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n272), .A2(G41), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G50), .B(new_n1163), .C1(new_n249), .C2(new_n463), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n739), .A2(G58), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n426), .A2(new_n756), .B1(new_n758), .B2(new_n477), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n979), .B(new_n1166), .C1(G77), .C2(new_n815), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1163), .B1(new_n768), .B2(new_n745), .C1(new_n753), .C2(new_n482), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n556), .B2(new_n750), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1164), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n741), .A2(new_n1125), .B1(new_n975), .B2(new_n759), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n762), .A2(G128), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n818), .B2(new_n751), .C1(new_n813), .C2(new_n753), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G125), .C2(new_n763), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT122), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n989), .C2(G124), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n738), .B2(new_n746), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT123), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .C1(new_n1179), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n733), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n730), .B1(new_n202), .B2(new_n825), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1157), .C2(new_n785), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1101), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1108), .B1(new_n1190), .B2(new_n1112), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n1161), .A3(new_n1160), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n687), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(KEYINPUT57), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1076), .A2(new_n784), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n729), .B1(new_n826), .B2(G68), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n753), .A2(new_n477), .B1(new_n766), .B2(new_n745), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n272), .B(new_n1201), .C1(G107), .C2(new_n750), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n768), .A2(new_n756), .B1(new_n758), .B2(new_n765), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G97), .B2(new_n815), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n972), .A3(new_n1018), .A4(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n753), .A2(new_n1125), .B1(new_n751), .B2(new_n975), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n329), .B(new_n1206), .C1(G128), .C2(new_n989), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n762), .A2(G137), .B1(new_n983), .B2(G50), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n815), .A2(G159), .B1(new_n763), .B2(G132), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1207), .A2(new_n1165), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1205), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1200), .B1(new_n1211), .B2(new_n733), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1198), .A2(new_n728), .B1(new_n1199), .B2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1084), .A2(new_n951), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1078), .A2(new_n1067), .A3(new_n1083), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1213), .B1(new_n1214), .B2(new_n1216), .ZN(G381));
  AND3_X1   g1017(.A1(new_n1119), .A2(KEYINPUT125), .A3(new_n1143), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT125), .B1(new_n1119), .B2(new_n1143), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1196), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1002), .A2(new_n791), .A3(new_n1036), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1223), .A2(new_n833), .A3(new_n968), .A4(new_n996), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G381), .A2(new_n1221), .A3(new_n1222), .A4(new_n1224), .ZN(G407));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G343), .C2(new_n1221), .ZN(G409));
  NAND2_X1  g1026(.A1(new_n662), .A2(G213), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1215), .B1(new_n1084), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(KEYINPUT126), .B(new_n1215), .C1(new_n1084), .C2(new_n1228), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n687), .B1(new_n1216), .B2(KEYINPUT60), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(G384), .A3(new_n1213), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G384), .B1(new_n1234), .B2(new_n1213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n687), .B1(new_n1190), .B2(new_n1112), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1142), .B1(new_n1239), .B2(new_n1107), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1240), .B(new_n1189), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1162), .B(new_n1188), .C1(new_n1192), .C2(new_n951), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT125), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G378), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1227), .B(new_n1238), .C1(new_n1241), .C2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT62), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1237), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1227), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G2897), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1235), .A3(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G2897), .B(new_n1250), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1196), .A2(G378), .B1(new_n1220), .B2(new_n1242), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1252), .B(new_n1253), .C1(new_n1254), .C2(new_n1250), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1220), .A2(new_n1242), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n686), .A3(new_n1195), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1189), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(G378), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1227), .A4(new_n1238), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1248), .A2(new_n1255), .A3(new_n1256), .A4(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G390), .A2(new_n968), .A3(new_n996), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G390), .B1(new_n968), .B2(new_n996), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1222), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n791), .B1(new_n1002), .B2(new_n1036), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1267), .A2(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(new_n1223), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1266), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1265), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1277), .B2(new_n1247), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1247), .A2(new_n1277), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1253), .A2(new_n1252), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1262), .A2(new_n1227), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1276), .A2(new_n1283), .ZN(G405));
  NAND2_X1  g1084(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1261), .B1(new_n1196), .B2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1238), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1275), .ZN(G402));
endmodule


