

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n411, n412, n413, n414, n415,
         n416, n417, n418, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n769, n770;

  XNOR2_X1 U372 ( .A(n466), .B(n350), .ZN(n560) );
  INV_X1 U373 ( .A(n423), .ZN(n350) );
  NOR2_X1 U374 ( .A1(n689), .A2(n386), .ZN(n468) );
  NOR2_X1 U375 ( .A1(n592), .A2(n686), .ZN(n594) );
  NOR2_X1 U376 ( .A1(n553), .A2(n691), .ZN(n414) );
  XNOR2_X1 U377 ( .A(n504), .B(n349), .ZN(n553) );
  XNOR2_X1 U378 ( .A(n505), .B(KEYINPUT1), .ZN(n349) );
  XNOR2_X1 U379 ( .A(n469), .B(KEYINPUT70), .ZN(n512) );
  XNOR2_X1 U380 ( .A(n482), .B(G953), .ZN(n497) );
  INV_X1 U381 ( .A(KEYINPUT64), .ZN(n482) );
  INV_X2 U382 ( .A(G125), .ZN(n421) );
  XNOR2_X1 U383 ( .A(n351), .B(n755), .ZN(n409) );
  NAND2_X1 U384 ( .A1(n525), .A2(G221), .ZN(n351) );
  XNOR2_X1 U385 ( .A(n352), .B(KEYINPUT96), .ZN(n589) );
  NOR2_X2 U386 ( .A1(n393), .A2(n691), .ZN(n352) );
  NAND2_X1 U387 ( .A1(n353), .A2(n681), .ZN(n588) );
  INV_X1 U388 ( .A(n574), .ZN(n353) );
  XNOR2_X2 U389 ( .A(n376), .B(n496), .ZN(n574) );
  XNOR2_X2 U390 ( .A(G119), .B(G113), .ZN(n399) );
  XNOR2_X2 U391 ( .A(n399), .B(n398), .ZN(n417) );
  NAND2_X2 U392 ( .A1(n415), .A2(n368), .ZN(n514) );
  XNOR2_X2 U393 ( .A(n370), .B(n400), .ZN(n415) );
  XNOR2_X2 U394 ( .A(n540), .B(n539), .ZN(n568) );
  NAND2_X1 U395 ( .A1(n693), .A2(n694), .ZN(n691) );
  XNOR2_X1 U396 ( .A(n451), .B(n450), .ZN(n595) );
  NOR2_X1 U397 ( .A1(G902), .A2(n646), .ZN(n540) );
  XNOR2_X1 U398 ( .A(n508), .B(n401), .ZN(n400) );
  XNOR2_X1 U399 ( .A(n509), .B(n512), .ZN(n401) );
  XNOR2_X1 U400 ( .A(n512), .B(G146), .ZN(n499) );
  NAND2_X1 U401 ( .A1(n427), .A2(n457), .ZN(n354) );
  NAND2_X1 U402 ( .A1(n427), .A2(n457), .ZN(n405) );
  AND2_X1 U403 ( .A1(n354), .A2(n463), .ZN(n760) );
  XNOR2_X1 U404 ( .A(n378), .B(n505), .ZN(n393) );
  XNOR2_X1 U405 ( .A(n466), .B(n423), .ZN(n355) );
  BUF_X1 U406 ( .A(n570), .Z(n356) );
  XNOR2_X2 U407 ( .A(n412), .B(n591), .ZN(n636) );
  BUF_X1 U408 ( .A(n415), .Z(n357) );
  NAND2_X1 U409 ( .A1(n746), .A2(n371), .ZN(n360) );
  NAND2_X1 U410 ( .A1(n358), .A2(n359), .ZN(n361) );
  NAND2_X1 U411 ( .A1(n360), .A2(n361), .ZN(n370) );
  INV_X1 U412 ( .A(n746), .ZN(n358) );
  INV_X1 U413 ( .A(n371), .ZN(n359) );
  XNOR2_X1 U414 ( .A(G137), .B(G140), .ZN(n502) );
  INV_X1 U415 ( .A(KEYINPUT8), .ZN(n411) );
  XNOR2_X1 U416 ( .A(n440), .B(G478), .ZN(n565) );
  OR2_X1 U417 ( .A1(n732), .A2(G902), .ZN(n440) );
  XNOR2_X1 U418 ( .A(n760), .B(n435), .ZN(n434) );
  NAND2_X1 U419 ( .A1(n383), .A2(n384), .ZN(n507) );
  INV_X1 U420 ( .A(KEYINPUT18), .ZN(n382) );
  XNOR2_X1 U421 ( .A(n569), .B(KEYINPUT104), .ZN(n685) );
  OR2_X1 U422 ( .A1(G237), .A2(G902), .ZN(n513) );
  XNOR2_X1 U423 ( .A(n418), .B(KEYINPUT3), .ZN(n416) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n418) );
  INV_X1 U425 ( .A(KEYINPUT45), .ZN(n442) );
  NAND2_X1 U426 ( .A1(n388), .A2(n458), .ZN(n457) );
  NOR2_X1 U427 ( .A1(n637), .A2(n462), .ZN(n461) );
  XNOR2_X1 U428 ( .A(n486), .B(KEYINPUT25), .ZN(n450) );
  XNOR2_X1 U429 ( .A(n449), .B(G128), .ZN(n448) );
  INV_X1 U430 ( .A(G119), .ZN(n449) );
  XNOR2_X1 U431 ( .A(n502), .B(n447), .ZN(n407) );
  XNOR2_X1 U432 ( .A(KEYINPUT75), .B(KEYINPUT24), .ZN(n447) );
  XNOR2_X1 U433 ( .A(n538), .B(n537), .ZN(n646) );
  XNOR2_X1 U434 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U435 ( .A(n531), .B(n530), .ZN(n538) );
  XNOR2_X1 U436 ( .A(n501), .B(n508), .ZN(n503) );
  XNOR2_X1 U437 ( .A(n499), .B(n498), .ZN(n501) );
  BUF_X1 U438 ( .A(n497), .Z(n762) );
  XNOR2_X1 U439 ( .A(n524), .B(n441), .ZN(n732) );
  XNOR2_X1 U440 ( .A(G116), .B(G122), .ZN(n522) );
  INV_X1 U441 ( .A(KEYINPUT17), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n439), .B(KEYINPUT79), .ZN(n626) );
  NAND2_X1 U443 ( .A1(n624), .A2(n625), .ZN(n439) );
  NOR2_X1 U444 ( .A1(n626), .A2(n367), .ZN(n458) );
  NOR2_X1 U445 ( .A1(G237), .A2(G953), .ZN(n487) );
  XNOR2_X1 U446 ( .A(G113), .B(G131), .ZN(n529) );
  XNOR2_X1 U447 ( .A(G143), .B(G122), .ZN(n533) );
  XOR2_X1 U448 ( .A(G140), .B(G104), .Z(n534) );
  XNOR2_X1 U449 ( .A(n511), .B(n372), .ZN(n371) );
  XNOR2_X1 U450 ( .A(n420), .B(n506), .ZN(n372) );
  XNOR2_X1 U451 ( .A(n507), .B(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U452 ( .A(n748), .B(n500), .ZN(n508) );
  INV_X1 U453 ( .A(KEYINPUT76), .ZN(n500) );
  XNOR2_X1 U454 ( .A(n414), .B(n554), .ZN(n570) );
  INV_X1 U455 ( .A(KEYINPUT92), .ZN(n515) );
  XOR2_X1 U456 ( .A(G137), .B(KEYINPUT5), .Z(n489) );
  INV_X1 U457 ( .A(n637), .ZN(n463) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n748) );
  XNOR2_X1 U459 ( .A(G107), .B(G104), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n404), .B(KEYINPUT95), .ZN(n403) );
  INV_X1 U461 ( .A(G110), .ZN(n404) );
  XNOR2_X1 U462 ( .A(G122), .B(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U463 ( .A(n437), .B(n436), .ZN(n523) );
  XNOR2_X1 U464 ( .A(G107), .B(KEYINPUT7), .ZN(n436) );
  XNOR2_X1 U465 ( .A(n438), .B(KEYINPUT101), .ZN(n437) );
  XNOR2_X1 U466 ( .A(KEYINPUT102), .B(KEYINPUT9), .ZN(n438) );
  INV_X1 U467 ( .A(KEYINPUT89), .ZN(n638) );
  INV_X1 U468 ( .A(KEYINPUT30), .ZN(n429) );
  INV_X1 U469 ( .A(KEYINPUT6), .ZN(n380) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n448), .B(n484), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U473 ( .A(n631), .B(n426), .ZN(n635) );
  XNOR2_X1 U474 ( .A(n632), .B(KEYINPUT108), .ZN(n426) );
  XNOR2_X1 U475 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n455) );
  INV_X1 U476 ( .A(KEYINPUT35), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n733), .B(n734), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n730), .B(n731), .ZN(n424) );
  INV_X1 U479 ( .A(KEYINPUT56), .ZN(n473) );
  AND2_X1 U480 ( .A1(G210), .A2(n513), .ZN(n362) );
  XOR2_X1 U481 ( .A(G131), .B(KEYINPUT4), .Z(n363) );
  NOR2_X1 U482 ( .A1(n614), .A2(n548), .ZN(n364) );
  INV_X1 U483 ( .A(n555), .ZN(n614) );
  XOR2_X1 U484 ( .A(KEYINPUT65), .B(KEYINPUT46), .Z(n365) );
  NAND2_X1 U485 ( .A1(n547), .A2(n470), .ZN(n658) );
  XOR2_X1 U486 ( .A(n546), .B(KEYINPUT22), .Z(n366) );
  XNOR2_X1 U487 ( .A(KEYINPUT71), .B(KEYINPUT48), .ZN(n367) );
  XNOR2_X1 U488 ( .A(G902), .B(KEYINPUT15), .ZN(n368) );
  NOR2_X1 U489 ( .A1(n762), .A2(G952), .ZN(n739) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n369) );
  INV_X1 U491 ( .A(KEYINPUT2), .ZN(n462) );
  XNOR2_X2 U492 ( .A(n510), .B(n479), .ZN(n746) );
  XNOR2_X2 U493 ( .A(n417), .B(n416), .ZN(n510) );
  AND2_X1 U494 ( .A1(n623), .A2(n675), .ZN(n388) );
  NAND2_X1 U495 ( .A1(n636), .A2(n669), .ZN(n456) );
  BUF_X1 U496 ( .A(n770), .Z(n373) );
  BUF_X1 U497 ( .A(n589), .Z(n374) );
  BUF_X1 U498 ( .A(n737), .Z(n375) );
  XNOR2_X1 U499 ( .A(n456), .B(KEYINPUT40), .ZN(n770) );
  NOR2_X1 U500 ( .A1(n642), .A2(G902), .ZN(n376) );
  BUF_X1 U501 ( .A(n609), .Z(n377) );
  XNOR2_X1 U502 ( .A(n396), .B(n366), .ZN(n446) );
  NOR2_X1 U503 ( .A1(n726), .A2(G902), .ZN(n378) );
  NOR2_X1 U504 ( .A1(n726), .A2(G902), .ZN(n504) );
  XNOR2_X1 U505 ( .A(n430), .B(n587), .ZN(n379) );
  XNOR2_X1 U506 ( .A(n430), .B(n587), .ZN(n682) );
  XNOR2_X1 U507 ( .A(n574), .B(n380), .ZN(n555) );
  NAND2_X1 U508 ( .A1(KEYINPUT17), .A2(n382), .ZN(n383) );
  NAND2_X1 U509 ( .A1(n381), .A2(KEYINPUT18), .ZN(n384) );
  BUF_X1 U510 ( .A(n618), .Z(n385) );
  INV_X1 U511 ( .A(n576), .ZN(n386) );
  XNOR2_X2 U512 ( .A(n476), .B(n641), .ZN(n387) );
  NAND2_X2 U513 ( .A1(n478), .A2(n477), .ZN(n476) );
  XNOR2_X1 U514 ( .A(n620), .B(KEYINPUT91), .ZN(n621) );
  NAND2_X1 U515 ( .A1(n633), .A2(n681), .ZN(n472) );
  INV_X2 U516 ( .A(n595), .ZN(n694) );
  XNOR2_X1 U517 ( .A(n409), .B(n406), .ZN(n737) );
  OR2_X2 U518 ( .A1(n737), .A2(G902), .ZN(n451) );
  INV_X1 U519 ( .A(n658), .ZN(n550) );
  XNOR2_X1 U520 ( .A(n685), .B(KEYINPUT87), .ZN(n624) );
  NOR2_X2 U521 ( .A1(n613), .A2(n612), .ZN(n623) );
  BUF_X1 U522 ( .A(n769), .Z(n389) );
  BUF_X1 U523 ( .A(n553), .Z(n390) );
  BUF_X1 U524 ( .A(n355), .Z(n391) );
  INV_X1 U525 ( .A(n433), .ZN(n392) );
  BUF_X1 U526 ( .A(n689), .Z(n394) );
  XNOR2_X1 U527 ( .A(n443), .B(n442), .ZN(n743) );
  XNOR2_X1 U528 ( .A(n588), .B(n429), .ZN(n428) );
  XNOR2_X1 U529 ( .A(n454), .B(n365), .ZN(n613) );
  NOR2_X1 U530 ( .A1(n743), .A2(n640), .ZN(n716) );
  XNOR2_X1 U531 ( .A(n395), .B(n493), .ZN(n494) );
  XNOR2_X2 U532 ( .A(n395), .B(n502), .ZN(n754) );
  XNOR2_X2 U533 ( .A(n413), .B(n363), .ZN(n395) );
  NOR2_X2 U534 ( .A1(n572), .A2(n545), .ZN(n396) );
  XNOR2_X2 U535 ( .A(n397), .B(n521), .ZN(n572) );
  NOR2_X2 U536 ( .A1(n609), .A2(n520), .ZN(n397) );
  XNOR2_X2 U537 ( .A(G116), .B(KEYINPUT73), .ZN(n398) );
  NAND2_X1 U538 ( .A1(n405), .A2(n461), .ZN(n639) );
  XNOR2_X2 U539 ( .A(n483), .B(n411), .ZN(n525) );
  NAND2_X1 U540 ( .A1(n602), .A2(n590), .ZN(n412) );
  AND2_X2 U541 ( .A1(n428), .A2(n589), .ZN(n602) );
  XNOR2_X1 U542 ( .A(n413), .B(n526), .ZN(n441) );
  XNOR2_X2 U543 ( .A(n511), .B(G134), .ZN(n413) );
  XNOR2_X1 U544 ( .A(n357), .B(n723), .ZN(n724) );
  NOR2_X1 U545 ( .A1(n600), .A2(n393), .ZN(n608) );
  XNOR2_X2 U546 ( .A(n421), .B(G146), .ZN(n506) );
  XNOR2_X2 U547 ( .A(n514), .B(n362), .ZN(n633) );
  NOR2_X1 U548 ( .A1(n716), .A2(n368), .ZN(n478) );
  NAND2_X1 U549 ( .A1(n445), .A2(n422), .ZN(n444) );
  NAND2_X1 U550 ( .A1(n560), .A2(n561), .ZN(n422) );
  NAND2_X1 U551 ( .A1(n729), .A2(G210), .ZN(n725) );
  XNOR2_X2 U552 ( .A(n476), .B(n641), .ZN(n729) );
  NAND2_X1 U553 ( .A1(n559), .A2(n355), .ZN(n445) );
  NOR2_X1 U554 ( .A1(n424), .A2(n739), .ZN(G54) );
  NOR2_X1 U555 ( .A1(n425), .A2(n739), .ZN(G63) );
  NAND2_X1 U556 ( .A1(n475), .A2(n645), .ZN(n474) );
  XNOR2_X1 U557 ( .A(n725), .B(n724), .ZN(n475) );
  NOR2_X2 U558 ( .A1(n666), .A2(n616), .ZN(n628) );
  XOR2_X2 U559 ( .A(KEYINPUT10), .B(n506), .Z(n755) );
  XNOR2_X1 U560 ( .A(n465), .B(n649), .ZN(n464) );
  NAND2_X1 U561 ( .A1(n464), .A2(n645), .ZN(n432) );
  NAND2_X1 U562 ( .A1(n444), .A2(n582), .ZN(n443) );
  XNOR2_X1 U563 ( .A(n644), .B(n643), .ZN(n453) );
  NAND2_X1 U564 ( .A1(n453), .A2(n645), .ZN(n452) );
  AND2_X2 U565 ( .A1(n460), .A2(n459), .ZN(n427) );
  XNOR2_X1 U566 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X2 U567 ( .A(n754), .B(n503), .ZN(n726) );
  BUF_X2 U568 ( .A(n633), .Z(n430) );
  NAND2_X1 U569 ( .A1(n431), .A2(n462), .ZN(n477) );
  NAND2_X1 U570 ( .A1(n433), .A2(n434), .ZN(n431) );
  XNOR2_X1 U571 ( .A(n432), .B(n369), .ZN(G60) );
  INV_X1 U572 ( .A(n743), .ZN(n433) );
  INV_X1 U573 ( .A(KEYINPUT83), .ZN(n435) );
  XNOR2_X2 U574 ( .A(n618), .B(KEYINPUT19), .ZN(n609) );
  XNOR2_X2 U575 ( .A(n472), .B(n515), .ZN(n618) );
  AND2_X2 U576 ( .A1(n446), .A2(n364), .ZN(n549) );
  AND2_X1 U577 ( .A1(n446), .A2(n390), .ZN(n547) );
  AND2_X1 U578 ( .A1(n446), .A2(n555), .ZN(n562) );
  XNOR2_X1 U579 ( .A(n452), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U580 ( .A(n474), .B(n473), .ZN(G51) );
  NAND2_X1 U581 ( .A1(n770), .A2(n767), .ZN(n454) );
  XNOR2_X2 U582 ( .A(n601), .B(n455), .ZN(n767) );
  NAND2_X1 U583 ( .A1(n626), .A2(n367), .ZN(n459) );
  NAND2_X1 U584 ( .A1(n627), .A2(n367), .ZN(n460) );
  NAND2_X1 U585 ( .A1(n387), .A2(G475), .ZN(n465) );
  NAND2_X1 U586 ( .A1(n467), .A2(n558), .ZN(n466) );
  XNOR2_X1 U587 ( .A(n468), .B(KEYINPUT34), .ZN(n467) );
  XNOR2_X2 U588 ( .A(KEYINPUT69), .B(G101), .ZN(n469) );
  NOR2_X1 U589 ( .A1(n694), .A2(n700), .ZN(n470) );
  XNOR2_X2 U590 ( .A(n549), .B(KEYINPUT32), .ZN(n769) );
  NOR2_X2 U591 ( .A1(n769), .A2(n550), .ZN(n552) );
  XOR2_X1 U592 ( .A(KEYINPUT86), .B(n607), .Z(n480) );
  NAND2_X1 U593 ( .A1(n603), .A2(n602), .ZN(n481) );
  INV_X1 U594 ( .A(KEYINPUT100), .ZN(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U597 ( .A(n739), .ZN(n645) );
  NAND2_X1 U598 ( .A1(n497), .A2(G234), .ZN(n483) );
  XNOR2_X1 U599 ( .A(G110), .B(KEYINPUT23), .ZN(n484) );
  NAND2_X1 U600 ( .A1(G234), .A2(n368), .ZN(n485) );
  XNOR2_X1 U601 ( .A(KEYINPUT20), .B(n485), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G217), .A2(n542), .ZN(n486) );
  XNOR2_X1 U603 ( .A(G472), .B(KEYINPUT98), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n487), .B(KEYINPUT84), .ZN(n532) );
  NAND2_X1 U605 ( .A1(G210), .A2(n532), .ZN(n488) );
  XNOR2_X1 U606 ( .A(n489), .B(n488), .ZN(n491) );
  INV_X1 U607 ( .A(n499), .ZN(n490) );
  XOR2_X1 U608 ( .A(n491), .B(n490), .Z(n495) );
  BUF_X1 U609 ( .A(n510), .Z(n493) );
  XNOR2_X2 U610 ( .A(G128), .B(KEYINPUT85), .ZN(n492) );
  XNOR2_X2 U611 ( .A(n492), .B(G143), .ZN(n511) );
  XNOR2_X1 U612 ( .A(n494), .B(n495), .ZN(n642) );
  XNOR2_X1 U613 ( .A(KEYINPUT72), .B(G469), .ZN(n505) );
  AND2_X1 U614 ( .A1(G227), .A2(n762), .ZN(n498) );
  INV_X1 U615 ( .A(n390), .ZN(n630) );
  NAND2_X1 U616 ( .A1(G214), .A2(n513), .ZN(n681) );
  NAND2_X1 U617 ( .A1(G224), .A2(n762), .ZN(n509) );
  NAND2_X1 U618 ( .A1(G234), .A2(G237), .ZN(n516) );
  XNOR2_X1 U619 ( .A(n516), .B(KEYINPUT14), .ZN(n517) );
  XNOR2_X1 U620 ( .A(KEYINPUT80), .B(n517), .ZN(n518) );
  NAND2_X1 U621 ( .A1(G952), .A2(n518), .ZN(n711) );
  NOR2_X1 U622 ( .A1(G953), .A2(n711), .ZN(n586) );
  INV_X1 U623 ( .A(G898), .ZN(n742) );
  NAND2_X1 U624 ( .A1(G953), .A2(n742), .ZN(n750) );
  NAND2_X1 U625 ( .A1(G902), .A2(n518), .ZN(n583) );
  NOR2_X1 U626 ( .A1(n750), .A2(n583), .ZN(n519) );
  NOR2_X1 U627 ( .A1(n586), .A2(n519), .ZN(n520) );
  XNOR2_X1 U628 ( .A(KEYINPUT93), .B(KEYINPUT0), .ZN(n521) );
  XNOR2_X1 U629 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U630 ( .A1(G217), .A2(n525), .ZN(n526) );
  XNOR2_X1 U631 ( .A(n755), .B(n527), .ZN(n531) );
  AND2_X1 U632 ( .A1(G214), .A2(n532), .ZN(n536) );
  XNOR2_X1 U633 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(G475), .ZN(n539) );
  NOR2_X1 U635 ( .A1(n565), .A2(n568), .ZN(n541) );
  INV_X1 U636 ( .A(n541), .ZN(n592) );
  NAND2_X1 U637 ( .A1(n542), .A2(G221), .ZN(n543) );
  XOR2_X1 U638 ( .A(KEYINPUT21), .B(n543), .Z(n693) );
  NAND2_X1 U639 ( .A1(n541), .A2(n693), .ZN(n544) );
  XOR2_X1 U640 ( .A(KEYINPUT105), .B(n544), .Z(n545) );
  INV_X1 U641 ( .A(KEYINPUT78), .ZN(n546) );
  INV_X1 U642 ( .A(n694), .ZN(n564) );
  NAND2_X1 U643 ( .A1(n564), .A2(n630), .ZN(n548) );
  INV_X1 U644 ( .A(KEYINPUT44), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n561), .A2(KEYINPUT90), .ZN(n551) );
  XNOR2_X1 U646 ( .A(n552), .B(n551), .ZN(n559) );
  NAND2_X1 U647 ( .A1(n565), .A2(n568), .ZN(n604) );
  INV_X1 U648 ( .A(n604), .ZN(n558) );
  INV_X1 U649 ( .A(KEYINPUT82), .ZN(n554) );
  XNOR2_X1 U650 ( .A(n570), .B(KEYINPUT106), .ZN(n556) );
  NOR2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U652 ( .A(n557), .B(KEYINPUT33), .ZN(n689) );
  NAND2_X1 U653 ( .A1(n562), .A2(n390), .ZN(n563) );
  NOR2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n650) );
  INV_X1 U655 ( .A(n565), .ZN(n567) );
  NAND2_X1 U656 ( .A1(n567), .A2(n568), .ZN(n566) );
  XNOR2_X2 U657 ( .A(n566), .B(KEYINPUT103), .ZN(n669) );
  NOR2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n671) );
  NOR2_X1 U659 ( .A1(n669), .A2(n671), .ZN(n569) );
  INV_X1 U660 ( .A(n624), .ZN(n580) );
  NOR2_X1 U661 ( .A1(n356), .A2(n574), .ZN(n571) );
  XOR2_X1 U662 ( .A(KEYINPUT99), .B(n571), .Z(n703) );
  INV_X1 U663 ( .A(n572), .ZN(n576) );
  NAND2_X1 U664 ( .A1(n703), .A2(n576), .ZN(n573) );
  XNOR2_X1 U665 ( .A(KEYINPUT31), .B(n573), .ZN(n672) );
  INV_X1 U666 ( .A(n574), .ZN(n700) );
  NAND2_X1 U667 ( .A1(n576), .A2(n374), .ZN(n577) );
  XOR2_X1 U668 ( .A(KEYINPUT97), .B(n577), .Z(n578) );
  NOR2_X1 U669 ( .A1(n700), .A2(n578), .ZN(n653) );
  NOR2_X1 U670 ( .A1(n672), .A2(n653), .ZN(n579) );
  NOR2_X1 U671 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U672 ( .A1(n650), .A2(n581), .ZN(n582) );
  XOR2_X1 U673 ( .A(KEYINPUT77), .B(KEYINPUT39), .Z(n591) );
  OR2_X1 U674 ( .A1(n762), .A2(n583), .ZN(n584) );
  NOR2_X1 U675 ( .A1(G900), .A2(n584), .ZN(n585) );
  NOR2_X1 U676 ( .A1(n586), .A2(n585), .ZN(n597) );
  INV_X1 U677 ( .A(n597), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT38), .B(KEYINPUT81), .ZN(n587) );
  AND2_X1 U679 ( .A1(n603), .A2(n379), .ZN(n590) );
  NAND2_X1 U680 ( .A1(n682), .A2(n681), .ZN(n686) );
  INV_X1 U681 ( .A(KEYINPUT41), .ZN(n593) );
  XNOR2_X1 U682 ( .A(n594), .B(n593), .ZN(n679) );
  NAND2_X1 U683 ( .A1(n564), .A2(n693), .ZN(n596) );
  NOR2_X1 U684 ( .A1(n597), .A2(n596), .ZN(n615) );
  AND2_X1 U685 ( .A1(n700), .A2(n615), .ZN(n599) );
  XNOR2_X1 U686 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n598) );
  XNOR2_X1 U687 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U688 ( .A1(n679), .A2(n608), .ZN(n601) );
  NOR2_X1 U689 ( .A1(n604), .A2(n481), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n430), .A2(n605), .ZN(n664) );
  NAND2_X1 U691 ( .A1(KEYINPUT47), .A2(n685), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n664), .A2(n606), .ZN(n607) );
  INV_X1 U693 ( .A(n377), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n608), .A2(n610), .ZN(n665) );
  NAND2_X1 U695 ( .A1(KEYINPUT47), .A2(n665), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n480), .A2(n611), .ZN(n612) );
  INV_X1 U697 ( .A(n669), .ZN(n666) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U699 ( .A(KEYINPUT111), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n628), .B(n617), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n619), .A2(n385), .ZN(n620) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT36), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n622), .A2(n630), .ZN(n675) );
  NAND2_X1 U704 ( .A1(n623), .A2(n675), .ZN(n627) );
  NOR2_X1 U705 ( .A1(KEYINPUT47), .A2(n665), .ZN(n625) );
  XNOR2_X1 U706 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n628), .A2(n681), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  INV_X1 U709 ( .A(n430), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n678) );
  NAND2_X1 U711 ( .A1(n671), .A2(n636), .ZN(n676) );
  NAND2_X1 U712 ( .A1(n678), .A2(n676), .ZN(n637) );
  INV_X1 U713 ( .A(KEYINPUT66), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n387), .A2(G472), .ZN(n644) );
  XOR2_X1 U715 ( .A(n642), .B(KEYINPUT62), .Z(n643) );
  XOR2_X1 U716 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n648) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT94), .ZN(n647) );
  XOR2_X1 U718 ( .A(G101), .B(n650), .Z(G3) );
  NAND2_X1 U719 ( .A1(n653), .A2(n669), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT112), .ZN(n652) );
  XNOR2_X1 U721 ( .A(G104), .B(n652), .ZN(G6) );
  XOR2_X1 U722 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n655) );
  NAND2_X1 U723 ( .A1(n653), .A2(n671), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(n657) );
  XOR2_X1 U725 ( .A(G107), .B(KEYINPUT27), .Z(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G9) );
  XOR2_X1 U727 ( .A(G110), .B(n550), .Z(G12) );
  INV_X1 U728 ( .A(n671), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n659), .A2(n665), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(G128), .B(n662), .ZN(G30) );
  XOR2_X1 U733 ( .A(G143), .B(KEYINPUT115), .Z(n663) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(G45) );
  NOR2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U736 ( .A(G146), .B(n667), .Z(n668) );
  XNOR2_X1 U737 ( .A(KEYINPUT116), .B(n668), .ZN(G48) );
  NAND2_X1 U738 ( .A1(n672), .A2(n669), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n670), .B(G113), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n673), .B(G116), .ZN(G18) );
  XOR2_X1 U742 ( .A(G125), .B(KEYINPUT37), .Z(n674) );
  XNOR2_X1 U743 ( .A(n675), .B(n674), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G134), .B(n676), .ZN(G36) );
  XOR2_X1 U745 ( .A(G140), .B(KEYINPUT117), .Z(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(G42) );
  INV_X1 U747 ( .A(n679), .ZN(n706) );
  NOR2_X1 U748 ( .A1(n394), .A2(n706), .ZN(n680) );
  NOR2_X1 U749 ( .A1(G953), .A2(n680), .ZN(n720) );
  NOR2_X1 U750 ( .A1(n379), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n683), .B(KEYINPUT120), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n592), .A2(n684), .ZN(n688) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n690), .A2(n394), .ZN(n708) );
  NAND2_X1 U756 ( .A1(n691), .A2(n390), .ZN(n692) );
  XNOR2_X1 U757 ( .A(KEYINPUT50), .B(n692), .ZN(n698) );
  XOR2_X1 U758 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n696) );
  OR2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT119), .B(n701), .Z(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U765 ( .A(KEYINPUT51), .B(n704), .Z(n705) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U768 ( .A(n709), .B(KEYINPUT52), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n718) );
  OR2_X1 U770 ( .A1(n760), .A2(KEYINPUT2), .ZN(n712) );
  XNOR2_X1 U771 ( .A(n712), .B(KEYINPUT88), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n392), .A2(n462), .ZN(n713) );
  NAND2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U777 ( .A(n721), .B(KEYINPUT53), .ZN(n722) );
  XNOR2_X1 U778 ( .A(KEYINPUT121), .B(n722), .ZN(G75) );
  XOR2_X1 U779 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n723) );
  XOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  XNOR2_X1 U781 ( .A(n726), .B(KEYINPUT122), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(n731) );
  BUF_X2 U783 ( .A(n729), .Z(n735) );
  NAND2_X1 U784 ( .A1(G469), .A2(n735), .ZN(n730) );
  XOR2_X1 U785 ( .A(n732), .B(KEYINPUT123), .Z(n734) );
  NAND2_X1 U786 ( .A1(G478), .A2(n735), .ZN(n733) );
  NAND2_X1 U787 ( .A1(n735), .A2(G217), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n736), .B(n375), .ZN(n738) );
  NOR2_X1 U789 ( .A1(n739), .A2(n738), .ZN(G66) );
  NAND2_X1 U790 ( .A1(G953), .A2(G224), .ZN(n740) );
  XOR2_X1 U791 ( .A(KEYINPUT61), .B(n740), .Z(n741) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(n745) );
  NOR2_X1 U793 ( .A1(G953), .A2(n392), .ZN(n744) );
  NOR2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n752) );
  XOR2_X1 U795 ( .A(G101), .B(n746), .Z(n747) );
  XNOR2_X1 U796 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U799 ( .A(KEYINPUT124), .B(n753), .ZN(G69) );
  XOR2_X1 U800 ( .A(n754), .B(n755), .Z(n759) );
  XNOR2_X1 U801 ( .A(G227), .B(n759), .ZN(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(G900), .ZN(n757) );
  XNOR2_X1 U803 ( .A(n757), .B(KEYINPUT126), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n758), .A2(G953), .ZN(n765) );
  XNOR2_X1 U805 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U806 ( .A(n761), .B(KEYINPUT125), .ZN(n763) );
  NAND2_X1 U807 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U808 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U809 ( .A(KEYINPUT127), .B(n766), .Z(G72) );
  XNOR2_X1 U810 ( .A(G137), .B(n767), .ZN(G39) );
  XNOR2_X1 U811 ( .A(n391), .B(G122), .ZN(G24) );
  XOR2_X1 U812 ( .A(n389), .B(G119), .Z(G21) );
  XNOR2_X1 U813 ( .A(n373), .B(G131), .ZN(G33) );
endmodule

