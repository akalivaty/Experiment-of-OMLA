//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n195));
  INV_X1    g009(.A(G110), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(new_n198), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n199), .A2(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G125), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(G146), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n206), .A2(KEYINPUT81), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(new_n211), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n202), .A2(new_n203), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n210), .B1(new_n215), .B2(new_n208), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n219), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n224), .B2(new_n211), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n194), .A2(new_n198), .A3(new_n195), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT78), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n194), .A2(new_n195), .A3(new_n228), .A4(new_n198), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(G110), .A3(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n225), .A2(KEYINPUT79), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT79), .B1(new_n225), .B2(new_n230), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n221), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND2_X1  g048(.A1(G221), .A2(G234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT82), .B1(new_n235), .B2(G953), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G221), .A4(G234), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n236), .B2(new_n239), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n234), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(G137), .A3(new_n241), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n233), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n225), .A2(new_n230), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n225), .A2(KEYINPUT79), .A3(new_n230), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n247), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n221), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n255), .A3(new_n188), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n248), .A2(new_n255), .A3(new_n188), .A4(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n190), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n248), .A2(new_n255), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n263), .A2(G902), .A3(new_n189), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G472), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n219), .A2(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n271), .B(new_n272), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n219), .A2(G143), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n267), .A2(G146), .ZN(new_n280));
  OAI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(new_n274), .B2(new_n273), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n272), .B1(new_n281), .B2(new_n271), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT11), .B1(new_n284), .B2(G137), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT11), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n234), .A3(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n234), .B2(G134), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(KEYINPUT64), .A3(G137), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT65), .A2(G131), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n288), .B2(new_n292), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT71), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n288), .A2(new_n292), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n293), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n283), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n191), .B1(new_n279), .B2(new_n280), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n268), .A3(new_n269), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n279), .A2(KEYINPUT1), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G131), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n234), .A2(G134), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n284), .A2(G137), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n285), .A2(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n311), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n304), .A2(KEYINPUT72), .A3(new_n306), .A4(new_n307), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT2), .B(G113), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  XOR2_X1   g135(.A(G116), .B(G119), .Z(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(KEYINPUT68), .ZN(new_n323));
  XNOR2_X1  g137(.A(G116), .B(G119), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT69), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n320), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(KEYINPUT68), .A3(new_n321), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT69), .B1(new_n324), .B2(new_n325), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n319), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n303), .A2(new_n318), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT76), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT76), .B1(new_n332), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n330), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n281), .A2(new_n271), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n299), .A2(new_n340), .A3(new_n301), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n288), .A2(new_n292), .A3(new_n311), .ZN(new_n342));
  INV_X1    g156(.A(new_n314), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n308), .A2(new_n342), .A3(KEYINPUT66), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT66), .B1(new_n316), .B2(new_n308), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n332), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT74), .B(KEYINPUT28), .Z(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n338), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n238), .A3(G210), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(G101), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(G101), .B1(new_n359), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n353), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT73), .A3(new_n361), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n349), .B1(new_n332), .B2(new_n347), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n338), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n337), .A2(new_n352), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n361), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n345), .B2(new_n346), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT67), .B(new_n373), .C1(new_n345), .C2(new_n346), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n303), .A2(KEYINPUT30), .A3(new_n318), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n376), .A2(new_n339), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n332), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n372), .B1(new_n380), .B2(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n332), .A2(new_n333), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n334), .ZN(new_n385));
  INV_X1    g199(.A(new_n332), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n331), .B1(new_n303), .B2(new_n318), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT28), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT77), .B(KEYINPUT28), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n371), .B(new_n381), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n266), .B1(new_n394), .B2(new_n188), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT31), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n386), .A2(new_n372), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n379), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n379), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n384), .B(new_n334), .C1(new_n338), .C2(new_n369), .ZN(new_n401));
  INV_X1    g215(.A(new_n370), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n367), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(G472), .A2(G902), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT32), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n405), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n367), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n351), .A2(new_n335), .A3(new_n336), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(new_n370), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n379), .A2(new_n397), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT31), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n379), .A2(new_n396), .A3(new_n397), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n410), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n265), .B1(new_n407), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT9), .B(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(G221), .B1(new_n420), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT84), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n238), .A2(G227), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND2_X1  g241(.A1(new_n297), .A2(new_n302), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n431));
  INV_X1    g245(.A(G107), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT85), .A2(G107), .ZN(new_n434));
  AOI21_X1  g248(.A(G104), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(G104), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G101), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n439));
  INV_X1    g253(.A(G104), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT3), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n433), .A3(new_n434), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT3), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(G104), .B2(new_n432), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(G101), .B1(new_n440), .B2(G107), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n438), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n439), .B1(new_n438), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n430), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n451));
  INV_X1    g265(.A(G101), .ZN(new_n452));
  AND2_X1   g266(.A1(KEYINPUT85), .A2(G107), .ZN(new_n453));
  NOR2_X1   g267(.A1(KEYINPUT85), .A2(G107), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n440), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n452), .B1(new_n455), .B2(new_n436), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT86), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n438), .A2(new_n447), .A3(new_n439), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(KEYINPUT87), .A3(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n310), .A2(new_n317), .A3(KEYINPUT10), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(G107), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n442), .A2(new_n445), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT4), .A3(G101), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n453), .A2(new_n454), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n444), .B1(new_n466), .B2(new_n441), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n452), .B1(new_n467), .B2(new_n463), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT4), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n467), .B2(new_n446), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n465), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT10), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n308), .A2(new_n438), .A3(new_n447), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n471), .A2(new_n283), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n461), .A2(new_n462), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n462), .B1(new_n461), .B2(new_n474), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n429), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT89), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n479), .B(new_n429), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n461), .A2(new_n428), .A3(new_n474), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n427), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR3_X1    g297(.A1(new_n448), .A2(new_n449), .A3(new_n308), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n473), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n485), .A2(KEYINPUT12), .A3(new_n299), .A4(new_n301), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n428), .B1(new_n484), .B2(new_n473), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(KEYINPUT12), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n482), .A2(new_n427), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n423), .B(new_n188), .C1(new_n483), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n423), .A2(new_n188), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n427), .B1(new_n488), .B2(new_n482), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n481), .B2(new_n490), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n496), .B2(G469), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n422), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G214), .B1(G237), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g315(.A(G113), .ZN(new_n502));
  INV_X1    g316(.A(G116), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n504), .B2(new_n197), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n501), .A2(new_n505), .B1(new_n319), .B2(new_n324), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n450), .A2(new_n459), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n471), .A2(new_n339), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G110), .B(G122), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT90), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n514), .ZN(new_n515));
  MUX2_X1   g329(.A(new_n340), .B(new_n308), .S(new_n213), .Z(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT91), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n238), .A2(G224), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n509), .A2(new_n520), .A3(new_n512), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n516), .B(new_n523), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n457), .A2(new_n458), .A3(new_n506), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n511), .B(KEYINPUT8), .Z(new_n526));
  NOR3_X1   g340(.A1(new_n506), .A2(new_n451), .A3(new_n456), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n524), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G902), .B1(new_n529), .B2(new_n514), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G210), .B1(G237), .B2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n530), .A3(new_n532), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n500), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n537));
  NOR2_X1   g351(.A1(G237), .A2(G953), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G214), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n267), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(G143), .A3(G214), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n537), .B1(new_n542), .B2(G131), .ZN(new_n543));
  AOI211_X1 g357(.A(KEYINPUT92), .B(new_n311), .C1(new_n540), .C2(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT17), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n541), .ZN(new_n546));
  AOI21_X1  g360(.A(G143), .B1(new_n538), .B2(G214), .ZN(new_n547));
  OAI21_X1  g361(.A(G131), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT92), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(new_n537), .A3(G131), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n540), .A2(new_n311), .A3(new_n541), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n211), .ZN(new_n554));
  AOI21_X1  g368(.A(G146), .B1(new_n207), .B2(new_n210), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n545), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G113), .B(G122), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n440), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n220), .B1(new_n219), .B2(new_n206), .ZN(new_n560));
  NAND2_X1  g374(.A1(KEYINPUT18), .A2(G131), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n540), .A2(new_n541), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n542), .A2(KEYINPUT18), .A3(G131), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n557), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n559), .B1(new_n557), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n188), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G475), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT19), .B1(new_n217), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT81), .B1(new_n571), .B2(KEYINPUT19), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n215), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n219), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n211), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n559), .B1(new_n576), .B2(new_n564), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n569), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT20), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT20), .ZN(new_n580));
  INV_X1    g394(.A(new_n577), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n557), .A2(new_n559), .A3(new_n564), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n583), .B2(new_n569), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n568), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n586));
  INV_X1    g400(.A(G122), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(G116), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n503), .A2(KEYINPUT94), .A3(G122), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT14), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(G116), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT14), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n593), .A3(new_n589), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G107), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n466), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n267), .A2(G128), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n191), .A2(G143), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G134), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n599), .A3(new_n284), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n503), .A2(KEYINPUT94), .A3(G122), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT94), .B1(new_n503), .B2(G122), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n592), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n466), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n597), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n602), .A2(KEYINPUT95), .ZN(new_n612));
  XNOR2_X1  g426(.A(G128), .B(G143), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n284), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(KEYINPUT13), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n191), .A2(G143), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT13), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n284), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n612), .A2(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(new_n611), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n611), .B1(new_n610), .B2(new_n620), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n604), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n420), .A2(new_n187), .A3(G953), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT97), .Z(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n610), .A2(new_n620), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n621), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n631), .B2(new_n604), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n188), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT15), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n634), .A3(G478), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n624), .A2(new_n626), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n631), .A2(new_n628), .A3(new_n604), .ZN(new_n637));
  AOI21_X1  g451(.A(G902), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G478), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(KEYINPUT15), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(G234), .A2(G237), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n642), .A2(G952), .A3(new_n238), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(G902), .A3(G953), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT98), .Z(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT21), .B(G898), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n585), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n536), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n419), .A2(new_n498), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G101), .ZN(G3));
  NAND2_X1  g466(.A1(new_n493), .A2(new_n497), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n266), .B1(new_n404), .B2(new_n188), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n408), .B1(new_n400), .B2(new_n403), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n265), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n653), .A2(new_n656), .A3(new_n421), .ZN(new_n657));
  INV_X1    g471(.A(new_n647), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n536), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n603), .A2(new_n597), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(G107), .B2(new_n595), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n630), .B2(new_n621), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n628), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n624), .A2(KEYINPUT99), .A3(new_n626), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT33), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n664), .A2(new_n665), .A3(new_n668), .A4(KEYINPUT33), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT33), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n627), .B2(new_n632), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n639), .A2(G902), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n669), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n633), .A2(new_n674), .A3(new_n639), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT101), .B1(new_n638), .B2(G478), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n578), .A2(KEYINPUT20), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n583), .A2(new_n580), .A3(new_n569), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n673), .A2(new_n677), .B1(new_n680), .B2(new_n568), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n659), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n657), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT34), .B(G104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G6));
  INV_X1    g502(.A(new_n641), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n585), .A3(new_n647), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n522), .A2(new_n532), .A3(new_n530), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n532), .B1(new_n522), .B2(new_n530), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n499), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n657), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT35), .B(G107), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  OR2_X1    g513(.A1(new_n654), .A2(new_n655), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n259), .A2(new_n261), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n189), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT36), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n254), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n233), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n253), .A2(new_n707), .A3(new_n221), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n189), .A2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT105), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n702), .A2(new_n703), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n710), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n714), .B2(new_n262), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n498), .A3(new_n650), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT37), .B(G110), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G12));
  NAND2_X1  g534(.A1(new_n394), .A2(new_n188), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  INV_X1    g536(.A(new_n406), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n418), .ZN(new_n724));
  INV_X1    g538(.A(G900), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n643), .B1(new_n645), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n689), .A2(new_n585), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n716), .A2(new_n695), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n498), .A2(new_n724), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G128), .ZN(G30));
  XOR2_X1   g544(.A(new_n726), .B(KEYINPUT39), .Z(new_n731));
  NAND2_X1  g545(.A1(new_n498), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT40), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n367), .B1(new_n386), .B2(new_n387), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n414), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n188), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G472), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n418), .B(new_n738), .C1(new_n655), .C2(KEYINPUT32), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n693), .A2(new_n694), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT38), .Z(new_n741));
  NOR2_X1   g555(.A1(new_n714), .A2(new_n262), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n680), .A2(new_n568), .B1(new_n635), .B2(new_n640), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n499), .A2(new_n741), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G143), .ZN(G45));
  NAND2_X1  g560(.A1(new_n673), .A2(new_n677), .ZN(new_n747));
  INV_X1    g561(.A(new_n726), .ZN(new_n748));
  AND4_X1   g562(.A1(KEYINPUT107), .A2(new_n747), .A3(new_n585), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n681), .B2(new_n748), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n498), .A2(new_n751), .A3(new_n724), .A4(new_n728), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  NAND2_X1  g567(.A1(new_n461), .A2(new_n474), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT88), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n461), .A2(new_n462), .A3(new_n474), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n479), .B1(new_n757), .B2(new_n429), .ZN(new_n758));
  INV_X1    g572(.A(new_n480), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n482), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n427), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n492), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n762), .B2(G902), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n764));
  INV_X1    g578(.A(new_n482), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n478), .B2(new_n480), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n491), .B1(new_n766), .B2(new_n427), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n423), .B1(new_n767), .B2(new_n188), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n493), .A2(new_n421), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n419), .A3(new_n683), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n772), .B1(new_n764), .B2(new_n770), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT109), .A3(new_n419), .A4(new_n683), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT41), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G113), .ZN(G15));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n419), .A3(new_n696), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G116), .ZN(G18));
  INV_X1    g597(.A(new_n410), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n400), .B2(new_n403), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n395), .A2(new_n406), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n716), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n777), .A2(new_n787), .A3(new_n648), .A4(new_n536), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G119), .ZN(G21));
  NAND2_X1  g603(.A1(new_n390), .A2(new_n391), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n411), .B1(new_n790), .B2(new_n337), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n405), .B1(new_n791), .B2(new_n417), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n262), .A2(new_n264), .ZN(new_n793));
  AOI21_X1  g607(.A(G902), .B1(new_n400), .B2(new_n403), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n266), .ZN(new_n795));
  INV_X1    g609(.A(new_n743), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n659), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n771), .A2(new_n797), .A3(new_n773), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G122), .ZN(G24));
  NAND2_X1  g613(.A1(new_n702), .A2(new_n711), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n792), .B(new_n800), .C1(new_n266), .C2(new_n794), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n749), .A3(new_n750), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n771), .A2(new_n536), .A3(new_n802), .A4(new_n773), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G125), .ZN(G27));
  NAND2_X1  g618(.A1(new_n740), .A2(new_n499), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n498), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n419), .A3(new_n751), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT42), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n785), .B(KEYINPUT110), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n265), .B1(new_n811), .B2(new_n407), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n807), .A2(KEYINPUT42), .A3(new_n751), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G131), .ZN(G33));
  NAND4_X1  g629(.A1(new_n419), .A2(new_n498), .A3(new_n727), .A4(new_n806), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G134), .ZN(G36));
  AOI21_X1  g631(.A(new_n585), .B1(new_n747), .B2(KEYINPUT112), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(KEYINPUT112), .B2(new_n747), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT43), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n585), .B(KEYINPUT113), .Z(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(KEYINPUT43), .A3(new_n747), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n700), .A3(new_n800), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT44), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n805), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n496), .A2(KEYINPUT45), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n496), .A2(KEYINPUT45), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(G469), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n831), .A2(KEYINPUT111), .A3(G469), .A4(new_n832), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n494), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(KEYINPUT46), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n493), .B1(new_n837), .B2(KEYINPUT46), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n421), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n828), .A2(new_n829), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n830), .A2(new_n731), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G137), .ZN(G39));
  NAND2_X1  g658(.A1(new_n840), .A2(KEYINPUT47), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT47), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n421), .C1(new_n838), .C2(new_n839), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n724), .A2(new_n793), .A3(new_n805), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n751), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G140), .ZN(G42));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n824), .A2(new_n643), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(new_n795), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(new_n805), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n847), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n771), .A2(new_n493), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n855), .A2(KEYINPUT119), .B1(new_n422), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n854), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n777), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n853), .A2(new_n499), .A3(new_n741), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n777), .A2(new_n806), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n868), .A2(new_n852), .A3(KEYINPUT122), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT122), .B1(new_n868), .B2(new_n852), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n801), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n643), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n739), .A2(new_n265), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n777), .A2(new_n806), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n585), .A3(new_n747), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n851), .B1(new_n861), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n768), .A2(new_n769), .ZN(new_n879));
  AOI211_X1 g693(.A(KEYINPUT108), .B(new_n423), .C1(new_n767), .C2(new_n188), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n773), .B(new_n536), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n853), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(G953), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n869), .A2(new_n870), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT48), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n812), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n885), .B2(new_n812), .ZN(new_n888));
  OAI221_X1 g702(.A(new_n884), .B1(new_n682), .B2(new_n874), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n871), .ZN(new_n890));
  INV_X1    g704(.A(new_n875), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT123), .B1(new_n871), .B2(new_n875), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n859), .A2(new_n422), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n854), .B1(new_n855), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT51), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n865), .B1(new_n866), .B2(new_n851), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n878), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n802), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n729), .B(new_n752), .C1(new_n881), .C2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n499), .B(new_n743), .C1(new_n693), .C2(new_n694), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n800), .A2(new_n726), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n906), .A2(new_n739), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n498), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT116), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n752), .A2(new_n729), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n803), .A4(new_n909), .ZN(new_n914));
  INV_X1    g728(.A(new_n803), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n498), .A2(new_n739), .A3(new_n906), .A4(new_n907), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n752), .A2(new_n729), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n904), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n911), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n585), .A2(new_n641), .A3(new_n726), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n740), .A2(new_n499), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT115), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n740), .A2(KEYINPUT115), .A3(new_n499), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n787), .A2(new_n925), .A3(new_n498), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n802), .A2(new_n498), .A3(new_n806), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n816), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n810), .B2(new_n813), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n788), .A2(new_n782), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n689), .A2(new_n585), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n681), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n659), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n498), .A3(new_n656), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n798), .A2(new_n651), .A3(new_n718), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n929), .A2(new_n936), .A3(new_n779), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT53), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n919), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n752), .A2(new_n729), .A3(new_n916), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT52), .B1(new_n940), .B2(new_n803), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n536), .A2(new_n715), .A3(new_n712), .A4(new_n727), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n786), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n498), .B1(new_n943), .B2(new_n908), .ZN(new_n944));
  AND4_X1   g758(.A1(KEYINPUT52), .A2(new_n803), .A3(new_n944), .A4(new_n752), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT117), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n776), .A2(new_n778), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n777), .A2(new_n797), .B1(new_n657), .B2(new_n933), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n498), .B(new_n650), .C1(new_n419), .C2(new_n717), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n782), .A3(new_n788), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT117), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n803), .A2(new_n944), .A3(KEYINPUT52), .A4(new_n752), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n918), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n946), .A2(new_n951), .A3(new_n929), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n939), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT54), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n955), .A2(KEYINPUT118), .A3(new_n938), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n938), .B1(new_n919), .B2(new_n937), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n938), .B2(new_n955), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT54), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  OAI22_X1  g779(.A1(new_n901), .A2(new_n965), .B1(G952), .B2(G953), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n265), .A2(new_n422), .A3(new_n500), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n747), .A3(new_n822), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n741), .A2(new_n970), .A3(new_n739), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n966), .A2(new_n972), .ZN(G75));
  NAND2_X1  g787(.A1(new_n956), .A2(new_n957), .ZN(new_n974));
  INV_X1    g788(.A(new_n939), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n960), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(G210), .A3(G902), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT56), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n515), .A2(new_n521), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n519), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT55), .Z(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n977), .B2(new_n978), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n238), .A2(G952), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(G51));
  XNOR2_X1  g799(.A(new_n494), .B(KEYINPUT57), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n959), .A2(new_n974), .A3(new_n960), .A4(new_n975), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n767), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n188), .B1(new_n958), .B2(new_n960), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n835), .A3(new_n836), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n984), .B1(new_n990), .B2(new_n992), .ZN(G54));
  NAND3_X1  g807(.A1(new_n991), .A2(KEYINPUT58), .A3(G475), .ZN(new_n994));
  INV_X1    g808(.A(new_n583), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n984), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n991), .A2(KEYINPUT58), .A3(G475), .A4(new_n583), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(G60));
  NAND3_X1  g813(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G478), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT59), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1001), .B1(new_n965), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n976), .A2(KEYINPUT54), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n961), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1005), .A2(new_n1008), .A3(new_n984), .ZN(G63));
  NAND2_X1  g823(.A1(G217), .A2(G902), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT60), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n976), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n984), .B1(new_n1013), .B2(new_n263), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1011), .B1(new_n958), .B2(new_n960), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n706), .A2(new_n708), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1014), .A2(KEYINPUT61), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT61), .ZN(new_n1019));
  INV_X1    g833(.A(new_n263), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n997), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n976), .A2(new_n1016), .A3(new_n1012), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1018), .A2(new_n1023), .ZN(G66));
  INV_X1    g838(.A(new_n951), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G224), .A2(G953), .ZN(new_n1026));
  OAI22_X1  g840(.A1(new_n1025), .A2(G953), .B1(new_n646), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(G898), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n979), .B1(new_n1028), .B2(G953), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1027), .B(new_n1029), .ZN(G69));
  INV_X1    g844(.A(new_n419), .ZN(new_n1031));
  NOR4_X1   g845(.A1(new_n1031), .A2(new_n732), .A3(new_n805), .A4(new_n932), .ZN(new_n1032));
  INV_X1    g846(.A(new_n903), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n745), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n745), .A2(new_n1033), .A3(KEYINPUT62), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n843), .A2(new_n1038), .A3(new_n849), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n238), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n572), .A2(new_n574), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(KEYINPUT124), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT124), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1040), .A2(new_n1047), .A3(new_n1044), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n841), .A2(new_n731), .A3(new_n812), .A4(new_n906), .ZN(new_n1049));
  AND4_X1   g863(.A1(new_n814), .A2(new_n1049), .A3(new_n816), .A4(new_n1033), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1050), .A2(new_n238), .A3(new_n843), .A4(new_n849), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1044), .B1(G900), .B2(G953), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1046), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n238), .B1(G227), .B2(G900), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1055), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1046), .A2(new_n1057), .A3(new_n1053), .A4(new_n1048), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1056), .A2(new_n1058), .ZN(G72));
  INV_X1    g873(.A(new_n380), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(new_n372), .ZN(new_n1061));
  NOR2_X1   g875(.A1(new_n1060), .A2(new_n372), .ZN(new_n1062));
  XNOR2_X1  g876(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n266), .A2(new_n188), .ZN(new_n1064));
  XNOR2_X1  g878(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NOR2_X1   g879(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n963), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g881(.A(new_n1067), .B(KEYINPUT127), .ZN(new_n1068));
  XNOR2_X1  g882(.A(new_n1061), .B(KEYINPUT126), .ZN(new_n1069));
  AND4_X1   g883(.A1(new_n843), .A2(new_n1050), .A3(new_n849), .A4(new_n951), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1069), .B1(new_n1070), .B2(new_n1065), .ZN(new_n1071));
  INV_X1    g885(.A(new_n1065), .ZN(new_n1072));
  OAI21_X1  g886(.A(new_n1072), .B1(new_n1039), .B2(new_n1025), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n984), .B1(new_n1073), .B2(new_n1062), .ZN(new_n1074));
  AND3_X1   g888(.A1(new_n1068), .A2(new_n1071), .A3(new_n1074), .ZN(G57));
endmodule


