

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764;

  OR2_X1 U378 ( .A1(G902), .A2(n723), .ZN(n356) );
  OR2_X1 U379 ( .A1(n634), .A2(G902), .ZN(n521) );
  INV_X1 U380 ( .A(G131), .ZN(n425) );
  NOR2_X1 U381 ( .A1(n719), .A2(G902), .ZN(n508) );
  INV_X1 U382 ( .A(G953), .ZN(n753) );
  XNOR2_X2 U383 ( .A(G478), .B(n356), .ZN(n543) );
  XNOR2_X2 U384 ( .A(n408), .B(n593), .ZN(n764) );
  INV_X2 U385 ( .A(n623), .ZN(n707) );
  XNOR2_X2 U386 ( .A(n427), .B(n426), .ZN(n623) );
  XNOR2_X2 U387 ( .A(n441), .B(KEYINPUT4), .ZN(n742) );
  NOR2_X1 U388 ( .A1(G953), .A2(n733), .ZN(n734) );
  NOR2_X1 U389 ( .A1(n532), .A2(n580), .ZN(n534) );
  NAND2_X2 U390 ( .A1(n707), .A2(n626), .ZN(n372) );
  AND2_X1 U391 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U392 ( .A(n534), .B(n533), .ZN(n762) );
  INV_X1 U393 ( .A(n672), .ZN(n367) );
  XNOR2_X1 U394 ( .A(n611), .B(n587), .ZN(n689) );
  OR2_X2 U395 ( .A1(n386), .A2(n385), .ZN(n679) );
  NOR2_X2 U396 ( .A1(n543), .A2(n423), .ZN(n663) );
  AND2_X1 U397 ( .A1(n403), .A2(n402), .ZN(n401) );
  OR2_X1 U398 ( .A1(n629), .A2(n398), .ZN(n397) );
  XNOR2_X1 U399 ( .A(n743), .B(G110), .ZN(n510) );
  XNOR2_X2 U400 ( .A(n431), .B(n430), .ZN(n757) );
  XNOR2_X2 U401 ( .A(n741), .B(n424), .ZN(n505) );
  XNOR2_X2 U402 ( .A(n425), .B(G134), .ZN(n741) );
  XNOR2_X2 U403 ( .A(n562), .B(KEYINPUT1), .ZN(n526) );
  XNOR2_X2 U404 ( .A(n508), .B(n507), .ZN(n562) );
  OR2_X1 U405 ( .A1(G237), .A2(G902), .ZN(n457) );
  INV_X1 U406 ( .A(KEYINPUT15), .ZN(n456) );
  NAND2_X2 U407 ( .A1(n379), .A2(n377), .ZN(n624) );
  NAND2_X1 U408 ( .A1(n378), .A2(KEYINPUT78), .ZN(n377) );
  INV_X1 U409 ( .A(KEYINPUT6), .ZN(n420) );
  XNOR2_X1 U410 ( .A(n503), .B(n445), .ZN(n498) );
  AND2_X1 U411 ( .A1(n560), .A2(n679), .ZN(n561) );
  XNOR2_X1 U412 ( .A(n410), .B(KEYINPUT47), .ZN(n409) );
  XNOR2_X1 U413 ( .A(n391), .B(KEYINPUT101), .ZN(n549) );
  NOR2_X1 U414 ( .A1(n535), .A2(n550), .ZN(n429) );
  OR2_X1 U415 ( .A1(n762), .A2(KEYINPUT44), .ZN(n535) );
  XOR2_X1 U416 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n462) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n491) );
  XNOR2_X1 U418 ( .A(G125), .B(G146), .ZN(n466) );
  NOR2_X1 U419 ( .A1(n419), .A2(n422), .ZN(n606) );
  NAND2_X1 U420 ( .A1(n663), .A2(n560), .ZN(n422) );
  AND2_X1 U421 ( .A1(n526), .A2(n367), .ZN(n537) );
  NAND2_X1 U422 ( .A1(n359), .A2(n619), .ZN(n402) );
  NAND2_X1 U423 ( .A1(n396), .A2(n401), .ZN(n559) );
  AND2_X1 U424 ( .A1(n397), .A2(n607), .ZN(n396) );
  INV_X1 U425 ( .A(G146), .ZN(n424) );
  XNOR2_X1 U426 ( .A(G137), .B(G113), .ZN(n493) );
  XNOR2_X1 U427 ( .A(n742), .B(n442), .ZN(n503) );
  INV_X1 U428 ( .A(G101), .ZN(n442) );
  NOR2_X1 U429 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U430 ( .A(KEYINPUT22), .ZN(n490) );
  NAND2_X1 U431 ( .A1(n387), .A2(n390), .ZN(n386) );
  NAND2_X1 U432 ( .A1(n421), .A2(G902), .ZN(n390) );
  NOR2_X1 U433 ( .A1(n523), .A2(n558), .ZN(n546) );
  AND2_X1 U434 ( .A1(n381), .A2(n617), .ZN(n380) );
  NAND2_X1 U435 ( .A1(n763), .A2(KEYINPUT78), .ZN(n381) );
  INV_X1 U436 ( .A(KEYINPUT45), .ZN(n426) );
  INV_X1 U437 ( .A(G234), .ZN(n486) );
  XOR2_X1 U438 ( .A(G113), .B(G104), .Z(n468) );
  XNOR2_X1 U439 ( .A(G143), .B(G122), .ZN(n461) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT83), .ZN(n446) );
  XOR2_X1 U441 ( .A(KEYINPUT71), .B(KEYINPUT17), .Z(n447) );
  NAND2_X1 U442 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U443 ( .A(n575), .B(KEYINPUT105), .ZN(n577) );
  AND2_X1 U444 ( .A1(n676), .A2(n360), .ZN(n560) );
  NAND2_X1 U445 ( .A1(n499), .A2(n389), .ZN(n388) );
  XNOR2_X1 U446 ( .A(KEYINPUT82), .B(KEYINPUT3), .ZN(n443) );
  XOR2_X1 U447 ( .A(G116), .B(G119), .Z(n444) );
  XNOR2_X1 U448 ( .A(G128), .B(G119), .ZN(n513) );
  XNOR2_X1 U449 ( .A(n510), .B(n509), .ZN(n412) );
  XNOR2_X1 U450 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n465) );
  XOR2_X1 U451 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n478) );
  XNOR2_X1 U452 ( .A(G116), .B(G134), .ZN(n477) );
  XNOR2_X1 U453 ( .A(n366), .B(n479), .ZN(n481) );
  XNOR2_X1 U454 ( .A(n404), .B(n480), .ZN(n366) );
  XOR2_X1 U455 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n480) );
  XNOR2_X1 U456 ( .A(n483), .B(KEYINPUT8), .ZN(n511) );
  XOR2_X1 U457 ( .A(G104), .B(KEYINPUT88), .Z(n501) );
  INV_X1 U458 ( .A(KEYINPUT102), .ZN(n527) );
  INV_X1 U459 ( .A(n559), .ZN(n375) );
  XNOR2_X1 U460 ( .A(n606), .B(KEYINPUT110), .ZN(n376) );
  NAND2_X1 U461 ( .A1(n367), .A2(n562), .ZN(n575) );
  XNOR2_X1 U462 ( .A(n498), .B(n497), .ZN(n637) );
  XNOR2_X1 U463 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U464 ( .A(n505), .B(n492), .ZN(n496) );
  AND2_X1 U465 ( .A1(n372), .A2(G475), .ZN(n406) );
  AND2_X1 U466 ( .A1(n372), .A2(G210), .ZN(n405) );
  NAND2_X1 U467 ( .A1(n711), .A2(n372), .ZN(n712) );
  XNOR2_X1 U468 ( .A(n599), .B(KEYINPUT40), .ZN(n643) );
  XNOR2_X1 U469 ( .A(n417), .B(KEYINPUT111), .ZN(n759) );
  NAND2_X1 U470 ( .A1(n418), .A2(n526), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n374), .B(n373), .ZN(n418) );
  INV_X1 U472 ( .A(KEYINPUT36), .ZN(n373) );
  XNOR2_X1 U473 ( .A(KEYINPUT32), .B(KEYINPUT64), .ZN(n430) );
  NAND2_X1 U474 ( .A1(n546), .A2(n522), .ZN(n431) );
  XNOR2_X1 U475 ( .A(n538), .B(n370), .ZN(n667) );
  XNOR2_X1 U476 ( .A(n371), .B(KEYINPUT95), .ZN(n370) );
  INV_X1 U477 ( .A(KEYINPUT31), .ZN(n371) );
  NOR2_X1 U478 ( .A1(n565), .A2(n590), .ZN(n662) );
  XNOR2_X1 U479 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U480 ( .A(n719), .B(n432), .ZN(n720) );
  XNOR2_X1 U481 ( .A(n559), .B(KEYINPUT19), .ZN(n564) );
  XNOR2_X1 U482 ( .A(n679), .B(n420), .ZN(n558) );
  INV_X1 U483 ( .A(n558), .ZN(n419) );
  AND2_X1 U484 ( .A1(n372), .A2(G472), .ZN(n357) );
  AND2_X1 U485 ( .A1(n372), .A2(G217), .ZN(n358) );
  NAND2_X1 U486 ( .A1(G210), .A2(n457), .ZN(n359) );
  AND2_X1 U487 ( .A1(n557), .A2(n576), .ZN(n360) );
  AND2_X1 U488 ( .A1(n673), .A2(n547), .ZN(n361) );
  INV_X1 U489 ( .A(G902), .ZN(n389) );
  XNOR2_X1 U490 ( .A(n456), .B(G902), .ZN(n619) );
  XOR2_X1 U491 ( .A(n629), .B(n628), .Z(n362) );
  XOR2_X1 U492 ( .A(n634), .B(n633), .Z(n363) );
  XOR2_X1 U493 ( .A(n637), .B(n636), .Z(n364) );
  XNOR2_X1 U494 ( .A(KEYINPUT79), .B(KEYINPUT56), .ZN(n365) );
  NAND2_X1 U495 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U496 ( .A1(n764), .A2(n643), .ZN(n601) );
  NAND2_X2 U497 ( .A1(n401), .A2(n397), .ZN(n611) );
  NAND2_X1 U498 ( .A1(n627), .A2(n405), .ZN(n630) );
  XNOR2_X1 U499 ( .A(n368), .B(n365), .ZN(G51) );
  NAND2_X1 U500 ( .A1(n632), .A2(n638), .ZN(n368) );
  XNOR2_X1 U501 ( .A(n369), .B(n504), .ZN(n719) );
  XNOR2_X1 U502 ( .A(n503), .B(n506), .ZN(n369) );
  NAND2_X1 U503 ( .A1(n564), .A2(n459), .ZN(n460) );
  AND2_X1 U504 ( .A1(n627), .A2(n372), .ZN(n407) );
  INV_X1 U505 ( .A(n384), .ZN(n378) );
  NAND2_X1 U506 ( .A1(n384), .A2(n383), .ZN(n382) );
  AND2_X1 U507 ( .A1(n614), .A2(n615), .ZN(n383) );
  XNOR2_X1 U508 ( .A(n605), .B(n604), .ZN(n384) );
  NOR2_X1 U509 ( .A1(n637), .A2(n388), .ZN(n385) );
  NAND2_X1 U510 ( .A1(n637), .A2(n421), .ZN(n387) );
  NAND2_X1 U511 ( .A1(n392), .A2(n644), .ZN(n391) );
  NAND2_X1 U512 ( .A1(n546), .A2(n361), .ZN(n644) );
  NAND2_X1 U513 ( .A1(n393), .A2(n693), .ZN(n392) );
  NAND2_X1 U514 ( .A1(n667), .A2(n652), .ZN(n393) );
  XNOR2_X1 U515 ( .A(n394), .B(n490), .ZN(n523) );
  NOR2_X1 U516 ( .A1(n539), .A2(n395), .ZN(n394) );
  NAND2_X1 U517 ( .A1(n691), .A2(n557), .ZN(n395) );
  INV_X1 U518 ( .A(n619), .ZN(n399) );
  INV_X1 U519 ( .A(n359), .ZN(n400) );
  NAND2_X1 U520 ( .A1(n629), .A2(n359), .ZN(n403) );
  NAND2_X1 U521 ( .A1(n627), .A2(n357), .ZN(n416) );
  INV_X1 U522 ( .A(n441), .ZN(n404) );
  NAND2_X1 U523 ( .A1(n627), .A2(n358), .ZN(n635) );
  NAND2_X1 U524 ( .A1(n627), .A2(n406), .ZN(n647) );
  NAND2_X1 U525 ( .A1(n407), .A2(G469), .ZN(n721) );
  NAND2_X1 U526 ( .A1(n407), .A2(G478), .ZN(n724) );
  NAND2_X1 U527 ( .A1(n687), .A2(n591), .ZN(n408) );
  XNOR2_X2 U528 ( .A(n589), .B(KEYINPUT41), .ZN(n687) );
  NAND2_X1 U529 ( .A1(n409), .A2(n566), .ZN(n569) );
  NAND2_X1 U530 ( .A1(n662), .A2(n693), .ZN(n410) );
  XNOR2_X1 U531 ( .A(n515), .B(n411), .ZN(n634) );
  XNOR2_X1 U532 ( .A(n413), .B(n412), .ZN(n411) );
  NAND2_X1 U533 ( .A1(n511), .A2(G221), .ZN(n413) );
  XNOR2_X2 U534 ( .A(n521), .B(n520), .ZN(n676) );
  XNOR2_X1 U535 ( .A(n414), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U536 ( .A1(n415), .A2(n638), .ZN(n414) );
  XNOR2_X1 U537 ( .A(n635), .B(n363), .ZN(n415) );
  XNOR2_X1 U538 ( .A(n416), .B(n364), .ZN(n639) );
  XNOR2_X1 U539 ( .A(n759), .B(KEYINPUT80), .ZN(n586) );
  INV_X1 U540 ( .A(n543), .ZN(n544) );
  INV_X1 U541 ( .A(n499), .ZN(n421) );
  INV_X1 U542 ( .A(n545), .ZN(n423) );
  NAND2_X1 U543 ( .A1(n552), .A2(n428), .ZN(n427) );
  XNOR2_X1 U544 ( .A(n429), .B(n536), .ZN(n428) );
  XOR2_X1 U545 ( .A(n718), .B(n717), .Z(n432) );
  AND2_X1 U546 ( .A1(n549), .A2(n548), .ZN(n433) );
  INV_X1 U547 ( .A(KEYINPUT46), .ZN(n600) );
  INV_X1 U548 ( .A(KEYINPUT68), .ZN(n536) );
  AND2_X1 U549 ( .A1(n433), .A2(n551), .ZN(n552) );
  INV_X1 U550 ( .A(n727), .ZN(n445) );
  INV_X1 U551 ( .A(KEYINPUT78), .ZN(n615) );
  INV_X1 U552 ( .A(KEYINPUT34), .ZN(n530) );
  INV_X1 U553 ( .A(n726), .ZN(n638) );
  INV_X1 U554 ( .A(KEYINPUT35), .ZN(n533) );
  NOR2_X1 U555 ( .A1(G898), .A2(n753), .ZN(n434) );
  XOR2_X1 U556 ( .A(KEYINPUT86), .B(n434), .Z(n731) );
  NAND2_X1 U557 ( .A1(G234), .A2(G237), .ZN(n435) );
  XNOR2_X1 U558 ( .A(n435), .B(KEYINPUT14), .ZN(n436) );
  XNOR2_X1 U559 ( .A(KEYINPUT70), .B(n436), .ZN(n438) );
  NAND2_X1 U560 ( .A1(G902), .A2(n438), .ZN(n553) );
  NOR2_X1 U561 ( .A1(n731), .A2(n553), .ZN(n437) );
  XNOR2_X1 U562 ( .A(KEYINPUT87), .B(n437), .ZN(n440) );
  NAND2_X1 U563 ( .A1(G952), .A2(n438), .ZN(n703) );
  NOR2_X1 U564 ( .A1(G953), .A2(n703), .ZN(n439) );
  XNOR2_X1 U565 ( .A(n439), .B(KEYINPUT85), .ZN(n556) );
  NAND2_X1 U566 ( .A1(n440), .A2(n556), .ZN(n459) );
  XNOR2_X2 U567 ( .A(G143), .B(G128), .ZN(n441) );
  XNOR2_X1 U568 ( .A(n444), .B(n443), .ZN(n727) );
  XNOR2_X1 U569 ( .A(n447), .B(n446), .ZN(n450) );
  NAND2_X1 U570 ( .A1(G224), .A2(n753), .ZN(n448) );
  XNOR2_X1 U571 ( .A(n466), .B(n448), .ZN(n449) );
  XNOR2_X1 U572 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U573 ( .A(n498), .B(n451), .ZN(n455) );
  XOR2_X1 U574 ( .A(KEYINPUT69), .B(G110), .Z(n453) );
  XOR2_X1 U575 ( .A(G122), .B(G107), .Z(n479) );
  XNOR2_X1 U576 ( .A(n479), .B(n468), .ZN(n452) );
  XNOR2_X1 U577 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U578 ( .A(KEYINPUT16), .B(n454), .ZN(n729) );
  XNOR2_X1 U579 ( .A(n455), .B(n729), .ZN(n629) );
  NAND2_X1 U580 ( .A1(n457), .A2(G214), .ZN(n458) );
  XNOR2_X1 U581 ( .A(n458), .B(KEYINPUT84), .ZN(n607) );
  INV_X1 U582 ( .A(n607), .ZN(n690) );
  XNOR2_X2 U583 ( .A(n460), .B(KEYINPUT0), .ZN(n539) );
  XNOR2_X1 U584 ( .A(n462), .B(n461), .ZN(n464) );
  NAND2_X1 U585 ( .A1(G214), .A2(n491), .ZN(n463) );
  XNOR2_X1 U586 ( .A(n464), .B(n463), .ZN(n467) );
  XNOR2_X1 U587 ( .A(n466), .B(n465), .ZN(n745) );
  XNOR2_X1 U588 ( .A(n467), .B(n745), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n468), .B(G140), .ZN(n472) );
  XOR2_X1 U590 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n470) );
  XNOR2_X1 U591 ( .A(G131), .B(KEYINPUT12), .ZN(n469) );
  XNOR2_X1 U592 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U593 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U594 ( .A(n474), .B(n473), .ZN(n645) );
  NAND2_X1 U595 ( .A1(n645), .A2(n389), .ZN(n476) );
  XOR2_X1 U596 ( .A(KEYINPUT13), .B(G475), .Z(n475) );
  XNOR2_X1 U597 ( .A(n476), .B(n475), .ZN(n545) );
  XNOR2_X1 U598 ( .A(n478), .B(n477), .ZN(n482) );
  XOR2_X1 U599 ( .A(n482), .B(n481), .Z(n485) );
  AND2_X1 U600 ( .A1(G234), .A2(n753), .ZN(n483) );
  NAND2_X1 U601 ( .A1(G217), .A2(n511), .ZN(n484) );
  XNOR2_X1 U602 ( .A(n485), .B(n484), .ZN(n723) );
  NOR2_X1 U603 ( .A1(n545), .A2(n543), .ZN(n691) );
  OR2_X1 U604 ( .A1(n619), .A2(n486), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n487), .B(KEYINPUT20), .ZN(n516) );
  NAND2_X1 U606 ( .A1(n516), .A2(G221), .ZN(n489) );
  INV_X1 U607 ( .A(KEYINPUT21), .ZN(n488) );
  XNOR2_X1 U608 ( .A(n489), .B(n488), .ZN(n557) );
  XNOR2_X1 U609 ( .A(G472), .B(KEYINPUT93), .ZN(n499) );
  NAND2_X1 U610 ( .A1(n491), .A2(G210), .ZN(n492) );
  XOR2_X1 U611 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n494) );
  XNOR2_X1 U612 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U613 ( .A1(G227), .A2(n753), .ZN(n500) );
  XNOR2_X1 U614 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X2 U615 ( .A(G140), .B(G137), .ZN(n743) );
  XOR2_X1 U616 ( .A(n502), .B(n510), .Z(n504) );
  XNOR2_X1 U617 ( .A(n505), .B(G107), .ZN(n506) );
  INV_X1 U618 ( .A(G469), .ZN(n507) );
  INV_X1 U619 ( .A(n526), .ZN(n673) );
  XNOR2_X1 U620 ( .A(KEYINPUT67), .B(KEYINPUT89), .ZN(n509) );
  XNOR2_X1 U621 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U623 ( .A(n745), .B(n514), .ZN(n515) );
  AND2_X1 U624 ( .A1(n516), .A2(G217), .ZN(n519) );
  XNOR2_X1 U625 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n517) );
  XNOR2_X1 U626 ( .A(n517), .B(KEYINPUT25), .ZN(n518) );
  XNOR2_X1 U627 ( .A(n519), .B(n518), .ZN(n520) );
  INV_X1 U628 ( .A(n676), .ZN(n547) );
  NOR2_X1 U629 ( .A1(n673), .A2(n547), .ZN(n522) );
  NOR2_X1 U630 ( .A1(n523), .A2(n526), .ZN(n525) );
  NOR2_X1 U631 ( .A1(n679), .A2(n547), .ZN(n524) );
  NAND2_X1 U632 ( .A1(n525), .A2(n524), .ZN(n657) );
  NAND2_X1 U633 ( .A1(n757), .A2(n657), .ZN(n550) );
  INV_X1 U634 ( .A(n557), .ZN(n675) );
  OR2_X1 U635 ( .A1(n676), .A2(n675), .ZN(n672) );
  XNOR2_X1 U636 ( .A(n537), .B(n527), .ZN(n528) );
  NOR2_X1 U637 ( .A1(n528), .A2(n419), .ZN(n529) );
  XNOR2_X1 U638 ( .A(KEYINPUT33), .B(n529), .ZN(n688) );
  NOR2_X1 U639 ( .A1(n688), .A2(n539), .ZN(n531) );
  XNOR2_X1 U640 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U641 ( .A1(n545), .A2(n543), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n679), .A2(n537), .ZN(n684) );
  NOR2_X1 U643 ( .A1(n539), .A2(n684), .ZN(n538) );
  NOR2_X1 U644 ( .A1(n679), .A2(n539), .ZN(n541) );
  INV_X1 U645 ( .A(n575), .ZN(n540) );
  NAND2_X1 U646 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U647 ( .A(n542), .B(KEYINPUT94), .ZN(n652) );
  OR2_X1 U648 ( .A1(n545), .A2(n544), .ZN(n668) );
  INV_X1 U649 ( .A(n663), .ZN(n665) );
  NAND2_X1 U650 ( .A1(n668), .A2(n665), .ZN(n693) );
  NAND2_X1 U651 ( .A1(KEYINPUT44), .A2(n762), .ZN(n548) );
  NAND2_X1 U652 ( .A1(n550), .A2(KEYINPUT44), .ZN(n551) );
  NOR2_X1 U653 ( .A1(n623), .A2(n399), .ZN(n618) );
  NOR2_X1 U654 ( .A1(G900), .A2(n553), .ZN(n554) );
  NAND2_X1 U655 ( .A1(n554), .A2(G953), .ZN(n555) );
  NAND2_X1 U656 ( .A1(n556), .A2(n555), .ZN(n576) );
  XNOR2_X1 U657 ( .A(KEYINPUT28), .B(n561), .ZN(n563) );
  NAND2_X1 U658 ( .A1(n563), .A2(n562), .ZN(n590) );
  INV_X1 U659 ( .A(n564), .ZN(n565) );
  INV_X1 U660 ( .A(KEYINPUT73), .ZN(n566) );
  NAND2_X1 U661 ( .A1(KEYINPUT47), .A2(n662), .ZN(n567) );
  NAND2_X1 U662 ( .A1(n567), .A2(KEYINPUT73), .ZN(n568) );
  NAND2_X1 U663 ( .A1(n569), .A2(n568), .ZN(n571) );
  AND2_X1 U664 ( .A1(n693), .A2(KEYINPUT73), .ZN(n570) );
  NOR2_X1 U665 ( .A1(n571), .A2(n570), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n679), .A2(n607), .ZN(n574) );
  INV_X1 U667 ( .A(KEYINPUT106), .ZN(n572) );
  XNOR2_X1 U668 ( .A(n572), .B(KEYINPUT30), .ZN(n573) );
  XNOR2_X1 U669 ( .A(n574), .B(n573), .ZN(n579) );
  AND2_X1 U670 ( .A1(n577), .A2(n576), .ZN(n578) );
  AND2_X1 U671 ( .A1(n579), .A2(n578), .ZN(n595) );
  NOR2_X1 U672 ( .A1(n611), .A2(n580), .ZN(n581) );
  NAND2_X1 U673 ( .A1(n595), .A2(n581), .ZN(n582) );
  XNOR2_X1 U674 ( .A(KEYINPUT107), .B(n582), .ZN(n758) );
  XOR2_X1 U675 ( .A(n758), .B(KEYINPUT74), .Z(n583) );
  NAND2_X1 U676 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U677 ( .A1(n586), .A2(n585), .ZN(n603) );
  INV_X1 U678 ( .A(KEYINPUT38), .ZN(n587) );
  NOR2_X1 U679 ( .A1(n689), .A2(n690), .ZN(n588) );
  XNOR2_X1 U680 ( .A(n588), .B(KEYINPUT108), .ZN(n694) );
  NAND2_X1 U681 ( .A1(n694), .A2(n691), .ZN(n589) );
  INV_X1 U682 ( .A(n590), .ZN(n591) );
  INV_X1 U683 ( .A(KEYINPUT109), .ZN(n592) );
  XNOR2_X1 U684 ( .A(n592), .B(KEYINPUT42), .ZN(n593) );
  INV_X1 U685 ( .A(n689), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n595), .A2(n594), .ZN(n598) );
  INV_X1 U687 ( .A(KEYINPUT81), .ZN(n596) );
  XNOR2_X1 U688 ( .A(n596), .B(KEYINPUT39), .ZN(n597) );
  XNOR2_X1 U689 ( .A(n598), .B(n597), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n616), .A2(n663), .ZN(n599) );
  XNOR2_X1 U691 ( .A(n601), .B(n600), .ZN(n602) );
  NAND2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U693 ( .A(KEYINPUT48), .ZN(n604) );
  NAND2_X1 U694 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U695 ( .A(KEYINPUT103), .B(n608), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n609), .A2(n673), .ZN(n610) );
  XNOR2_X1 U697 ( .A(n610), .B(KEYINPUT43), .ZN(n612) );
  AND2_X1 U698 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U699 ( .A(n613), .B(KEYINPUT104), .ZN(n763) );
  INV_X1 U700 ( .A(n763), .ZN(n614) );
  INV_X1 U701 ( .A(n668), .ZN(n659) );
  AND2_X1 U702 ( .A1(n616), .A2(n659), .ZN(n641) );
  INV_X1 U703 ( .A(n641), .ZN(n617) );
  XNOR2_X2 U704 ( .A(n624), .B(KEYINPUT77), .ZN(n751) );
  NAND2_X1 U705 ( .A1(n618), .A2(n751), .ZN(n622) );
  XNOR2_X1 U706 ( .A(n619), .B(KEYINPUT76), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n620), .A2(KEYINPUT2), .ZN(n621) );
  NAND2_X2 U708 ( .A1(n622), .A2(n621), .ZN(n627) );
  INV_X1 U709 ( .A(KEYINPUT2), .ZN(n625) );
  XOR2_X1 U710 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n628) );
  XNOR2_X1 U711 ( .A(n630), .B(n362), .ZN(n632) );
  INV_X1 U712 ( .A(G952), .ZN(n631) );
  AND2_X1 U713 ( .A1(n631), .A2(G953), .ZN(n726) );
  XOR2_X1 U714 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n633) );
  XNOR2_X1 U715 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U718 ( .A(G134), .B(KEYINPUT116), .ZN(n642) );
  XOR2_X1 U719 ( .A(n642), .B(n641), .Z(G36) );
  XNOR2_X1 U720 ( .A(n643), .B(G131), .ZN(G33) );
  XNOR2_X1 U721 ( .A(n644), .B(G101), .ZN(G3) );
  XNOR2_X1 U722 ( .A(n645), .B(KEYINPUT59), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U724 ( .A1(n648), .A2(n726), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n649) );
  XNOR2_X1 U726 ( .A(n650), .B(n649), .ZN(G60) );
  NOR2_X1 U727 ( .A1(n652), .A2(n665), .ZN(n651) );
  XOR2_X1 U728 ( .A(G104), .B(n651), .Z(G6) );
  NOR2_X1 U729 ( .A1(n668), .A2(n652), .ZN(n656) );
  XOR2_X1 U730 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n654) );
  XNOR2_X1 U731 ( .A(G107), .B(KEYINPUT113), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(G9) );
  XNOR2_X1 U734 ( .A(G110), .B(KEYINPUT114), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(n657), .ZN(G12) );
  XOR2_X1 U736 ( .A(G128), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U737 ( .A1(n662), .A2(n659), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n661), .B(n660), .ZN(G30) );
  NAND2_X1 U739 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U740 ( .A(G146), .B(n664), .ZN(G48) );
  NOR2_X1 U741 ( .A1(n665), .A2(n667), .ZN(n666) );
  XOR2_X1 U742 ( .A(G113), .B(n666), .Z(G15) );
  NOR2_X1 U743 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U744 ( .A(G116), .B(n669), .Z(G18) );
  INV_X1 U745 ( .A(n687), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n670), .A2(n688), .ZN(n671) );
  NOR2_X1 U747 ( .A1(G953), .A2(n671), .ZN(n706) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n674), .B(KEYINPUT50), .ZN(n682) );
  XNOR2_X1 U750 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U752 ( .A(n678), .B(n677), .Z(n680) );
  NOR2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U756 ( .A(KEYINPUT51), .B(n685), .Z(n686) );
  NAND2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n700) );
  INV_X1 U758 ( .A(n688), .ZN(n698) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U765 ( .A(KEYINPUT52), .B(n701), .Z(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U767 ( .A(KEYINPUT118), .B(n704), .Z(n705) );
  NAND2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n715) );
  XOR2_X1 U769 ( .A(KEYINPUT2), .B(KEYINPUT72), .Z(n709) );
  INV_X1 U770 ( .A(n707), .ZN(n733) );
  NAND2_X1 U771 ( .A1(n709), .A2(n733), .ZN(n708) );
  XNOR2_X1 U772 ( .A(KEYINPUT75), .B(n708), .ZN(n713) );
  INV_X1 U773 ( .A(n751), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U777 ( .A(KEYINPUT53), .B(n716), .ZN(G75) );
  XOR2_X1 U778 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n718) );
  XNOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n726), .A2(n722), .ZN(G54) );
  XNOR2_X1 U781 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(G63) );
  XOR2_X1 U783 ( .A(n727), .B(KEYINPUT125), .Z(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U785 ( .A(G101), .B(n730), .ZN(n732) );
  NAND2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n740) );
  XOR2_X1 U787 ( .A(KEYINPUT124), .B(n734), .Z(n738) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n735) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n735), .ZN(n736) );
  NAND2_X1 U790 ( .A1(n736), .A2(G898), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U792 ( .A(n740), .B(n739), .Z(G69) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(n747) );
  XNOR2_X1 U794 ( .A(n743), .B(KEYINPUT88), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n752) );
  XNOR2_X1 U797 ( .A(G227), .B(n752), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n749), .A2(G953), .ZN(n750) );
  XNOR2_X1 U800 ( .A(n750), .B(KEYINPUT126), .ZN(n756) );
  XOR2_X1 U801 ( .A(n752), .B(n751), .Z(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(G72) );
  XNOR2_X1 U804 ( .A(n757), .B(G119), .ZN(G21) );
  XOR2_X1 U805 ( .A(G143), .B(n758), .Z(G45) );
  XOR2_X1 U806 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n761) );
  XNOR2_X1 U807 ( .A(G125), .B(n759), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(G27) );
  XOR2_X1 U809 ( .A(n762), .B(G122), .Z(G24) );
  XOR2_X1 U810 ( .A(G140), .B(n763), .Z(G42) );
  XNOR2_X1 U811 ( .A(G137), .B(n764), .ZN(G39) );
endmodule

