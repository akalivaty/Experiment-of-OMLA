

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U323 ( .A1(n371), .A2(n370), .ZN(n372) );
  XOR2_X1 U324 ( .A(n339), .B(n338), .Z(n291) );
  NOR2_X1 U325 ( .A1(n575), .A2(n569), .ZN(n365) );
  XNOR2_X1 U326 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n329) );
  XNOR2_X1 U327 ( .A(n330), .B(n329), .ZN(n363) );
  INV_X1 U328 ( .A(KEYINPUT81), .ZN(n431) );
  XNOR2_X1 U329 ( .A(n389), .B(n388), .ZN(n411) );
  XNOR2_X1 U330 ( .A(n432), .B(n431), .ZN(n433) );
  NOR2_X1 U331 ( .A1(n411), .A2(n514), .ZN(n449) );
  XNOR2_X1 U332 ( .A(n434), .B(n433), .ZN(n435) );
  AND2_X1 U333 ( .A1(n550), .A2(n449), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U335 ( .A(n310), .B(n309), .ZN(n542) );
  XOR2_X1 U336 ( .A(n344), .B(n343), .Z(n581) );
  INV_X1 U337 ( .A(G190GAT), .ZN(n443) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n474) );
  XNOR2_X1 U339 ( .A(n441), .B(n440), .ZN(n527) );
  XNOR2_X1 U340 ( .A(n453), .B(KEYINPUT126), .ZN(n454) );
  XNOR2_X1 U341 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U342 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U343 ( .A(n455), .B(n454), .ZN(G1355GAT) );
  XNOR2_X1 U344 ( .A(n446), .B(n445), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT9), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n292), .B(KEYINPUT7), .ZN(n351) );
  XNOR2_X1 U349 ( .A(n351), .B(G218GAT), .ZN(n293) );
  NAND2_X1 U350 ( .A1(n294), .A2(n293), .ZN(n296) );
  OR2_X1 U351 ( .A1(n294), .A2(n293), .ZN(n295) );
  NAND2_X1 U352 ( .A1(n296), .A2(n295), .ZN(n300) );
  XOR2_X1 U353 ( .A(G36GAT), .B(G92GAT), .Z(n298) );
  NAND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XOR2_X1 U355 ( .A(n298), .B(n297), .Z(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n310) );
  XOR2_X1 U357 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n302) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G162GAT), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U360 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n304) );
  XNOR2_X1 U361 ( .A(G190GAT), .B(G99GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U363 ( .A(n306), .B(n305), .Z(n308) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(G50GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(G134GAT), .B(n542), .ZN(n561) );
  XOR2_X1 U366 ( .A(G57GAT), .B(G78GAT), .Z(n312) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U369 ( .A(KEYINPUT13), .B(G64GAT), .Z(n314) );
  XNOR2_X1 U370 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n328) );
  XOR2_X1 U373 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n318) );
  XNOR2_X1 U374 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n326) );
  NAND2_X1 U376 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XOR2_X1 U377 ( .A(G155GAT), .B(G71GAT), .Z(n320) );
  XNOR2_X1 U378 ( .A(G22GAT), .B(G127GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G183GAT), .Z(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n558) );
  XOR2_X1 U385 ( .A(KEYINPUT36), .B(n561), .Z(n471) );
  NAND2_X1 U386 ( .A1(n558), .A2(n471), .ZN(n330) );
  XOR2_X1 U387 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n332) );
  XNOR2_X1 U388 ( .A(G176GAT), .B(KEYINPUT33), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n344) );
  XNOR2_X1 U390 ( .A(G204GAT), .B(G92GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n333), .B(G64GAT), .ZN(n377) );
  XOR2_X1 U392 ( .A(G85GAT), .B(G57GAT), .Z(n400) );
  XOR2_X1 U393 ( .A(n377), .B(n400), .Z(n335) );
  NAND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n337) );
  XNOR2_X1 U397 ( .A(KEYINPUT13), .B(KEYINPUT74), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G71GAT), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n340), .B(G120GAT), .ZN(n434) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n341), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U403 ( .A(n434), .B(n419), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n291), .B(n342), .ZN(n343) );
  XOR2_X1 U405 ( .A(G36GAT), .B(G8GAT), .Z(n373) );
  XOR2_X1 U406 ( .A(KEYINPUT67), .B(G1GAT), .Z(n346) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G197GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U409 ( .A(n373), .B(n347), .Z(n349) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U412 ( .A(n350), .B(KEYINPUT68), .Z(n353) );
  XNOR2_X1 U413 ( .A(n351), .B(KEYINPUT66), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U415 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n355) );
  XNOR2_X1 U416 ( .A(KEYINPUT30), .B(KEYINPUT70), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U418 ( .A(n357), .B(n356), .Z(n361) );
  XNOR2_X1 U419 ( .A(G43GAT), .B(G15GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n358), .B(G113GAT), .ZN(n437) );
  XNOR2_X1 U421 ( .A(G50GAT), .B(G22GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n359), .B(G141GAT), .ZN(n420) );
  XNOR2_X1 U423 ( .A(n437), .B(n420), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n575) );
  XOR2_X1 U425 ( .A(n575), .B(KEYINPUT71), .Z(n564) );
  AND2_X1 U426 ( .A1(n581), .A2(n564), .ZN(n362) );
  AND2_X1 U427 ( .A1(n363), .A2(n362), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n364), .B(KEYINPUT110), .ZN(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n369) );
  XNOR2_X1 U430 ( .A(KEYINPUT41), .B(n581), .ZN(n533) );
  INV_X1 U431 ( .A(n533), .ZN(n569) );
  XNOR2_X1 U432 ( .A(n365), .B(KEYINPUT46), .ZN(n366) );
  NOR2_X1 U433 ( .A1(n558), .A2(n366), .ZN(n367) );
  NAND2_X1 U434 ( .A1(n367), .A2(n561), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U436 ( .A(KEYINPUT48), .B(n372), .ZN(n549) );
  XOR2_X1 U437 ( .A(KEYINPUT77), .B(n373), .Z(n375) );
  NAND2_X1 U438 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n379) );
  XNOR2_X1 U442 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U444 ( .A(n380), .B(G183GAT), .Z(n382) );
  XNOR2_X1 U445 ( .A(G169GAT), .B(G176GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n430) );
  XOR2_X1 U447 ( .A(G211GAT), .B(KEYINPUT21), .Z(n384) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(G218GAT), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n424) );
  XNOR2_X1 U450 ( .A(n430), .B(n424), .ZN(n385) );
  XOR2_X1 U451 ( .A(n386), .B(n385), .Z(n516) );
  XNOR2_X1 U452 ( .A(KEYINPUT117), .B(n516), .ZN(n387) );
  NOR2_X1 U453 ( .A1(n549), .A2(n387), .ZN(n389) );
  INV_X1 U454 ( .A(KEYINPUT54), .ZN(n388) );
  XOR2_X1 U455 ( .A(G120GAT), .B(G29GAT), .Z(n391) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(G141GAT), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n393) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(G148GAT), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U461 ( .A(n395), .B(n394), .Z(n406) );
  XOR2_X1 U462 ( .A(KEYINPUT87), .B(KEYINPUT1), .Z(n397) );
  XNOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n404) );
  XOR2_X1 U465 ( .A(G155GAT), .B(KEYINPUT3), .Z(n399) );
  XNOR2_X1 U466 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n412) );
  XOR2_X1 U468 ( .A(n412), .B(n400), .Z(n402) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U473 ( .A(n407), .B(KEYINPUT86), .Z(n410) );
  XNOR2_X1 U474 ( .A(G134GAT), .B(G127GAT), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n408), .B(KEYINPUT0), .ZN(n436) );
  XNOR2_X1 U476 ( .A(n436), .B(KEYINPUT88), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n514) );
  XOR2_X1 U478 ( .A(G204GAT), .B(n412), .Z(n414) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n416) );
  XNOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n415) );
  XOR2_X1 U483 ( .A(n416), .B(n415), .Z(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n464) );
  NAND2_X1 U488 ( .A1(n449), .A2(n464), .ZN(n426) );
  XNOR2_X1 U489 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n442) );
  XOR2_X1 U491 ( .A(KEYINPUT80), .B(KEYINPUT64), .Z(n428) );
  XNOR2_X1 U492 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n441) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XOR2_X1 U496 ( .A(n435), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U499 ( .A1(n442), .A2(n527), .ZN(n563) );
  NOR2_X1 U500 ( .A1(n561), .A2(n563), .ZN(n446) );
  XNOR2_X1 U501 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n444) );
  INV_X1 U502 ( .A(KEYINPUT123), .ZN(n451) );
  NOR2_X1 U503 ( .A1(n527), .A2(n464), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT91), .B(n447), .Z(n448) );
  XNOR2_X1 U505 ( .A(KEYINPUT26), .B(n448), .ZN(n550) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n574) );
  NAND2_X1 U507 ( .A1(n574), .A2(n471), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT127), .ZN(n455) );
  XOR2_X1 U509 ( .A(G218GAT), .B(KEYINPUT62), .Z(n453) );
  XNOR2_X1 U510 ( .A(n516), .B(KEYINPUT27), .ZN(n465) );
  NAND2_X1 U511 ( .A1(n465), .A2(n550), .ZN(n460) );
  NAND2_X1 U512 ( .A1(n527), .A2(n516), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n456), .A2(n464), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n457), .Z(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT92), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n461), .B(KEYINPUT93), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n514), .A2(n462), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT94), .ZN(n469) );
  XOR2_X1 U520 ( .A(n464), .B(KEYINPUT28), .Z(n521) );
  NAND2_X1 U521 ( .A1(n514), .A2(n465), .ZN(n548) );
  NOR2_X1 U522 ( .A1(n521), .A2(n548), .ZN(n530) );
  XOR2_X1 U523 ( .A(n527), .B(KEYINPUT84), .Z(n466) );
  NAND2_X1 U524 ( .A1(n530), .A2(n466), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT90), .B(n467), .Z(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n480) );
  NOR2_X1 U527 ( .A1(n558), .A2(n480), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT37), .B(n472), .Z(n513) );
  INV_X1 U530 ( .A(n564), .ZN(n531) );
  NAND2_X1 U531 ( .A1(n531), .A2(n581), .ZN(n483) );
  OR2_X1 U532 ( .A1(n513), .A2(n483), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT38), .B(n473), .Z(n498) );
  NAND2_X1 U534 ( .A1(n527), .A2(n498), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n479) );
  NAND2_X1 U537 ( .A1(n561), .A2(n558), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(KEYINPUT95), .ZN(n501) );
  NOR2_X1 U541 ( .A1(n483), .A2(n501), .ZN(n491) );
  NAND2_X1 U542 ( .A1(n514), .A2(n491), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n516), .A2(n491), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT96), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT35), .B(KEYINPUT97), .Z(n489) );
  NAND2_X1 U549 ( .A1(n491), .A2(n527), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NAND2_X1 U552 ( .A1(n491), .A2(n521), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n498), .A2(n514), .ZN(n495) );
  XOR2_X1 U558 ( .A(n496), .B(n495), .Z(G1328GAT) );
  NAND2_X1 U559 ( .A1(n498), .A2(n516), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT101), .Z(n500) );
  NAND2_X1 U562 ( .A1(n521), .A2(n498), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  NAND2_X1 U564 ( .A1(n575), .A2(n533), .ZN(n512) );
  NOR2_X1 U565 ( .A1(n512), .A2(n501), .ZN(n502) );
  XNOR2_X1 U566 ( .A(KEYINPUT102), .B(n502), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n508), .A2(n514), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n516), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U572 ( .A(G71GAT), .B(KEYINPUT103), .Z(n507) );
  NAND2_X1 U573 ( .A1(n527), .A2(n508), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n510) );
  NAND2_X1 U576 ( .A1(n521), .A2(n508), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n514), .A2(n522), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n522), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n519) );
  NAND2_X1 U585 ( .A1(n522), .A2(n527), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n520), .ZN(G1338GAT) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n526) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n524) );
  NAND2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  INV_X1 U593 ( .A(n527), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n528), .A2(n549), .ZN(n529) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n544) );
  INV_X1 U596 ( .A(n544), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n531), .A2(n543), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G113GAT), .ZN(G1340GAT) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n535) );
  NAND2_X1 U601 ( .A1(n543), .A2(n533), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT111), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n540) );
  NAND2_X1 U606 ( .A1(n543), .A2(n558), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U610 ( .A1(G134GAT), .A2(n544), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n560) );
  NOR2_X1 U615 ( .A1(n575), .A2(n560), .ZN(n553) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n555) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n569), .A2(n560), .ZN(n556) );
  XOR2_X1 U622 ( .A(n557), .B(n556), .Z(G1345GAT) );
  INV_X1 U623 ( .A(n558), .ZN(n585) );
  NOR2_X1 U624 ( .A1(n585), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n568) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n571) );
  NOR2_X1 U634 ( .A1(n569), .A2(n563), .ZN(n570) );
  XOR2_X1 U635 ( .A(n571), .B(n570), .Z(G1349GAT) );
  NOR2_X1 U636 ( .A1(n585), .A2(n563), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  INV_X1 U639 ( .A(n574), .ZN(n584) );
  NOR2_X1 U640 ( .A1(n575), .A2(n584), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
endmodule

