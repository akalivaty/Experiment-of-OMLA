

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733;

  INV_X1 U363 ( .A(n348), .ZN(n672) );
  XNOR2_X1 U364 ( .A(n718), .B(n456), .ZN(n485) );
  NAND2_X1 U365 ( .A1(n678), .A2(n395), .ZN(n348) );
  XNOR2_X2 U366 ( .A(n400), .B(G134), .ZN(n454) );
  NAND2_X1 U367 ( .A1(n729), .A2(n733), .ZN(n542) );
  XOR2_X1 U368 ( .A(n466), .B(KEYINPUT23), .Z(n343) );
  INV_X2 U369 ( .A(G953), .ZN(n720) );
  INV_X1 U370 ( .A(G472), .ZN(n463) );
  AND2_X1 U371 ( .A1(n719), .A2(n382), .ZN(n351) );
  NAND2_X1 U372 ( .A1(n406), .A2(n544), .ZN(n595) );
  NOR2_X1 U373 ( .A1(n731), .A2(n730), .ZN(n583) );
  XNOR2_X1 U374 ( .A(n513), .B(KEYINPUT35), .ZN(n728) );
  XNOR2_X1 U375 ( .A(n418), .B(n417), .ZN(n730) );
  AND2_X1 U376 ( .A1(n409), .A2(n408), .ZN(n632) );
  XNOR2_X1 U377 ( .A(n398), .B(n533), .ZN(n629) );
  XNOR2_X1 U378 ( .A(n506), .B(n345), .ZN(n378) );
  XOR2_X1 U379 ( .A(n694), .B(KEYINPUT123), .Z(n696) );
  XNOR2_X1 U380 ( .A(n709), .B(n396), .ZN(n499) );
  XNOR2_X1 U381 ( .A(n489), .B(G104), .ZN(n709) );
  XNOR2_X1 U382 ( .A(n458), .B(n457), .ZN(n503) );
  BUF_X1 U383 ( .A(n699), .Z(n344) );
  AND2_X2 U384 ( .A1(n348), .A2(n599), .ZN(n699) );
  XNOR2_X2 U385 ( .A(n454), .B(n366), .ZN(n718) );
  NOR2_X1 U386 ( .A1(n600), .A2(G902), .ZN(n465) );
  XNOR2_X1 U387 ( .A(n397), .B(n499), .ZN(n606) );
  XNOR2_X1 U388 ( .A(n500), .B(n504), .ZN(n397) );
  XNOR2_X1 U389 ( .A(n386), .B(n498), .ZN(n500) );
  NOR2_X1 U390 ( .A1(n404), .A2(n403), .ZN(n402) );
  INV_X1 U391 ( .A(n634), .ZN(n403) );
  XNOR2_X1 U392 ( .A(n595), .B(KEYINPUT45), .ZN(n405) );
  NAND2_X1 U393 ( .A1(n514), .A2(n528), .ZN(n564) );
  XNOR2_X1 U394 ( .A(KEYINPUT105), .B(n520), .ZN(n522) );
  XNOR2_X1 U395 ( .A(n425), .B(G131), .ZN(n455) );
  INV_X1 U396 ( .A(KEYINPUT69), .ZN(n425) );
  XNOR2_X1 U397 ( .A(n728), .B(n389), .ZN(n526) );
  INV_X1 U398 ( .A(KEYINPUT44), .ZN(n389) );
  XNOR2_X1 U399 ( .A(n459), .B(n350), .ZN(n349) );
  INV_X1 U400 ( .A(G101), .ZN(n350) );
  NOR2_X1 U401 ( .A1(G953), .A2(G237), .ZN(n461) );
  XNOR2_X1 U402 ( .A(G119), .B(KEYINPUT3), .ZN(n457) );
  XOR2_X1 U403 ( .A(G113), .B(G116), .Z(n458) );
  XOR2_X1 U404 ( .A(G146), .B(G125), .Z(n497) );
  XOR2_X1 U405 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n443) );
  XNOR2_X1 U406 ( .A(G143), .B(G113), .ZN(n439) );
  XOR2_X1 U407 ( .A(G122), .B(G104), .Z(n440) );
  XNOR2_X1 U408 ( .A(n455), .B(n367), .ZN(n366) );
  XNOR2_X1 U409 ( .A(n424), .B(n368), .ZN(n367) );
  INV_X1 U410 ( .A(KEYINPUT4), .ZN(n424) );
  NOR2_X1 U411 ( .A1(n553), .A2(n627), .ZN(n586) );
  XNOR2_X1 U412 ( .A(n497), .B(n360), .ZN(n717) );
  XNOR2_X1 U413 ( .A(KEYINPUT10), .B(G140), .ZN(n360) );
  XNOR2_X1 U414 ( .A(G119), .B(G110), .ZN(n466) );
  XNOR2_X1 U415 ( .A(G137), .B(G128), .ZN(n467) );
  XNOR2_X1 U416 ( .A(n450), .B(n393), .ZN(n392) );
  INV_X1 U417 ( .A(KEYINPUT7), .ZN(n393) );
  XOR2_X1 U418 ( .A(G122), .B(KEYINPUT9), .Z(n450) );
  XNOR2_X1 U419 ( .A(G116), .B(G107), .ZN(n451) );
  XNOR2_X1 U420 ( .A(n449), .B(n355), .ZN(n470) );
  INV_X1 U421 ( .A(KEYINPUT8), .ZN(n355) );
  INV_X1 U422 ( .A(KEYINPUT71), .ZN(n396) );
  INV_X1 U423 ( .A(G146), .ZN(n456) );
  INV_X1 U424 ( .A(KEYINPUT39), .ZN(n423) );
  XNOR2_X1 U425 ( .A(n586), .B(KEYINPUT112), .ZN(n413) );
  INV_X1 U426 ( .A(n587), .ZN(n412) );
  INV_X1 U427 ( .A(n522), .ZN(n375) );
  INV_X1 U428 ( .A(n538), .ZN(n372) );
  NAND2_X1 U429 ( .A1(n358), .A2(n357), .ZN(n362) );
  INV_X1 U430 ( .A(n564), .ZN(n358) );
  INV_X1 U431 ( .A(n563), .ZN(n357) );
  XNOR2_X1 U432 ( .A(n453), .B(G478), .ZN(n529) );
  XNOR2_X1 U433 ( .A(n447), .B(n448), .ZN(n528) );
  XNOR2_X1 U434 ( .A(n587), .B(n508), .ZN(n573) );
  XNOR2_X1 U435 ( .A(n516), .B(n515), .ZN(n521) );
  XNOR2_X1 U436 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n515) );
  XNOR2_X1 U437 ( .A(n391), .B(n390), .ZN(n430) );
  INV_X1 U438 ( .A(n588), .ZN(n408) );
  NAND2_X1 U439 ( .A1(n521), .A2(n401), .ZN(n538) );
  NAND2_X1 U440 ( .A1(n381), .A2(n347), .ZN(n599) );
  INV_X1 U441 ( .A(G137), .ZN(n368) );
  XNOR2_X1 U442 ( .A(n400), .B(n432), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n434), .B(n433), .ZN(n432) );
  XNOR2_X1 U444 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n434) );
  NAND2_X1 U445 ( .A1(n720), .A2(G224), .ZN(n433) );
  INV_X1 U446 ( .A(KEYINPUT64), .ZN(n428) );
  OR2_X1 U447 ( .A1(G237), .A2(G902), .ZN(n507) );
  XOR2_X1 U448 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n474) );
  XNOR2_X2 U449 ( .A(G110), .B(KEYINPUT86), .ZN(n486) );
  XNOR2_X1 U450 ( .A(G902), .B(KEYINPUT15), .ZN(n593) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n493) );
  XNOR2_X1 U452 ( .A(n352), .B(KEYINPUT102), .ZN(n657) );
  NOR2_X1 U453 ( .A1(n657), .A2(n641), .ZN(n391) );
  INV_X1 U454 ( .A(KEYINPUT103), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n485), .B(n414), .ZN(n600) );
  XNOR2_X1 U456 ( .A(n503), .B(n349), .ZN(n460) );
  XNOR2_X1 U457 ( .A(n595), .B(KEYINPUT45), .ZN(n395) );
  INV_X1 U458 ( .A(KEYINPUT16), .ZN(n501) );
  XNOR2_X1 U459 ( .A(n446), .B(n359), .ZN(n688) );
  XNOR2_X1 U460 ( .A(n441), .B(n717), .ZN(n359) );
  XNOR2_X1 U461 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n431) );
  XNOR2_X1 U462 ( .A(n600), .B(KEYINPUT62), .ZN(n601) );
  AND2_X1 U463 ( .A1(n395), .A2(n720), .ZN(n707) );
  XNOR2_X1 U464 ( .A(n471), .B(n388), .ZN(n472) );
  XNOR2_X1 U465 ( .A(n469), .B(n343), .ZN(n388) );
  XNOR2_X1 U466 ( .A(n356), .B(n354), .ZN(n452) );
  NAND2_X1 U467 ( .A1(n470), .A2(G217), .ZN(n354) );
  XNOR2_X1 U468 ( .A(n392), .B(n451), .ZN(n356) );
  XNOR2_X1 U469 ( .A(n485), .B(n426), .ZN(n684) );
  XNOR2_X1 U470 ( .A(n499), .B(n484), .ZN(n426) );
  XNOR2_X1 U471 ( .A(n608), .B(n607), .ZN(n610) );
  NOR2_X1 U472 ( .A1(G952), .A2(n720), .ZN(n703) );
  XNOR2_X1 U473 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n417) );
  NAND2_X1 U474 ( .A1(n420), .A2(n419), .ZN(n418) );
  INV_X1 U475 ( .A(n582), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n731) );
  INV_X1 U477 ( .A(KEYINPUT40), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n409) );
  INV_X1 U479 ( .A(KEYINPUT36), .ZN(n410) );
  NOR2_X1 U480 ( .A1(n380), .A2(n564), .ZN(n513) );
  XNOR2_X1 U481 ( .A(n512), .B(n511), .ZN(n380) );
  NAND2_X1 U482 ( .A1(n373), .A2(n370), .ZN(n729) );
  NAND2_X1 U483 ( .A1(n372), .A2(n346), .ZN(n370) );
  AND2_X1 U484 ( .A1(n376), .A2(n374), .ZN(n373) );
  INV_X1 U485 ( .A(KEYINPUT110), .ZN(n384) );
  NOR2_X2 U486 ( .A1(n573), .A2(n582), .ZN(n625) );
  NOR2_X1 U487 ( .A1(n369), .A2(n394), .ZN(n679) );
  XNOR2_X1 U488 ( .A(n505), .B(KEYINPUT87), .ZN(n345) );
  AND2_X1 U489 ( .A1(n522), .A2(n371), .ZN(n346) );
  XNOR2_X1 U490 ( .A(KEYINPUT66), .B(n594), .ZN(n347) );
  INV_X1 U491 ( .A(n562), .ZN(n363) );
  XNOR2_X1 U492 ( .A(n558), .B(KEYINPUT30), .ZN(n562) );
  NAND2_X1 U493 ( .A1(n405), .A2(n719), .ZN(n369) );
  NAND2_X1 U494 ( .A1(n351), .A2(n405), .ZN(n381) );
  INV_X1 U495 ( .A(n529), .ZN(n514) );
  NAND2_X1 U496 ( .A1(n529), .A2(n353), .ZN(n352) );
  INV_X1 U497 ( .A(n528), .ZN(n353) );
  NAND2_X1 U498 ( .A1(n363), .A2(n361), .ZN(n385) );
  NOR2_X1 U499 ( .A1(n415), .A2(n362), .ZN(n361) );
  NOR2_X1 U500 ( .A1(n562), .A2(n415), .ZN(n364) );
  AND2_X1 U501 ( .A1(n364), .A2(n655), .ZN(n580) );
  NAND2_X1 U502 ( .A1(n365), .A2(n638), .ZN(n416) );
  XNOR2_X1 U503 ( .A(n365), .B(KEYINPUT1), .ZN(n637) );
  NAND2_X1 U504 ( .A1(n572), .A2(n365), .ZN(n582) );
  XNOR2_X2 U505 ( .A(n490), .B(G469), .ZN(n365) );
  XNOR2_X2 U506 ( .A(n435), .B(G143), .ZN(n400) );
  NAND2_X1 U507 ( .A1(n538), .A2(n523), .ZN(n376) );
  INV_X1 U508 ( .A(n523), .ZN(n371) );
  NAND2_X1 U509 ( .A1(n375), .A2(n523), .ZN(n374) );
  NAND2_X1 U510 ( .A1(n378), .A2(n654), .ZN(n587) );
  INV_X1 U511 ( .A(n378), .ZN(n563) );
  XNOR2_X1 U512 ( .A(n563), .B(KEYINPUT38), .ZN(n655) );
  OR2_X1 U513 ( .A1(n557), .A2(n378), .ZN(n377) );
  XNOR2_X1 U514 ( .A(n609), .B(n610), .ZN(n611) );
  XNOR2_X1 U515 ( .A(n695), .B(n696), .ZN(n697) );
  INV_X1 U516 ( .A(n677), .ZN(n678) );
  NAND2_X1 U517 ( .A1(n597), .A2(n598), .ZN(n677) );
  NAND2_X1 U518 ( .A1(n379), .A2(n526), .ZN(n544) );
  NAND2_X1 U519 ( .A1(n525), .A2(n728), .ZN(n379) );
  NAND2_X1 U520 ( .A1(n542), .A2(KEYINPUT44), .ZN(n429) );
  INV_X1 U521 ( .A(n593), .ZN(n382) );
  XNOR2_X1 U522 ( .A(n429), .B(n428), .ZN(n427) );
  NOR2_X1 U523 ( .A1(n401), .A2(n570), .ZN(n552) );
  NAND2_X1 U524 ( .A1(n413), .A2(n412), .ZN(n411) );
  NOR2_X2 U525 ( .A1(n603), .A2(n703), .ZN(n605) );
  NOR2_X2 U526 ( .A1(n697), .A2(n703), .ZN(n698) );
  NOR2_X2 U527 ( .A1(n691), .A2(n703), .ZN(n693) );
  INV_X1 U528 ( .A(n653), .ZN(n420) );
  NAND2_X1 U529 ( .A1(n655), .A2(n654), .ZN(n658) );
  XNOR2_X1 U530 ( .A(n383), .B(n613), .ZN(G51) );
  NOR2_X2 U531 ( .A1(n611), .A2(n703), .ZN(n383) );
  XNOR2_X2 U532 ( .A(n385), .B(n384), .ZN(n732) );
  NAND2_X1 U533 ( .A1(n387), .A2(n566), .ZN(n568) );
  XNOR2_X1 U534 ( .A(n732), .B(KEYINPUT81), .ZN(n387) );
  NOR2_X2 U535 ( .A1(n590), .A2(n589), .ZN(n591) );
  AND2_X2 U536 ( .A1(n407), .A2(n402), .ZN(n719) );
  XNOR2_X1 U537 ( .A(n460), .B(n462), .ZN(n414) );
  NOR2_X1 U538 ( .A1(n427), .A2(n543), .ZN(n406) );
  XNOR2_X2 U539 ( .A(n479), .B(n478), .ZN(n642) );
  INV_X1 U540 ( .A(n677), .ZN(n394) );
  NOR2_X1 U541 ( .A1(n694), .A2(G902), .ZN(n453) );
  NAND2_X1 U542 ( .A1(n535), .A2(n649), .ZN(n398) );
  XNOR2_X2 U543 ( .A(n399), .B(n431), .ZN(n535) );
  NOR2_X2 U544 ( .A1(n573), .A2(n509), .ZN(n399) );
  NOR2_X1 U545 ( .A1(n401), .A2(n532), .ZN(n492) );
  XNOR2_X2 U546 ( .A(n647), .B(KEYINPUT6), .ZN(n401) );
  AND2_X1 U547 ( .A1(n407), .A2(n377), .ZN(n597) );
  INV_X1 U548 ( .A(n377), .ZN(n404) );
  XNOR2_X1 U549 ( .A(n591), .B(KEYINPUT48), .ZN(n407) );
  NAND2_X1 U550 ( .A1(n535), .A2(n430), .ZN(n516) );
  NAND2_X1 U551 ( .A1(n561), .A2(n560), .ZN(n415) );
  XNOR2_X2 U552 ( .A(n416), .B(KEYINPUT93), .ZN(n561) );
  NAND2_X1 U553 ( .A1(n592), .A2(n624), .ZN(n422) );
  XNOR2_X1 U554 ( .A(n580), .B(n423), .ZN(n592) );
  XNOR2_X2 U555 ( .A(G128), .B(KEYINPUT78), .ZN(n435) );
  INV_X2 U556 ( .A(n569), .ZN(n647) );
  XNOR2_X1 U557 ( .A(n542), .B(n524), .ZN(n525) );
  OR2_X2 U558 ( .A1(n684), .A2(G902), .ZN(n490) );
  XOR2_X1 U559 ( .A(n683), .B(n682), .Z(n436) );
  OR2_X1 U560 ( .A1(n647), .A2(n517), .ZN(n437) );
  XNOR2_X1 U561 ( .A(KEYINPUT59), .B(KEYINPUT85), .ZN(n438) );
  INV_X1 U562 ( .A(KEYINPUT80), .ZN(n567) );
  XNOR2_X1 U563 ( .A(n568), .B(n567), .ZN(n577) );
  INV_X1 U564 ( .A(KEYINPUT83), .ZN(n524) );
  INV_X1 U565 ( .A(n710), .ZN(n504) );
  INV_X1 U566 ( .A(n642), .ZN(n517) );
  XNOR2_X1 U567 ( .A(n501), .B(G122), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n463), .B(KEYINPUT95), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n688), .B(n438), .ZN(n689) );
  NOR2_X1 U570 ( .A1(n408), .A2(n437), .ZN(n518) );
  XNOR2_X1 U571 ( .A(n690), .B(n689), .ZN(n691) );
  INV_X1 U572 ( .A(KEYINPUT63), .ZN(n604) );
  XNOR2_X1 U573 ( .A(KEYINPUT13), .B(G475), .ZN(n448) );
  XNOR2_X1 U574 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U575 ( .A(n455), .B(KEYINPUT98), .ZN(n445) );
  NAND2_X1 U576 ( .A1(G214), .A2(n461), .ZN(n442) );
  XNOR2_X1 U577 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U578 ( .A(n445), .B(n444), .ZN(n446) );
  NOR2_X1 U579 ( .A1(G902), .A2(n688), .ZN(n447) );
  NAND2_X1 U580 ( .A1(G234), .A2(n720), .ZN(n449) );
  XNOR2_X1 U581 ( .A(n454), .B(n452), .ZN(n694) );
  XOR2_X1 U582 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n459) );
  NAND2_X1 U583 ( .A1(n461), .A2(G210), .ZN(n462) );
  XNOR2_X2 U584 ( .A(n465), .B(n464), .ZN(n569) );
  XOR2_X1 U585 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n468) );
  XNOR2_X1 U586 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U587 ( .A1(G221), .A2(n470), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n472), .B(n717), .ZN(n701) );
  NOR2_X1 U589 ( .A1(G902), .A2(n701), .ZN(n479) );
  XOR2_X1 U590 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n476) );
  NAND2_X1 U591 ( .A1(G234), .A2(n593), .ZN(n473) );
  XNOR2_X1 U592 ( .A(n474), .B(n473), .ZN(n480) );
  NAND2_X1 U593 ( .A1(n480), .A2(G217), .ZN(n475) );
  XNOR2_X1 U594 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U595 ( .A(KEYINPUT90), .B(n477), .ZN(n478) );
  NAND2_X1 U596 ( .A1(n480), .A2(G221), .ZN(n481) );
  XNOR2_X1 U597 ( .A(n481), .B(KEYINPUT21), .ZN(n641) );
  NOR2_X1 U598 ( .A1(n642), .A2(n641), .ZN(n638) );
  XOR2_X1 U599 ( .A(G140), .B(KEYINPUT76), .Z(n483) );
  NAND2_X1 U600 ( .A1(G227), .A2(n720), .ZN(n482) );
  XNOR2_X1 U601 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U602 ( .A(n486), .ZN(n488) );
  XNOR2_X1 U603 ( .A(G101), .B(G107), .ZN(n487) );
  XNOR2_X1 U604 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U605 ( .A1(n638), .A2(n637), .ZN(n532) );
  XNOR2_X1 U606 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n491) );
  XNOR2_X1 U607 ( .A(n492), .B(n491), .ZN(n664) );
  XOR2_X1 U608 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n494) );
  XNOR2_X1 U609 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U610 ( .A1(G952), .A2(n495), .ZN(n670) );
  NOR2_X1 U611 ( .A1(G953), .A2(n670), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G902), .A2(n495), .ZN(n546) );
  XOR2_X1 U613 ( .A(G898), .B(KEYINPUT88), .Z(n706) );
  NAND2_X1 U614 ( .A1(G953), .A2(n706), .ZN(n712) );
  NOR2_X1 U615 ( .A1(n546), .A2(n712), .ZN(n496) );
  NOR2_X1 U616 ( .A1(n549), .A2(n496), .ZN(n509) );
  XNOR2_X1 U617 ( .A(KEYINPUT4), .B(n497), .ZN(n498) );
  XNOR2_X1 U618 ( .A(n503), .B(n502), .ZN(n710) );
  NAND2_X1 U619 ( .A1(n606), .A2(n593), .ZN(n506) );
  NAND2_X1 U620 ( .A1(n507), .A2(G210), .ZN(n505) );
  NAND2_X1 U621 ( .A1(G214), .A2(n507), .ZN(n654) );
  XNOR2_X1 U622 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n508) );
  INV_X1 U623 ( .A(n535), .ZN(n510) );
  NOR2_X1 U624 ( .A1(n664), .A2(n510), .ZN(n512) );
  XNOR2_X1 U625 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n511) );
  INV_X1 U626 ( .A(n637), .ZN(n588) );
  NAND2_X1 U627 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U628 ( .A(n519), .B(KEYINPUT106), .ZN(n733) );
  NAND2_X1 U629 ( .A1(n642), .A2(n408), .ZN(n520) );
  XOR2_X1 U630 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n523) );
  NOR2_X1 U631 ( .A1(n529), .A2(n528), .ZN(n527) );
  XNOR2_X1 U632 ( .A(n527), .B(KEYINPUT100), .ZN(n621) );
  NAND2_X1 U633 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U634 ( .A(n530), .B(KEYINPUT99), .ZN(n624) );
  NOR2_X1 U635 ( .A1(n621), .A2(n624), .ZN(n531) );
  XNOR2_X1 U636 ( .A(n531), .B(KEYINPUT101), .ZN(n565) );
  XOR2_X1 U637 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n533) );
  NOR2_X1 U638 ( .A1(n569), .A2(n532), .ZN(n649) );
  AND2_X1 U639 ( .A1(n561), .A2(n569), .ZN(n534) );
  NAND2_X1 U640 ( .A1(n535), .A2(n534), .ZN(n616) );
  NAND2_X1 U641 ( .A1(n629), .A2(n616), .ZN(n536) );
  XOR2_X1 U642 ( .A(KEYINPUT97), .B(n536), .Z(n537) );
  NAND2_X1 U643 ( .A1(n565), .A2(n537), .ZN(n540) );
  NOR2_X1 U644 ( .A1(n642), .A2(n538), .ZN(n539) );
  NAND2_X1 U645 ( .A1(n588), .A2(n539), .ZN(n614) );
  NAND2_X1 U646 ( .A1(n540), .A2(n614), .ZN(n541) );
  XNOR2_X1 U647 ( .A(n541), .B(KEYINPUT104), .ZN(n543) );
  XOR2_X1 U648 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n545) );
  XNOR2_X1 U649 ( .A(KEYINPUT108), .B(n545), .ZN(n556) );
  OR2_X1 U650 ( .A1(n720), .A2(n546), .ZN(n547) );
  NOR2_X1 U651 ( .A1(G900), .A2(n547), .ZN(n548) );
  NOR2_X1 U652 ( .A1(n549), .A2(n548), .ZN(n559) );
  NOR2_X1 U653 ( .A1(n641), .A2(n559), .ZN(n550) );
  NAND2_X1 U654 ( .A1(n642), .A2(n550), .ZN(n551) );
  XNOR2_X1 U655 ( .A(KEYINPUT70), .B(n551), .ZN(n570) );
  XNOR2_X1 U656 ( .A(n552), .B(KEYINPUT107), .ZN(n553) );
  INV_X1 U657 ( .A(n624), .ZN(n627) );
  NAND2_X1 U658 ( .A1(n586), .A2(n654), .ZN(n554) );
  NOR2_X1 U659 ( .A1(n408), .A2(n554), .ZN(n555) );
  XNOR2_X1 U660 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U661 ( .A1(n647), .A2(n654), .ZN(n558) );
  INV_X1 U662 ( .A(n559), .ZN(n560) );
  INV_X1 U663 ( .A(n565), .ZN(n659) );
  NAND2_X1 U664 ( .A1(n659), .A2(KEYINPUT47), .ZN(n566) );
  NOR2_X1 U665 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U666 ( .A(KEYINPUT28), .B(n571), .ZN(n572) );
  XOR2_X1 U667 ( .A(n625), .B(KEYINPUT47), .Z(n575) );
  NAND2_X1 U668 ( .A1(n625), .A2(n659), .ZN(n574) );
  NAND2_X1 U669 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U670 ( .A1(n577), .A2(n576), .ZN(n579) );
  INV_X1 U671 ( .A(KEYINPUT74), .ZN(n578) );
  XNOR2_X1 U672 ( .A(n579), .B(n578), .ZN(n585) );
  NOR2_X1 U673 ( .A1(n657), .A2(n658), .ZN(n581) );
  XNOR2_X1 U674 ( .A(KEYINPUT41), .B(n581), .ZN(n653) );
  XNOR2_X1 U675 ( .A(n583), .B(KEYINPUT46), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n585), .A2(n584), .ZN(n590) );
  XNOR2_X1 U677 ( .A(n632), .B(KEYINPUT82), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n592), .A2(n621), .ZN(n634) );
  INV_X1 U679 ( .A(KEYINPUT2), .ZN(n671) );
  OR2_X1 U680 ( .A1(n593), .A2(n671), .ZN(n594) );
  NAND2_X1 U681 ( .A1(KEYINPUT2), .A2(n634), .ZN(n596) );
  XNOR2_X1 U682 ( .A(KEYINPUT79), .B(n596), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n699), .A2(G472), .ZN(n602) );
  XNOR2_X1 U684 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U685 ( .A(n605), .B(n604), .ZN(G57) );
  XNOR2_X1 U686 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n606), .B(KEYINPUT84), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n699), .A2(G210), .ZN(n609) );
  INV_X1 U689 ( .A(KEYINPUT119), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT56), .ZN(n613) );
  XNOR2_X1 U691 ( .A(G101), .B(n614), .ZN(G3) );
  NOR2_X1 U692 ( .A1(n627), .A2(n616), .ZN(n615) );
  XOR2_X1 U693 ( .A(G104), .B(n615), .Z(G6) );
  INV_X1 U694 ( .A(n621), .ZN(n630) );
  NOR2_X1 U695 ( .A1(n616), .A2(n630), .ZN(n620) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n618) );
  XNOR2_X1 U697 ( .A(G107), .B(KEYINPUT26), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n620), .B(n619), .ZN(G9) );
  XOR2_X1 U700 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U701 ( .A1(n625), .A2(n621), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n623), .B(n622), .ZN(G30) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(G146), .ZN(G48) );
  NOR2_X1 U705 ( .A1(n629), .A2(n627), .ZN(n628) );
  XOR2_X1 U706 ( .A(G113), .B(n628), .Z(G15) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U708 ( .A(G116), .B(n631), .Z(G18) );
  XNOR2_X1 U709 ( .A(G125), .B(n632), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U711 ( .A(G134), .B(n634), .ZN(G36) );
  XOR2_X1 U712 ( .A(G140), .B(n404), .Z(n635) );
  XNOR2_X1 U713 ( .A(KEYINPUT114), .B(n635), .ZN(G42) );
  NOR2_X1 U714 ( .A1(n664), .A2(n653), .ZN(n636) );
  NOR2_X1 U715 ( .A1(G953), .A2(n636), .ZN(n676) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U717 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n640), .B(n639), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT49), .B(n643), .Z(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U724 ( .A(n650), .B(KEYINPUT51), .Z(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT116), .B(n651), .ZN(n652) );
  NOR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n666) );
  NOR2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U730 ( .A(KEYINPUT117), .B(n660), .Z(n661) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT52), .ZN(n668) );
  XNOR2_X1 U735 ( .A(KEYINPUT118), .B(n668), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n680) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U741 ( .A(n681), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U742 ( .A1(n344), .A2(G469), .ZN(n686) );
  XOR2_X1 U743 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n683) );
  XNOR2_X1 U744 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n684), .B(n436), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U747 ( .A1(n703), .A2(n687), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n699), .A2(G475), .ZN(n690) );
  XNOR2_X1 U749 ( .A(KEYINPUT60), .B(KEYINPUT122), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(G60) );
  NAND2_X1 U751 ( .A1(n699), .A2(G478), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n698), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U753 ( .A1(G217), .A2(n344), .ZN(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(G66) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n704) );
  XOR2_X1 U757 ( .A(KEYINPUT61), .B(n704), .Z(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n708) );
  NOR2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n715) );
  XNOR2_X1 U760 ( .A(KEYINPUT126), .B(n709), .ZN(n711) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U764 ( .A(KEYINPUT125), .B(n716), .Z(G69) );
  XOR2_X1 U765 ( .A(n718), .B(n717), .Z(n722) );
  XNOR2_X1 U766 ( .A(n722), .B(n719), .ZN(n721) );
  NAND2_X1 U767 ( .A1(n721), .A2(n720), .ZN(n727) );
  XNOR2_X1 U768 ( .A(n722), .B(G227), .ZN(n723) );
  XNOR2_X1 U769 ( .A(n723), .B(KEYINPUT127), .ZN(n724) );
  NAND2_X1 U770 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(G953), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n727), .A2(n726), .ZN(G72) );
  XNOR2_X1 U773 ( .A(G122), .B(n728), .ZN(G24) );
  XNOR2_X1 U774 ( .A(n729), .B(G119), .ZN(G21) );
  XOR2_X1 U775 ( .A(G137), .B(n730), .Z(G39) );
  XOR2_X1 U776 ( .A(G131), .B(n731), .Z(G33) );
  XOR2_X1 U777 ( .A(n732), .B(G143), .Z(G45) );
  XNOR2_X1 U778 ( .A(G110), .B(n733), .ZN(G12) );
endmodule

