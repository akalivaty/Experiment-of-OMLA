//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT1), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT66), .Z(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n218));
  AND3_X1   g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n207), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n203), .A2(G50), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n213), .B2(new_n220), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n220), .A2(new_n213), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT67), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n240), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT74), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(new_n249), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G238), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(new_n254), .B2(new_n249), .ZN(new_n258));
  OAI211_X1 g0058(.A(KEYINPUT75), .B(new_n252), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n249), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT74), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G238), .A3(new_n256), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT75), .B1(new_n263), .B2(new_n252), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G97), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(G226), .A4(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n266), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n274), .A2(KEYINPUT73), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT73), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n260), .A2(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n263), .A2(new_n252), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT75), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n259), .ZN(new_n284));
  INV_X1    g0084(.A(new_n277), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n274), .A2(KEYINPUT73), .A3(new_n275), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n280), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G169), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT14), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n284), .A2(new_n287), .A3(new_n280), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n290), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n268), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n241), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n221), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(KEYINPUT11), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n202), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT12), .ZN(new_n312));
  INV_X1    g0112(.A(new_n307), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G1), .B2(new_n300), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n308), .B(new_n312), .C1(new_n202), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT11), .B1(new_n305), .B2(new_n307), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n299), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n297), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n319), .B2(G190), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n324));
  INV_X1    g0124(.A(G150), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n304), .ZN(new_n326));
  OR2_X1    g0126(.A1(KEYINPUT68), .A2(G58), .ZN(new_n327));
  NAND2_X1  g0127(.A1(KEYINPUT68), .A2(G58), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT8), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT69), .B1(new_n201), .B2(KEYINPUT8), .ZN(new_n331));
  OR3_X1    g0131(.A1(new_n201), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n326), .B1(new_n333), .B2(new_n302), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n313), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n310), .A2(new_n241), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n314), .B2(new_n241), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n335), .A2(new_n340), .A3(new_n337), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n338), .A2(KEYINPUT71), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT72), .B(KEYINPUT9), .C1(new_n346), .C2(new_n343), .ZN(new_n347));
  INV_X1    g0147(.A(G226), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n252), .B1(new_n261), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n265), .A2(G222), .A3(new_n272), .ZN(new_n350));
  INV_X1    g0150(.A(G77), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n265), .A2(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G223), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n350), .B1(new_n351), .B2(new_n265), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n354), .B2(new_n275), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n321), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(G190), .B2(new_n355), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n345), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT10), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n345), .A2(new_n347), .A3(new_n360), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n339), .B1(G169), .B2(new_n355), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n355), .A2(new_n298), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n327), .A2(G68), .A3(new_n328), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n300), .B1(new_n368), .B2(new_n203), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n369), .A2(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(KEYINPUT78), .ZN(new_n371));
  INV_X1    g0171(.A(new_n304), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G159), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n269), .A2(new_n271), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n300), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT76), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT76), .B1(new_n269), .B2(new_n271), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n300), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n202), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT76), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n270), .A2(G33), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT76), .ZN(new_n390));
  AOI21_X1  g0190(.A(G20), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n377), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT77), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT16), .B(new_n375), .C1(new_n385), .C2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n376), .B2(new_n300), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n202), .B1(new_n397), .B2(new_n377), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n395), .B1(new_n374), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n399), .A3(new_n307), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT79), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n265), .A2(G223), .A3(new_n272), .ZN(new_n402));
  INV_X1    g0202(.A(G87), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n402), .B1(new_n268), .B2(new_n403), .C1(new_n352), .C2(new_n348), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n275), .ZN(new_n405));
  INV_X1    g0205(.A(new_n261), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n251), .B1(new_n406), .B2(G232), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n401), .B1(new_n408), .B2(G190), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n410), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n321), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n333), .A2(new_n310), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n314), .B2(new_n333), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n400), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n417), .A2(KEYINPUT17), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n400), .A2(new_n416), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n408), .A2(new_n298), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n291), .B1(new_n405), .B2(new_n407), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT18), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  AOI211_X1 g0226(.A(new_n426), .B(new_n423), .C1(new_n400), .C2(new_n416), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n418), .A2(new_n419), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n310), .A2(new_n351), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT8), .B(G58), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n304), .B1(new_n300), .B2(new_n351), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT15), .B(G87), .Z(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n302), .B2(new_n432), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n429), .B1(new_n351), .B2(new_n314), .C1(new_n433), .C2(new_n313), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT70), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n406), .A2(G244), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n265), .A2(G232), .A3(new_n272), .ZN(new_n437));
  INV_X1    g0237(.A(G107), .ZN(new_n438));
  INV_X1    g0238(.A(G238), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n437), .B1(new_n438), .B2(new_n265), .C1(new_n352), .C2(new_n439), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n251), .B(new_n436), .C1(new_n440), .C2(new_n275), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G190), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n435), .B(new_n442), .C1(new_n321), .C2(new_n441), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n441), .A2(new_n298), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n434), .B1(new_n441), .B2(G169), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NOR4_X1   g0247(.A1(new_n323), .A2(new_n367), .A3(new_n428), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n269), .A2(new_n271), .A3(new_n300), .A4(G87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT22), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT22), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n265), .A2(new_n451), .A3(new_n300), .A4(G87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n300), .B2(G107), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n438), .A2(KEYINPUT23), .A3(G20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G116), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(G20), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n453), .A2(KEYINPUT24), .A3(new_n460), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n307), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(new_n272), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n265), .A2(new_n468), .A3(G250), .A4(new_n272), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n275), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(G274), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n275), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G264), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n473), .A2(G190), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n309), .B1(G1), .B2(new_n268), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n307), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n310), .A2(KEYINPUT25), .A3(new_n438), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n309), .B2(G107), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n484), .A2(G107), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n465), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n472), .A2(new_n275), .B1(G264), .B2(new_n480), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n321), .B1(new_n490), .B2(new_n479), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT87), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  INV_X1    g0293(.A(new_n488), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n313), .B1(new_n461), .B2(new_n462), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n464), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT87), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .A4(new_n482), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  AND4_X1   g0300(.A1(G179), .A2(new_n473), .A3(new_n479), .A4(new_n481), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n291), .B1(new_n490), .B2(new_n479), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n496), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n490), .A2(G179), .A3(new_n479), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(KEYINPUT86), .C1(new_n506), .C2(new_n291), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n438), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT6), .A2(G97), .ZN(new_n515));
  OR3_X1    g0315(.A1(new_n515), .A2(KEYINPUT80), .A3(G107), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT80), .B1(new_n515), .B2(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G20), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n372), .A2(G77), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n438), .B1(new_n397), .B2(new_n377), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n307), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n309), .A2(G97), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n484), .B2(G97), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(KEYINPUT81), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n372), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n378), .B2(new_n396), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n313), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n525), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(new_n272), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n275), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n248), .A2(G45), .A3(G274), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n474), .B2(new_n475), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n480), .B2(G257), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(KEYINPUT82), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT82), .B1(new_n541), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g0347(.A(G190), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(new_n544), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n533), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n291), .A3(new_n545), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n541), .A2(new_n298), .A3(new_n544), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n523), .A2(new_n525), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n300), .B1(new_n267), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n513), .A2(new_n403), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n269), .A2(new_n271), .A3(new_n300), .A4(G68), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n558), .B1(new_n301), .B2(new_n511), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n432), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n564), .A2(new_n307), .B1(new_n310), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n484), .A2(G87), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n269), .A2(new_n271), .A3(G238), .A4(new_n272), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n458), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n275), .ZN(new_n572));
  OAI21_X1  g0372(.A(G250), .B1(new_n477), .B2(G1), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n542), .B1(new_n275), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n568), .B(new_n577), .C1(new_n410), .C2(new_n576), .ZN(new_n578));
  INV_X1    g0378(.A(new_n484), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n566), .B1(new_n565), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n291), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n574), .B1(new_n571), .B2(new_n275), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n298), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n551), .A2(new_n557), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n543), .B1(new_n480), .B2(G270), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n272), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n590));
  INV_X1    g0390(.A(G303), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n265), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n275), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n291), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(KEYINPUT5), .A2(G41), .ZN(new_n595));
  NOR2_X1   g0395(.A1(KEYINPUT5), .A2(G41), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n478), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(G270), .A3(new_n254), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n479), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n275), .B2(new_n592), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n594), .A2(KEYINPUT21), .B1(new_n600), .B2(G179), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n309), .A2(G116), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n484), .B2(G116), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G20), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(G33), .B2(G283), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n268), .A2(G97), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT83), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT83), .B1(new_n607), .B2(new_n608), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n307), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT84), .B1(new_n601), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n611), .B(new_n612), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n603), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT84), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n600), .A2(new_n620), .A3(new_n291), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n588), .A2(new_n593), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n298), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n618), .B(new_n619), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n594), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n620), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(G200), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n615), .B(new_n628), .C1(new_n410), .C2(new_n622), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n509), .A2(new_n587), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n448), .A2(new_n631), .ZN(G372));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n425), .B2(new_n427), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n384), .B1(new_n383), .B2(new_n202), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n392), .A2(KEYINPUT77), .A3(G68), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n374), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n313), .B1(new_n637), .B2(KEYINPUT16), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n415), .B1(new_n638), .B2(new_n399), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n426), .B1(new_n639), .B2(new_n423), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n420), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(KEYINPUT90), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n446), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n322), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n318), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n417), .B(KEYINPUT17), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n646), .A2(new_n647), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n365), .B1(new_n652), .B2(new_n362), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n557), .A2(new_n585), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(KEYINPUT26), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n554), .A2(new_n555), .A3(new_n532), .A4(new_n526), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n566), .B(new_n567), .C1(new_n582), .C2(new_n321), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n576), .A2(new_n410), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT88), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n578), .A2(new_n662), .A3(new_n584), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n657), .A2(KEYINPUT89), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(new_n533), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT89), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n554), .A4(new_n555), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n618), .B1(new_n621), .B2(new_n623), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n627), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n504), .B1(new_n502), .B2(new_n501), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n661), .A2(new_n663), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n499), .A2(new_n674), .A3(new_n557), .A4(new_n551), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n656), .B(new_n669), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n448), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n653), .A2(new_n677), .ZN(G369));
  NOR2_X1   g0478(.A1(new_n208), .A2(G20), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n248), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n504), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT92), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n499), .A3(new_n508), .ZN(new_n688));
  INV_X1    g0488(.A(new_n685), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n508), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n671), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n615), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n630), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n625), .A2(new_n627), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n689), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n688), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n685), .B(KEYINPUT93), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n672), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n697), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n209), .A2(G41), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n560), .A2(G116), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n704), .A2(new_n248), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n225), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n704), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n622), .B2(new_n298), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(new_n490), .A3(new_n582), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n553), .A2(new_n545), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n600), .A2(KEYINPUT94), .A3(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n713), .A2(new_n716), .A3(new_n490), .A4(new_n582), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n546), .A2(new_n547), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n600), .A2(G179), .A3(new_n582), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n490), .A2(new_n479), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(new_n723), .A3(new_n549), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n717), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n717), .A2(new_n721), .A3(KEYINPUT96), .A4(new_n724), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n685), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  INV_X1    g0530(.A(new_n701), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(new_n730), .B1(new_n631), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT95), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n711), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n557), .A2(new_n585), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n654), .B1(new_n736), .B2(new_n665), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n508), .A2(new_n625), .A3(new_n627), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n675), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n665), .B1(new_n664), .B2(new_n668), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n689), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT98), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n551), .A2(new_n557), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n508), .A2(new_n625), .A3(new_n627), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n499), .A4(new_n674), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n664), .A2(new_n668), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n746), .B(new_n737), .C1(new_n747), .C2(new_n665), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT98), .B1(new_n748), .B2(new_n689), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT29), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n676), .A2(new_n731), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n735), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n710), .B1(new_n754), .B2(G1), .ZN(G364));
  OR2_X1    g0555(.A1(new_n695), .A2(G330), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT99), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n248), .B1(new_n679), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n704), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(KEYINPUT99), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n757), .A2(new_n696), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n221), .B1(G20), .B2(new_n291), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n300), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n321), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n265), .B1(new_n768), .B2(new_n438), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n298), .A2(new_n321), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n766), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n298), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G68), .A2(new_n772), .B1(new_n775), .B2(G77), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n300), .A2(new_n410), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n767), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n773), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n776), .B1(new_n403), .B2(new_n778), .C1(new_n329), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n770), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT102), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(KEYINPUT102), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n769), .B(new_n780), .C1(G50), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G179), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n766), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT103), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT32), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n300), .B1(new_n788), .B2(G190), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n792), .A2(new_n793), .B1(G97), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n787), .B(new_n799), .C1(new_n793), .C2(new_n792), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n778), .A2(new_n591), .B1(new_n768), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n772), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n779), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n265), .B1(new_n805), .B2(G322), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G311), .A2(new_n775), .B1(new_n790), .B2(G329), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n786), .A2(G326), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n797), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n765), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n765), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n389), .A2(new_n390), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n210), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT101), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n708), .A2(new_n477), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n477), .C2(new_n246), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n210), .A2(new_n265), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT100), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G355), .B1(new_n605), .B2(new_n209), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n817), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n812), .A2(new_n826), .A3(new_n761), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n695), .B2(new_n816), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT105), .Z(new_n829));
  NAND2_X1  g0629(.A1(new_n763), .A2(new_n829), .ZN(G396));
  OAI22_X1  g0630(.A1(new_n801), .A2(new_n771), .B1(new_n779), .B2(new_n810), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n778), .A2(new_n438), .B1(new_n768), .B2(new_n403), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n376), .B1(new_n774), .B2(new_n605), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n789), .A2(new_n834), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n511), .B2(new_n797), .C1(new_n591), .C2(new_n785), .ZN(new_n837));
  XOR2_X1   g0637(.A(KEYINPUT106), .B(G143), .Z(new_n838));
  AOI22_X1  g0638(.A1(new_n805), .A2(new_n838), .B1(new_n775), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n325), .B2(new_n771), .C1(new_n785), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n778), .A2(new_n241), .B1(new_n789), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n768), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n818), .B(new_n845), .C1(G68), .C2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n843), .B(new_n847), .C1(new_n329), .C2(new_n797), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n841), .A2(new_n842), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n764), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n764), .A2(new_n813), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n761), .B1(new_n351), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n446), .A2(new_n685), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n434), .A2(new_n685), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n443), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n856), .B2(new_n446), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n851), .B(new_n853), .C1(new_n857), .C2(new_n814), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n751), .B(new_n857), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n735), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n760), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(new_n224), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(G116), .C1(KEYINPUT35), .C2(new_n518), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(KEYINPUT35), .B2(new_n518), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  AND3_X1   g0669(.A1(new_n708), .A2(G77), .A3(new_n368), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n242), .B(KEYINPUT107), .ZN(new_n871));
  OAI211_X1 g0671(.A(G1), .B(new_n208), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT108), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n294), .A2(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n289), .A2(KEYINPUT14), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n317), .B(new_n685), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT109), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n299), .A2(KEYINPUT109), .A3(new_n317), .A4(new_n685), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n317), .A2(new_n685), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n318), .A2(new_n322), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n729), .A2(new_n730), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n631), .A2(new_n731), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n685), .A4(new_n728), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n857), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  INV_X1    g0689(.A(new_n683), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n420), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n643), .B2(new_n649), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT90), .A3(new_n417), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n420), .A2(new_n424), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n891), .A3(new_n417), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n891), .A2(new_n417), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(new_n633), .A3(KEYINPUT37), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n889), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n637), .A2(KEYINPUT16), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n415), .B1(new_n902), .B2(new_n638), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n428), .A2(new_n890), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n423), .A2(new_n683), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n639), .B2(new_n413), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n906), .A2(new_n896), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n888), .B1(new_n901), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n896), .A2(new_n906), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n909), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n904), .A2(new_n890), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n640), .A2(new_n641), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n649), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n889), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n911), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n913), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n912), .A2(new_n913), .B1(new_n888), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G330), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n711), .B1(new_n732), .B2(new_n886), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n448), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n448), .A3(new_n887), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n299), .A2(new_n317), .A3(new_n689), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n901), .A2(new_n931), .A3(new_n911), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n921), .A2(KEYINPUT39), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n676), .A2(new_n731), .A3(new_n857), .ZN(new_n935));
  INV_X1    g0735(.A(new_n854), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n921), .A2(new_n937), .A3(new_n883), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n643), .B2(new_n890), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n929), .B(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n750), .A2(new_n448), .A3(new_n753), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT110), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n750), .A2(new_n945), .A3(new_n448), .A4(new_n753), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n653), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n942), .A2(new_n948), .B1(new_n248), .B2(new_n679), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n942), .A2(new_n948), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n869), .B(new_n873), .C1(new_n949), .C2(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n789), .A2(new_n840), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n768), .A2(new_n351), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G159), .C2(new_n772), .ZN(new_n954));
  INV_X1    g0754(.A(new_n778), .ZN(new_n955));
  INV_X1    g0755(.A(new_n329), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n376), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G150), .A2(new_n805), .B1(new_n775), .B2(G50), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n838), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n202), .B2(new_n797), .C1(new_n785), .C2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n797), .A2(new_n438), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G294), .A2(new_n772), .B1(new_n790), .B2(G317), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n801), .B2(new_n774), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G311), .B2(new_n786), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n768), .A2(new_n511), .ZN(new_n966));
  INV_X1    g0766(.A(new_n818), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(G303), .C2(new_n805), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n955), .A2(G116), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT46), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n961), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT47), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n765), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n973), .B2(new_n972), .ZN(new_n975));
  INV_X1    g0775(.A(new_n236), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n820), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n817), .B1(new_n209), .B2(new_n432), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n761), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n568), .A2(new_n689), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n654), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n674), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n981), .B1(new_n982), .B2(new_n980), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n975), .B(new_n979), .C1(new_n983), .C2(new_n816), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n551), .B(new_n557), .C1(new_n533), .C2(new_n731), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT111), .ZN(new_n986));
  INV_X1    g0786(.A(new_n657), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n986), .B1(new_n987), .B2(new_n701), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n702), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n702), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n702), .A2(KEYINPUT44), .A3(new_n988), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT44), .B1(new_n702), .B2(new_n988), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n990), .A2(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n697), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n691), .A2(new_n699), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n700), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(new_n696), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n754), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n704), .B(KEYINPUT41), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n759), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n983), .B(KEYINPUT43), .Z(new_n1003));
  OR3_X1    g0803(.A1(new_n988), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT42), .B1(new_n988), .B2(new_n700), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n557), .B1(new_n988), .B2(new_n508), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1007), .A2(new_n731), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1003), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT112), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n1006), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(KEYINPUT112), .B(new_n1003), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n988), .A2(new_n696), .A3(new_n691), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1015), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n984), .B1(new_n1002), .B2(new_n1018), .ZN(G387));
  AOI22_X1  g0819(.A1(new_n786), .A2(G159), .B1(new_n333), .B2(new_n772), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n798), .A2(new_n432), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n779), .A2(new_n241), .B1(new_n789), .B2(new_n325), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G77), .B2(new_n955), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n966), .B(new_n818), .C1(G68), .C2(new_n775), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G116), .A2(new_n846), .B1(new_n790), .B2(G326), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G311), .A2(new_n772), .B1(new_n775), .B2(G303), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(new_n779), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G322), .B2(new_n786), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n797), .A2(new_n801), .B1(new_n810), .B2(new_n778), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n818), .B(new_n1026), .C1(new_n1033), .C2(KEYINPUT49), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n764), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n430), .A2(G50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n477), .B1(new_n202), .B2(new_n351), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n705), .B2(KEYINPUT113), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(KEYINPUT113), .C2(new_n705), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n820), .B(new_n1042), .C1(new_n477), .C2(new_n233), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n824), .A2(new_n706), .B1(new_n438), .B2(new_n209), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n817), .B1(new_n1045), .B2(KEYINPUT114), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n761), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1037), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n691), .B2(new_n815), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n999), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n759), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n754), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n704), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1051), .A2(new_n754), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(G393));
  NAND2_X1  g0856(.A1(new_n988), .A2(new_n815), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n778), .A2(new_n202), .B1(new_n774), .B2(new_n430), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n967), .B1(new_n403), .B2(new_n768), .C1(new_n789), .C2(new_n960), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G50), .C2(new_n772), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n786), .A2(G150), .B1(G159), .B2(new_n805), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n798), .A2(G77), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n376), .B1(new_n768), .B2(new_n438), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G294), .A2(new_n775), .B1(new_n790), .B2(G322), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n801), .B2(new_n778), .C1(new_n591), .C2(new_n771), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G116), .C2(new_n798), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n785), .A2(new_n1028), .B1(new_n834), .B2(new_n779), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n765), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n820), .A2(new_n240), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n817), .B1(new_n209), .B2(G97), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n761), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1057), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n996), .B2(new_n758), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n996), .A2(new_n1053), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n704), .B1(new_n996), .B2(new_n1053), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(G390));
  AND4_X1   g0883(.A1(G330), .A2(new_n883), .A3(new_n857), .A4(new_n887), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n883), .B1(new_n735), .B2(new_n857), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n937), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n887), .A2(G330), .A3(new_n857), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n882), .A3(new_n880), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n741), .A2(new_n742), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n748), .A2(KEYINPUT98), .A3(new_n689), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n936), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n856), .A2(new_n446), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n735), .A2(new_n857), .A3(new_n883), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1088), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1096));
  AND4_X1   g0896(.A1(new_n653), .A2(new_n947), .A3(new_n1096), .A4(new_n926), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n937), .A2(new_n883), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n930), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n932), .A2(new_n1100), .A3(new_n933), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n930), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n901), .B2(new_n911), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1091), .A2(new_n1092), .A3(new_n883), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1103), .A2(KEYINPUT116), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT116), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1101), .B(new_n1094), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n932), .A2(new_n933), .A3(new_n1100), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n425), .A2(new_n427), .A3(new_n633), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT90), .B1(new_n640), .B2(new_n641), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n649), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n891), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n897), .A2(new_n899), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT38), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n911), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n930), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1091), .A2(new_n1092), .A3(new_n883), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1109), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1103), .A2(KEYINPUT116), .A3(new_n1104), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1108), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1084), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1107), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1098), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1084), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1097), .A2(new_n1127), .A3(new_n1107), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n704), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1127), .A2(new_n759), .A3(new_n1107), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT119), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n932), .A2(new_n933), .A3(new_n813), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n852), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n760), .B1(new_n333), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT117), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n786), .A2(G283), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n779), .A2(new_n605), .B1(new_n768), .B2(new_n202), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n265), .B(new_n1138), .C1(G87), .C2(new_n955), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n771), .A2(new_n438), .B1(new_n774), .B2(new_n511), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G294), .B2(new_n790), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1065), .A4(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT54), .B(G143), .Z(new_n1143));
  AOI22_X1  g0943(.A1(G137), .A2(new_n772), .B1(new_n775), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G132), .A2(new_n805), .B1(new_n790), .B2(G125), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n786), .B2(G128), .ZN(new_n1147));
  INV_X1    g0947(.A(G159), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n797), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n778), .A2(new_n325), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n265), .B1(new_n768), .B2(new_n241), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT118), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1142), .B1(new_n1149), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1136), .B1(new_n1157), .B2(new_n764), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1133), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1131), .A2(new_n1132), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1132), .B1(new_n1131), .B2(new_n1159), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1130), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G378));
  NAND3_X1  g0963(.A1(new_n341), .A2(new_n344), .A3(new_n890), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n367), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n367), .A2(new_n1165), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n813), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n760), .B1(G50), .B2(new_n1134), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n967), .A2(G41), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1176), .B(new_n241), .C1(G33), .C2(G41), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT120), .Z(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(G116), .B2(new_n786), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n846), .A2(new_n956), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n511), .B2(new_n771), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n351), .A2(new_n778), .B1(new_n779), .B2(new_n438), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n565), .A2(new_n774), .B1(new_n801), .B2(new_n789), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1179), .B(new_n1184), .C1(new_n202), .C2(new_n797), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1178), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n786), .A2(G125), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n798), .A2(G150), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n772), .B1(new_n775), .B2(G137), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1143), .A2(new_n955), .B1(new_n805), .B2(G128), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n846), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1188), .B1(new_n1186), .B2(new_n1185), .C1(new_n1194), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1174), .B1(new_n1199), .B2(new_n764), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1173), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1172), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n923), .A2(G330), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n923), .B2(G330), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n941), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n924), .A2(new_n1172), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n923), .A2(G330), .A3(new_n1203), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n940), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1202), .B1(new_n1210), .B2(new_n759), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT121), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n947), .A2(new_n653), .A3(new_n926), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1096), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1216), .B1(new_n1124), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT57), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1128), .A2(new_n1216), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n704), .B1(new_n1221), .B2(KEYINPUT57), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1211), .B1(new_n1220), .B2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1098), .A2(new_n1001), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n880), .A2(new_n813), .A3(new_n882), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1134), .A2(G68), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G97), .A2(new_n955), .B1(new_n772), .B2(G116), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n438), .B2(new_n774), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n779), .A2(new_n801), .B1(new_n789), .B2(new_n591), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1229), .A2(new_n265), .A3(new_n953), .A4(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n1021), .C1(new_n810), .C2(new_n785), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT122), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n840), .A2(new_n779), .B1(new_n778), .B2(new_n1148), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n772), .A2(new_n1143), .B1(new_n790), .B2(G128), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n325), .B2(new_n774), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(G132), .C2(new_n786), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n967), .A2(new_n1180), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1238), .A2(new_n1239), .B1(new_n798), .B2(G50), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1237), .B(new_n1240), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1232), .A2(KEYINPUT122), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1233), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n761), .B(new_n1227), .C1(new_n1243), .C2(new_n764), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1096), .A2(new_n759), .B1(new_n1226), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1225), .A2(new_n1245), .ZN(G381));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  INV_X1    g1048(.A(G396), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1052), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1251), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1252), .A2(G387), .A3(G381), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT124), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1211), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n704), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1218), .A2(new_n1210), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT57), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(KEYINPUT57), .B(new_n1218), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1255), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1254), .A2(new_n1162), .A3(new_n1261), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1162), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G407), .B(G213), .C1(G343), .C2(new_n1263), .ZN(G409));
  NAND2_X1  g1064(.A1(new_n684), .A2(G213), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1202), .B1(new_n1221), .B2(new_n1001), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n759), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1129), .A4(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1265), .B(new_n1269), .C1(new_n1261), .C2(new_n1162), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1224), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1215), .A2(KEYINPUT60), .A3(new_n1217), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1098), .A3(new_n704), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1245), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1248), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(G384), .A3(new_n1245), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT62), .B1(new_n1270), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1276), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1269), .A2(new_n1265), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G375), .A2(G378), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1278), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1279), .A2(new_n1284), .A3(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(new_n1251), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1292), .A2(KEYINPUT125), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(KEYINPUT125), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1247), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G390), .B(new_n984), .C1(new_n1002), .C2(new_n1018), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1301), .A3(new_n1295), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1298), .A2(new_n1292), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1290), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1270), .B2(new_n1278), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1285), .A2(new_n1286), .A3(KEYINPUT63), .A4(new_n1288), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1304), .A2(new_n1308), .A3(new_n1284), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1306), .A2(new_n1310), .ZN(G405));
  NAND2_X1  g1111(.A1(new_n1286), .A2(new_n1263), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1288), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1286), .A2(new_n1263), .A3(new_n1278), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1304), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1305), .A2(new_n1314), .A3(new_n1313), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


