

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753;

  NOR2_X1 U369 ( .A1(n717), .A2(n723), .ZN(n718) );
  XNOR2_X2 U370 ( .A(G128), .B(G143), .ZN(n471) );
  NOR2_X2 U371 ( .A1(n624), .A2(n723), .ZN(n625) );
  XNOR2_X2 U372 ( .A(n394), .B(n393), .ZN(n731) );
  XNOR2_X1 U373 ( .A(n385), .B(n384), .ZN(n708) );
  XNOR2_X1 U374 ( .A(G472), .B(n508), .ZN(n614) );
  NOR2_X1 U375 ( .A1(n631), .A2(n723), .ZN(n634) );
  NOR2_X1 U376 ( .A1(n639), .A2(n723), .ZN(n641) );
  INV_X1 U377 ( .A(n398), .ZN(n348) );
  NOR2_X1 U378 ( .A1(n708), .A2(n596), .ZN(n597) );
  NOR2_X1 U379 ( .A1(n594), .A2(n593), .ZN(n449) );
  NOR2_X1 U380 ( .A1(n713), .A2(G902), .ZN(n520) );
  INV_X1 U381 ( .A(KEYINPUT110), .ZN(n455) );
  INV_X1 U382 ( .A(KEYINPUT66), .ZN(n448) );
  INV_X1 U383 ( .A(n398), .ZN(n349) );
  XNOR2_X1 U384 ( .A(n456), .B(n455), .ZN(n697) );
  XNOR2_X1 U385 ( .A(n449), .B(n447), .ZN(n616) );
  NAND2_X1 U386 ( .A1(n692), .A2(n691), .ZN(n456) );
  XNOR2_X1 U387 ( .A(n406), .B(n356), .ZN(n692) );
  XNOR2_X1 U388 ( .A(n527), .B(n526), .ZN(n557) );
  XOR2_X1 U389 ( .A(n714), .B(KEYINPUT59), .Z(n716) );
  XNOR2_X1 U390 ( .A(n404), .B(n481), .ZN(n719) );
  XNOR2_X1 U391 ( .A(n383), .B(n417), .ZN(n513) );
  XNOR2_X1 U392 ( .A(n500), .B(n499), .ZN(n383) );
  XNOR2_X1 U393 ( .A(n473), .B(n472), .ZN(n500) );
  INV_X1 U394 ( .A(n489), .ZN(n744) );
  XNOR2_X1 U395 ( .A(n595), .B(n448), .ZN(n447) );
  XNOR2_X1 U396 ( .A(KEYINPUT64), .B(G953), .ZN(n489) );
  XNOR2_X1 U397 ( .A(KEYINPUT4), .B(KEYINPUT68), .ZN(n499) );
  NAND2_X1 U398 ( .A1(n650), .A2(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U399 ( .A(n411), .B(n410), .ZN(n479) );
  INV_X1 U400 ( .A(KEYINPUT8), .ZN(n410) );
  NAND2_X1 U401 ( .A1(n744), .A2(G234), .ZN(n411) );
  XNOR2_X1 U402 ( .A(KEYINPUT65), .B(KEYINPUT79), .ZN(n472) );
  XNOR2_X1 U403 ( .A(G125), .B(G146), .ZN(n522) );
  XNOR2_X1 U404 ( .A(G137), .B(G140), .ZN(n512) );
  XNOR2_X1 U405 ( .A(n355), .B(n414), .ZN(n573) );
  XNOR2_X1 U406 ( .A(n415), .B(G478), .ZN(n414) );
  INV_X1 U407 ( .A(KEYINPUT99), .ZN(n415) );
  XNOR2_X1 U408 ( .A(n459), .B(KEYINPUT39), .ZN(n585) );
  NAND2_X1 U409 ( .A1(n571), .A2(n692), .ZN(n459) );
  XNOR2_X1 U410 ( .A(n354), .B(KEYINPUT82), .ZN(n558) );
  XNOR2_X1 U411 ( .A(n400), .B(n399), .ZN(n463) );
  INV_X1 U412 ( .A(KEYINPUT81), .ZN(n399) );
  NOR2_X1 U413 ( .A1(n612), .A2(n392), .ZN(n388) );
  NOR2_X1 U414 ( .A1(n642), .A2(n364), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n620), .B(n365), .ZN(n364) );
  INV_X1 U416 ( .A(KEYINPUT101), .ZN(n365) );
  INV_X1 U417 ( .A(KEYINPUT45), .ZN(n393) );
  NAND2_X1 U418 ( .A1(n366), .A2(n361), .ZN(n394) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n361) );
  NOR2_X1 U420 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U421 ( .A(n408), .B(n407), .ZN(n577) );
  XNOR2_X1 U422 ( .A(n446), .B(n445), .ZN(n444) );
  XNOR2_X1 U423 ( .A(n522), .B(KEYINPUT78), .ZN(n445) );
  XOR2_X1 U424 ( .A(G902), .B(KEYINPUT15), .Z(n525) );
  OR2_X1 U425 ( .A1(n589), .A2(n676), .ZN(n416) );
  XNOR2_X1 U426 ( .A(n435), .B(n350), .ZN(n673) );
  OR2_X1 U427 ( .A1(n719), .A2(G902), .ZN(n435) );
  XNOR2_X1 U428 ( .A(n566), .B(KEYINPUT1), .ZN(n589) );
  XNOR2_X1 U429 ( .A(n530), .B(n529), .ZN(n594) );
  XNOR2_X1 U430 ( .A(G101), .B(G146), .ZN(n504) );
  XOR2_X1 U431 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n461) );
  XNOR2_X1 U432 ( .A(G119), .B(G110), .ZN(n482) );
  XOR2_X1 U433 ( .A(G131), .B(G104), .Z(n536) );
  XNOR2_X1 U434 ( .A(G122), .B(G113), .ZN(n535) );
  XOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n538) );
  XNOR2_X1 U436 ( .A(n522), .B(KEYINPUT10), .ZN(n736) );
  NAND2_X1 U437 ( .A1(n423), .A2(n525), .ZN(n422) );
  NAND2_X1 U438 ( .A1(n731), .A2(n426), .ZN(n423) );
  XNOR2_X1 U439 ( .A(n513), .B(n512), .ZN(n737) );
  NOR2_X1 U440 ( .A1(n422), .A2(n375), .ZN(n374) );
  INV_X1 U441 ( .A(G210), .ZN(n375) );
  AND2_X1 U442 ( .A1(n436), .A2(n352), .ZN(n576) );
  INV_X1 U443 ( .A(n570), .ZN(n406) );
  AND2_X1 U444 ( .A1(n555), .A2(n556), .ZN(n571) );
  XNOR2_X1 U445 ( .A(n554), .B(KEYINPUT77), .ZN(n555) );
  INV_X1 U446 ( .A(n673), .ZN(n613) );
  BUF_X1 U447 ( .A(n589), .Z(n677) );
  XNOR2_X1 U448 ( .A(G475), .B(n545), .ZN(n572) );
  INV_X1 U449 ( .A(n677), .ZN(n371) );
  INV_X1 U450 ( .A(n613), .ZN(n437) );
  BUF_X1 U451 ( .A(n744), .Z(n403) );
  BUF_X1 U452 ( .A(G953), .Z(n409) );
  XNOR2_X1 U453 ( .A(n369), .B(n368), .ZN(n623) );
  XNOR2_X1 U454 ( .A(n470), .B(KEYINPUT9), .ZN(n368) );
  XNOR2_X1 U455 ( .A(n474), .B(n475), .ZN(n369) );
  NOR2_X1 U456 ( .A1(n422), .A2(n381), .ZN(n380) );
  INV_X1 U457 ( .A(G478), .ZN(n381) );
  XNOR2_X1 U458 ( .A(n737), .B(n460), .ZN(n713) );
  XNOR2_X1 U459 ( .A(n516), .B(n524), .ZN(n460) );
  XNOR2_X1 U460 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U461 ( .A(G146), .ZN(n514) );
  NOR2_X1 U462 ( .A1(n403), .A2(G952), .ZN(n723) );
  INV_X1 U463 ( .A(n409), .ZN(n359) );
  INV_X1 U464 ( .A(KEYINPUT44), .ZN(n392) );
  NOR2_X1 U465 ( .A1(n558), .A2(n433), .ZN(n431) );
  INV_X1 U466 ( .A(KEYINPUT103), .ZN(n362) );
  NAND2_X1 U467 ( .A1(n357), .A2(n390), .ZN(n366) );
  NAND2_X1 U468 ( .A1(n389), .A2(n388), .ZN(n390) );
  AND2_X1 U469 ( .A1(n367), .A2(n391), .ZN(n357) );
  INV_X1 U470 ( .A(KEYINPUT46), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n521), .B(n353), .ZN(n446) );
  NAND2_X1 U472 ( .A1(G224), .A2(n744), .ZN(n521) );
  XOR2_X1 U473 ( .A(n494), .B(KEYINPUT21), .Z(n674) );
  XOR2_X1 U474 ( .A(G137), .B(KEYINPUT5), .Z(n502) );
  NOR2_X1 U475 ( .A1(n409), .A2(G237), .ZN(n532) );
  NOR2_X1 U476 ( .A1(n426), .A2(n420), .ZN(n419) );
  XNOR2_X1 U477 ( .A(G134), .B(G131), .ZN(n417) );
  OR2_X1 U478 ( .A1(G902), .A2(G237), .ZN(n528) );
  XNOR2_X1 U479 ( .A(n497), .B(n401), .ZN(n562) );
  INV_X1 U480 ( .A(KEYINPUT70), .ZN(n401) );
  NOR2_X1 U481 ( .A1(n673), .A2(n496), .ZN(n497) );
  XNOR2_X1 U482 ( .A(G107), .B(G134), .ZN(n464) );
  XNOR2_X1 U483 ( .A(n360), .B(KEYINPUT97), .ZN(n465) );
  INV_X1 U484 ( .A(KEYINPUT98), .ZN(n360) );
  XNOR2_X1 U485 ( .A(n467), .B(n466), .ZN(n468) );
  INV_X1 U486 ( .A(KEYINPUT96), .ZN(n466) );
  XNOR2_X1 U487 ( .A(G122), .B(G116), .ZN(n467) );
  XNOR2_X1 U488 ( .A(n511), .B(n510), .ZN(n524) );
  BUF_X1 U489 ( .A(n731), .Z(n402) );
  XOR2_X1 U490 ( .A(KEYINPUT88), .B(n677), .Z(n601) );
  INV_X1 U491 ( .A(KEYINPUT33), .ZN(n384) );
  NAND2_X1 U492 ( .A1(n576), .A2(n531), .ZN(n650) );
  NAND2_X1 U493 ( .A1(n349), .A2(n376), .ZN(n638) );
  NOR2_X1 U494 ( .A1(n422), .A2(n377), .ZN(n376) );
  INV_X1 U495 ( .A(G472), .ZN(n377) );
  XNOR2_X1 U496 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U497 ( .A(n440), .B(n524), .ZN(n724) );
  XNOR2_X1 U498 ( .A(n523), .B(n441), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n442), .B(KEYINPUT75), .ZN(n441) );
  XNOR2_X1 U500 ( .A(G122), .B(KEYINPUT16), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n480), .B(n483), .ZN(n404) );
  XNOR2_X1 U502 ( .A(n541), .B(n397), .ZN(n714) );
  XNOR2_X1 U503 ( .A(n542), .B(n736), .ZN(n397) );
  NAND2_X1 U504 ( .A1(n348), .A2(n378), .ZN(n715) );
  NOR2_X1 U505 ( .A1(n422), .A2(n379), .ZN(n378) );
  INV_X1 U506 ( .A(G475), .ZN(n379) );
  XNOR2_X1 U507 ( .A(n628), .B(n627), .ZN(n629) );
  NAND2_X1 U508 ( .A1(n349), .A2(n374), .ZN(n630) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n752) );
  XNOR2_X1 U510 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(n753) );
  INV_X1 U512 ( .A(KEYINPUT40), .ZN(n457) );
  AND2_X1 U513 ( .A1(n598), .A2(n406), .ZN(n405) );
  AND2_X1 U514 ( .A1(n438), .A2(n437), .ZN(n642) );
  NOR2_X1 U515 ( .A1(n386), .A2(n371), .ZN(n370) );
  NAND2_X1 U516 ( .A1(n348), .A2(n380), .ZN(n622) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n452) );
  XNOR2_X1 U518 ( .A(n713), .B(n712), .ZN(n453) );
  NAND2_X1 U519 ( .A1(n711), .A2(n359), .ZN(n358) );
  XOR2_X1 U520 ( .A(n486), .B(n485), .Z(n350) );
  XOR2_X1 U521 ( .A(G113), .B(G119), .Z(n351) );
  XNOR2_X1 U522 ( .A(n566), .B(KEYINPUT109), .ZN(n352) );
  XNOR2_X1 U523 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n353) );
  AND2_X1 U524 ( .A1(n571), .A2(n405), .ZN(n354) );
  NOR2_X1 U525 ( .A1(n623), .A2(G902), .ZN(n355) );
  XOR2_X1 U526 ( .A(KEYINPUT38), .B(KEYINPUT76), .Z(n356) );
  INV_X1 U527 ( .A(n525), .ZN(n621) );
  INV_X1 U528 ( .A(KEYINPUT2), .ZN(n426) );
  NAND2_X1 U529 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U530 ( .A1(n672), .A2(n358), .ZN(n395) );
  NAND2_X1 U531 ( .A1(n748), .A2(n392), .ZN(n367) );
  NOR2_X1 U532 ( .A1(n610), .A2(n386), .ZN(n373) );
  NAND2_X1 U533 ( .A1(n372), .A2(n370), .ZN(n439) );
  INV_X1 U534 ( .A(n610), .ZN(n372) );
  NAND2_X1 U535 ( .A1(n373), .A2(n607), .ZN(n608) );
  NOR2_X1 U536 ( .A1(n398), .A2(n422), .ZN(n382) );
  NAND2_X1 U537 ( .A1(n382), .A2(G217), .ZN(n720) );
  NAND2_X1 U538 ( .A1(n382), .A2(G469), .ZN(n454) );
  XNOR2_X1 U539 ( .A(n383), .B(n444), .ZN(n443) );
  NAND2_X1 U540 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U541 ( .A(n606), .ZN(n386) );
  XNOR2_X1 U542 ( .A(n416), .B(KEYINPUT105), .ZN(n387) );
  INV_X1 U543 ( .A(n748), .ZN(n389) );
  NAND2_X1 U544 ( .A1(n612), .A2(n392), .ZN(n391) );
  XNOR2_X1 U545 ( .A(n715), .B(n716), .ZN(n717) );
  XNOR2_X1 U546 ( .A(n395), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U547 ( .A1(n396), .A2(n616), .ZN(n605) );
  XNOR2_X1 U548 ( .A(n604), .B(KEYINPUT102), .ZN(n396) );
  XNOR2_X1 U549 ( .A(n439), .B(KEYINPUT85), .ZN(n438) );
  XNOR2_X1 U550 ( .A(n443), .B(n724), .ZN(n626) );
  NOR2_X1 U551 ( .A1(n753), .A2(n752), .ZN(n408) );
  XNOR2_X1 U552 ( .A(n579), .B(KEYINPUT48), .ZN(n588) );
  NAND2_X1 U553 ( .A1(n425), .A2(n424), .ZN(n398) );
  XNOR2_X2 U554 ( .A(n600), .B(KEYINPUT35), .ZN(n748) );
  NOR2_X1 U555 ( .A1(n562), .A2(n614), .ZN(n509) );
  XNOR2_X1 U556 ( .A(n434), .B(n569), .ZN(n578) );
  NOR2_X2 U557 ( .A1(n676), .A2(n566), .ZN(n617) );
  XNOR2_X2 U558 ( .A(n608), .B(KEYINPUT32), .ZN(n750) );
  XNOR2_X1 U559 ( .A(n412), .B(n477), .ZN(n478) );
  XNOR2_X1 U560 ( .A(n461), .B(n476), .ZN(n412) );
  NAND2_X1 U561 ( .A1(n585), .A2(n657), .ZN(n458) );
  NAND2_X1 U562 ( .A1(n427), .A2(n462), .ZN(n434) );
  AND2_X1 U563 ( .A1(n413), .A2(n432), .ZN(n429) );
  NAND2_X1 U564 ( .A1(n558), .A2(n433), .ZN(n413) );
  XNOR2_X1 U565 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U566 ( .A1(n416), .A2(n614), .ZN(n686) );
  NAND2_X1 U567 ( .A1(n588), .A2(n587), .ZN(n743) );
  NAND2_X1 U568 ( .A1(n421), .A2(n418), .ZN(n425) );
  AND2_X1 U569 ( .A1(n588), .A2(n419), .ZN(n418) );
  INV_X1 U570 ( .A(n587), .ZN(n420) );
  INV_X1 U571 ( .A(n731), .ZN(n421) );
  NOR2_X1 U572 ( .A1(n743), .A2(n402), .ZN(n667) );
  NAND2_X1 U573 ( .A1(n743), .A2(n426), .ZN(n424) );
  NAND2_X1 U574 ( .A1(n429), .A2(n428), .ZN(n427) );
  NAND2_X1 U575 ( .A1(n430), .A2(n431), .ZN(n428) );
  INV_X1 U576 ( .A(n559), .ZN(n430) );
  NAND2_X1 U577 ( .A1(n559), .A2(n433), .ZN(n432) );
  INV_X1 U578 ( .A(KEYINPUT80), .ZN(n433) );
  XNOR2_X1 U579 ( .A(n509), .B(KEYINPUT28), .ZN(n436) );
  XNOR2_X1 U580 ( .A(n478), .B(n736), .ZN(n481) );
  NAND2_X1 U581 ( .A1(n688), .A2(n576), .ZN(n451) );
  NOR2_X1 U582 ( .A1(n452), .A2(n723), .ZN(G54) );
  INV_X1 U583 ( .A(n557), .ZN(n570) );
  AND2_X1 U584 ( .A1(n568), .A2(n663), .ZN(n462) );
  INV_X1 U585 ( .A(KEYINPUT69), .ZN(n569) );
  INV_X1 U586 ( .A(KEYINPUT19), .ZN(n529) );
  INV_X1 U587 ( .A(n551), .ZN(n552) );
  INV_X1 U588 ( .A(n664), .ZN(n586) );
  INV_X1 U589 ( .A(KEYINPUT0), .ZN(n595) );
  NOR2_X1 U590 ( .A1(n665), .A2(n586), .ZN(n587) );
  INV_X1 U591 ( .A(n573), .ZN(n546) );
  NAND2_X1 U592 ( .A1(n479), .A2(G217), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n465), .B(n464), .ZN(n469) );
  INV_X1 U594 ( .A(n471), .ZN(n473) );
  XNOR2_X1 U595 ( .A(n500), .B(KEYINPUT7), .ZN(n474) );
  XOR2_X1 U596 ( .A(KEYINPUT90), .B(KEYINPUT83), .Z(n477) );
  XNOR2_X1 U597 ( .A(G128), .B(KEYINPUT89), .ZN(n476) );
  NAND2_X1 U598 ( .A1(G221), .A2(n479), .ZN(n480) );
  XNOR2_X1 U599 ( .A(n482), .B(n512), .ZN(n483) );
  XOR2_X1 U600 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n486) );
  NAND2_X1 U601 ( .A1(G234), .A2(n621), .ZN(n484) );
  XNOR2_X1 U602 ( .A(KEYINPUT20), .B(n484), .ZN(n493) );
  NAND2_X1 U603 ( .A1(n493), .A2(G217), .ZN(n485) );
  NAND2_X1 U604 ( .A1(G237), .A2(G234), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n487), .B(KEYINPUT14), .ZN(n488) );
  NAND2_X1 U606 ( .A1(G952), .A2(n488), .ZN(n706) );
  NOR2_X1 U607 ( .A1(n409), .A2(n706), .ZN(n592) );
  NAND2_X1 U608 ( .A1(G902), .A2(n488), .ZN(n590) );
  NOR2_X1 U609 ( .A1(G900), .A2(n590), .ZN(n490) );
  NAND2_X1 U610 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U611 ( .A(KEYINPUT106), .B(n491), .Z(n492) );
  NOR2_X1 U612 ( .A1(n592), .A2(n492), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G221), .A2(n493), .ZN(n494) );
  INV_X1 U614 ( .A(n674), .ZN(n603) );
  NOR2_X1 U615 ( .A1(n551), .A2(n603), .ZN(n495) );
  XNOR2_X1 U616 ( .A(n495), .B(KEYINPUT71), .ZN(n496) );
  XNOR2_X1 U617 ( .A(G116), .B(KEYINPUT3), .ZN(n498) );
  XNOR2_X1 U618 ( .A(n351), .B(n498), .ZN(n523) );
  XNOR2_X1 U619 ( .A(n513), .B(n523), .ZN(n507) );
  NAND2_X1 U620 ( .A1(n532), .A2(G210), .ZN(n501) );
  XNOR2_X1 U621 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U622 ( .A(n503), .B(KEYINPUT92), .Z(n505) );
  XNOR2_X1 U623 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U624 ( .A(n507), .B(n506), .ZN(n636) );
  NOR2_X1 U625 ( .A1(G902), .A2(n636), .ZN(n508) );
  XOR2_X1 U626 ( .A(G101), .B(G104), .Z(n511) );
  XNOR2_X1 U627 ( .A(G107), .B(G110), .ZN(n510) );
  NAND2_X1 U628 ( .A1(G227), .A2(n403), .ZN(n515) );
  XOR2_X1 U629 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n518) );
  XNOR2_X1 U630 ( .A(KEYINPUT72), .B(G469), .ZN(n517) );
  XNOR2_X1 U631 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X2 U632 ( .A(n520), .B(n519), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n525), .A2(n626), .ZN(n527) );
  NAND2_X1 U634 ( .A1(G210), .A2(n528), .ZN(n526) );
  NAND2_X1 U635 ( .A1(G214), .A2(n528), .ZN(n691) );
  NAND2_X1 U636 ( .A1(n557), .A2(n691), .ZN(n530) );
  INV_X1 U637 ( .A(n594), .ZN(n531) );
  XNOR2_X1 U638 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n544) );
  XOR2_X1 U639 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n534) );
  NAND2_X1 U640 ( .A1(n532), .A2(G214), .ZN(n533) );
  XNOR2_X1 U641 ( .A(n534), .B(n533), .ZN(n542) );
  XNOR2_X1 U642 ( .A(n536), .B(n535), .ZN(n540) );
  XNOR2_X1 U643 ( .A(G143), .B(G140), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n537), .B(n538), .ZN(n539) );
  XOR2_X1 U645 ( .A(n540), .B(n539), .Z(n541) );
  NOR2_X1 U646 ( .A1(G902), .A2(n714), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n544), .B(n543), .ZN(n545) );
  NOR2_X1 U648 ( .A1(n572), .A2(n546), .ZN(n657) );
  AND2_X1 U649 ( .A1(n572), .A2(n546), .ZN(n659) );
  XNOR2_X1 U650 ( .A(KEYINPUT100), .B(n659), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n657), .A2(n584), .ZN(n695) );
  NAND2_X1 U652 ( .A1(n695), .A2(KEYINPUT47), .ZN(n547) );
  NAND2_X1 U653 ( .A1(n463), .A2(n547), .ZN(n559) );
  XOR2_X1 U654 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n549) );
  INV_X1 U655 ( .A(n614), .ZN(n684) );
  NAND2_X1 U656 ( .A1(n684), .A2(n691), .ZN(n548) );
  XNOR2_X1 U657 ( .A(n549), .B(n548), .ZN(n556) );
  NAND2_X1 U658 ( .A1(n674), .A2(n673), .ZN(n676) );
  INV_X1 U659 ( .A(KEYINPUT107), .ZN(n550) );
  XNOR2_X1 U660 ( .A(n617), .B(n550), .ZN(n553) );
  NAND2_X1 U661 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U662 ( .A1(n573), .A2(n572), .ZN(n598) );
  XNOR2_X1 U663 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n561) );
  NOR2_X1 U664 ( .A1(n695), .A2(n650), .ZN(n560) );
  NAND2_X1 U665 ( .A1(n561), .A2(n560), .ZN(n568) );
  XOR2_X1 U666 ( .A(n614), .B(KEYINPUT6), .Z(n606) );
  NOR2_X1 U667 ( .A1(n562), .A2(n606), .ZN(n563) );
  AND2_X1 U668 ( .A1(n563), .A2(n691), .ZN(n564) );
  NAND2_X1 U669 ( .A1(n657), .A2(n564), .ZN(n580) );
  NOR2_X1 U670 ( .A1(n570), .A2(n580), .ZN(n565) );
  XNOR2_X1 U671 ( .A(KEYINPUT36), .B(n565), .ZN(n567) );
  NAND2_X1 U672 ( .A1(n567), .A2(n601), .ZN(n663) );
  NAND2_X1 U673 ( .A1(n573), .A2(n572), .ZN(n694) );
  INV_X1 U674 ( .A(n694), .ZN(n574) );
  NAND2_X1 U675 ( .A1(n697), .A2(n574), .ZN(n575) );
  XOR2_X1 U676 ( .A(n575), .B(KEYINPUT41), .Z(n707) );
  INV_X1 U677 ( .A(n707), .ZN(n688) );
  INV_X1 U678 ( .A(n580), .ZN(n581) );
  NAND2_X1 U679 ( .A1(n677), .A2(n581), .ZN(n582) );
  XOR2_X1 U680 ( .A(KEYINPUT43), .B(n582), .Z(n583) );
  NOR2_X1 U681 ( .A1(n557), .A2(n583), .ZN(n665) );
  NAND2_X1 U682 ( .A1(n585), .A2(n584), .ZN(n664) );
  INV_X1 U683 ( .A(G898), .ZN(n730) );
  NAND2_X1 U684 ( .A1(n409), .A2(n730), .ZN(n725) );
  NOR2_X1 U685 ( .A1(n590), .A2(n725), .ZN(n591) );
  NOR2_X1 U686 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U687 ( .A(n616), .ZN(n596) );
  XNOR2_X1 U688 ( .A(n597), .B(KEYINPUT34), .ZN(n599) );
  AND2_X1 U689 ( .A1(n613), .A2(n601), .ZN(n602) );
  XNOR2_X1 U690 ( .A(KEYINPUT104), .B(n602), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n603), .A2(n694), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n605), .B(KEYINPUT22), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n613), .A2(n677), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n611), .A2(n614), .ZN(n649) );
  NAND2_X1 U696 ( .A1(n750), .A2(n649), .ZN(n612) );
  NAND2_X1 U697 ( .A1(n686), .A2(n616), .ZN(n615) );
  XNOR2_X1 U698 ( .A(n615), .B(KEYINPUT31), .ZN(n660) );
  NAND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U700 ( .A1(n684), .A2(n618), .ZN(n645) );
  NOR2_X1 U701 ( .A1(n660), .A2(n645), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n695), .A2(n619), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n622), .B(n623), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n625), .B(KEYINPUT120), .ZN(G63) );
  XOR2_X1 U705 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n628) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT86), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n630), .B(n629), .ZN(n631) );
  INV_X1 U708 ( .A(KEYINPUT119), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT56), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(G51) );
  XOR2_X1 U711 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n635) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(n639) );
  INV_X1 U713 ( .A(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G57) );
  XOR2_X1 U715 ( .A(G101), .B(n642), .Z(n643) );
  XNOR2_X1 U716 ( .A(KEYINPUT112), .B(n643), .ZN(G3) );
  NAND2_X1 U717 ( .A1(n645), .A2(n657), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(G104), .ZN(G6) );
  XOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n647) );
  NAND2_X1 U720 ( .A1(n645), .A2(n659), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U722 ( .A(G107), .B(n648), .ZN(G9) );
  XNOR2_X1 U723 ( .A(G110), .B(n649), .ZN(G12) );
  XOR2_X1 U724 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n652) );
  INV_X1 U725 ( .A(n650), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n654), .A2(n659), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U728 ( .A(G128), .B(n653), .Z(G30) );
  XOR2_X1 U729 ( .A(n354), .B(G143), .Z(G45) );
  NAND2_X1 U730 ( .A1(n654), .A2(n657), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n655), .B(KEYINPUT114), .ZN(n656) );
  XNOR2_X1 U732 ( .A(G146), .B(n656), .ZN(G48) );
  NAND2_X1 U733 ( .A1(n660), .A2(n657), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n658), .B(G113), .ZN(G15) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(G116), .ZN(G18) );
  XOR2_X1 U737 ( .A(G125), .B(KEYINPUT37), .Z(n662) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(G27) );
  XNOR2_X1 U739 ( .A(G134), .B(n664), .ZN(G36) );
  XOR2_X1 U740 ( .A(G140), .B(n665), .Z(G42) );
  NAND2_X1 U741 ( .A1(n426), .A2(n402), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(KEYINPUT84), .ZN(n669) );
  NAND2_X1 U743 ( .A1(KEYINPUT2), .A2(n667), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n671) );
  AND2_X1 U745 ( .A1(n426), .A2(n743), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n674), .A2(n437), .ZN(n675) );
  XNOR2_X1 U748 ( .A(KEYINPUT49), .B(n675), .ZN(n682) );
  XOR2_X1 U749 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n679) );
  NAND2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U752 ( .A(KEYINPUT115), .B(n680), .ZN(n681) );
  NAND2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U756 ( .A(KEYINPUT51), .B(n687), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n690), .B(KEYINPUT117), .ZN(n703) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n700) );
  INV_X1 U761 ( .A(n695), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U763 ( .A(KEYINPUT118), .B(n698), .Z(n699) );
  NOR2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n708), .A2(n701), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  XNOR2_X1 U772 ( .A(n718), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U773 ( .A(n719), .B(KEYINPUT121), .Z(n721) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n723), .A2(n722), .ZN(G66) );
  NAND2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n735) );
  XOR2_X1 U777 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n727) );
  NAND2_X1 U778 ( .A1(G224), .A2(n409), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U780 ( .A(KEYINPUT122), .B(n728), .Z(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n733) );
  NOR2_X1 U782 ( .A1(n409), .A2(n402), .ZN(n732) );
  NOR2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(G69) );
  XOR2_X1 U785 ( .A(n737), .B(n736), .Z(n738) );
  XNOR2_X1 U786 ( .A(KEYINPUT124), .B(n738), .ZN(n742) );
  XNOR2_X1 U787 ( .A(KEYINPUT125), .B(n742), .ZN(n739) );
  XNOR2_X1 U788 ( .A(G227), .B(n739), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(n409), .ZN(n747) );
  XOR2_X1 U791 ( .A(n743), .B(n742), .Z(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(n403), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n747), .A2(n746), .ZN(G72) );
  XOR2_X1 U794 ( .A(n748), .B(G122), .Z(n749) );
  XNOR2_X1 U795 ( .A(KEYINPUT126), .B(n749), .ZN(G24) );
  XOR2_X1 U796 ( .A(n750), .B(G119), .Z(n751) );
  XNOR2_X1 U797 ( .A(KEYINPUT127), .B(n751), .ZN(G21) );
  XOR2_X1 U798 ( .A(G137), .B(n752), .Z(G39) );
  XOR2_X1 U799 ( .A(G131), .B(n753), .Z(G33) );
endmodule

