//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G128), .B(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT13), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n188), .B(G134), .C1(KEYINPUT13), .C2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G122), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G122), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(KEYINPUT96), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(KEYINPUT96), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(G107), .B1(new_n199), .B2(new_n200), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n191), .B(new_n193), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n196), .A2(G122), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(KEYINPUT14), .B2(new_n197), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n207), .B(KEYINPUT97), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n197), .A2(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g023(.A(G107), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n204), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n187), .B(new_n192), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT9), .B(G234), .Z(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G217), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n216), .A2(new_n217), .A3(G953), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT98), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n205), .A2(new_n213), .A3(new_n218), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G902), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n205), .A2(new_n213), .A3(KEYINPUT98), .A4(new_n218), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n223), .A2(KEYINPUT99), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G478), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT15), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n226), .A2(new_n228), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G475), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n189), .ZN(new_n234));
  NOR2_X1   g048(.A1(G237), .A2(G953), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(G214), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G237), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G214), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT92), .A2(G143), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT17), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n240), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n234), .A2(G214), .A3(new_n235), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n243), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT94), .ZN(new_n249));
  INV_X1    g063(.A(G125), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n250), .A2(KEYINPUT16), .A3(G140), .ZN(new_n251));
  XNOR2_X1  g065(.A(G125), .B(G140), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(KEYINPUT16), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n244), .A2(new_n245), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT17), .A3(G131), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT94), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n242), .A2(new_n258), .A3(new_n243), .A4(new_n247), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n249), .A2(new_n255), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G113), .B(G122), .ZN(new_n261));
  INV_X1    g075(.A(G104), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT78), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(new_n264), .A3(new_n254), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n252), .B2(new_n254), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n266), .A2(new_n267), .B1(new_n254), .B2(new_n252), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT18), .A2(G131), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n256), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n272));
  INV_X1    g086(.A(new_n256), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n269), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n256), .A2(KEYINPUT93), .A3(new_n270), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n268), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n260), .A2(new_n263), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT95), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT95), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n260), .A2(new_n279), .A3(new_n263), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n260), .A2(new_n276), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n263), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n232), .B1(new_n283), .B2(new_n224), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n263), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n242), .A2(new_n247), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n253), .A2(G146), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n252), .B(KEYINPUT19), .Z(new_n289));
  OAI211_X1 g103(.A(new_n287), .B(new_n288), .C1(new_n289), .C2(G146), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n276), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n278), .A2(new_n280), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n292), .A2(G475), .A3(G902), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n286), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n281), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n294), .A3(new_n232), .A4(new_n224), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n231), .B(new_n285), .C1(new_n295), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT11), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n192), .B2(G137), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT66), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n192), .A2(G137), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT11), .ZN(new_n306));
  INV_X1    g120(.A(G137), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G134), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n310), .B(new_n302), .C1(new_n192), .C2(G137), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n304), .A2(new_n306), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n303), .B2(KEYINPUT66), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n314), .A2(new_n246), .A3(new_n306), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n262), .B2(G107), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n202), .A2(KEYINPUT3), .A3(G104), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n319), .B1(new_n262), .B2(G107), .ZN(new_n320));
  INV_X1    g134(.A(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n202), .B2(G104), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n202), .A2(G104), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n323), .A2(new_n202), .A3(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(G101), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n254), .A2(G143), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n189), .A2(G146), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT1), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .A4(G128), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n330), .A2(new_n331), .ZN(new_n334));
  INV_X1    g148(.A(G128), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n189), .A2(G146), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT64), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n254), .B2(G143), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n189), .A2(KEYINPUT64), .A3(G146), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n333), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n329), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n316), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT12), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n238), .A2(G227), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(G140), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT82), .B(G110), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n320), .A2(new_n321), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n353));
  OR3_X1    g167(.A1(new_n320), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n189), .A2(KEYINPUT64), .A3(G146), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT64), .B1(new_n189), .B2(G146), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n330), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G128), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT0), .A4(G128), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n355), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n355), .B(new_n362), .C1(new_n343), .C2(new_n359), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n353), .B(new_n354), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT70), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n344), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT70), .B(new_n333), .C1(new_n343), .C2(new_n336), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT10), .A3(new_n329), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n329), .A2(new_n337), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n316), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n366), .A2(new_n371), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT12), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n316), .C1(new_n338), .C2(new_n345), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n347), .A2(new_n351), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n379), .A2(KEYINPUT85), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n371), .A3(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n316), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(new_n351), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(KEYINPUT85), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n224), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n347), .A2(new_n376), .A3(new_n378), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n347), .A2(KEYINPUT84), .A3(new_n376), .A4(new_n378), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n351), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n382), .B2(new_n376), .ZN(new_n395));
  OAI21_X1  g209(.A(G469), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(G469), .A2(G902), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G221), .B1(new_n216), .B2(G902), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT101), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n402), .B(KEYINPUT86), .Z(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n404));
  INV_X1    g218(.A(G119), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(G116), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(KEYINPUT88), .A3(G116), .A4(new_n405), .ZN(new_n409));
  XNOR2_X1  g223(.A(G116), .B(G119), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n408), .A2(G113), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n410), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT2), .B(G113), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n329), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n408), .A2(G113), .A3(new_n409), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n410), .A2(KEYINPUT68), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n410), .A2(KEYINPUT68), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n420), .A2(new_n421), .A3(new_n404), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n415), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n329), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n412), .A2(new_n329), .A3(KEYINPUT90), .A4(new_n415), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(G110), .B(G122), .Z(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT8), .Z(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n415), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n353), .A2(new_n432), .A3(new_n354), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n329), .B(new_n415), .C1(new_n419), .C2(new_n422), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n428), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n362), .B1(new_n343), .B2(new_n359), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G125), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(G125), .B2(new_n344), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n238), .A2(G224), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT7), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n440), .A2(new_n442), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n430), .A2(new_n437), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n435), .A2(new_n428), .B1(KEYINPUT89), .B2(KEYINPUT6), .ZN(new_n448));
  INV_X1    g262(.A(new_n428), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT89), .A2(KEYINPUT6), .ZN(new_n450));
  AOI211_X1 g264(.A(new_n449), .B(new_n450), .C1(new_n433), .C2(new_n434), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n448), .A2(new_n451), .A3(new_n436), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n440), .B(new_n441), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n447), .B(new_n224), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n435), .A2(new_n428), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n450), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n435), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n428), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n437), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n453), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n455), .A3(new_n447), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n403), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(G234), .A2(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(G902), .A3(G953), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT100), .Z(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(G898), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n466), .A2(G952), .A3(new_n238), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n301), .A2(new_n400), .A3(new_n401), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT65), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n438), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT65), .B(new_n362), .C1(new_n343), .C2(new_n359), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(new_n375), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n308), .B2(new_n305), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n315), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n344), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n316), .A2(KEYINPUT67), .A3(new_n479), .A4(new_n480), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n484), .B1(new_n368), .B2(new_n369), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n438), .A2(KEYINPUT69), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n492), .A2(new_n364), .B1(new_n313), .B2(new_n315), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n491), .A2(new_n493), .A3(new_n489), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n490), .A2(new_n432), .A3(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n491), .A2(new_n493), .A3(new_n432), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n235), .A2(G210), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n321), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n501), .B(new_n502), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n491), .B2(new_n493), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n370), .A2(new_n485), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n316), .B1(new_n363), .B2(new_n365), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT73), .ZN(new_n510));
  INV_X1    g324(.A(new_n432), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n497), .B1(new_n488), .B2(new_n432), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n505), .B1(new_n504), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n432), .B1(new_n491), .B2(new_n493), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n498), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n514), .B1(new_n520), .B2(new_n513), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n503), .A2(KEYINPUT29), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n517), .B(new_n224), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G472), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n516), .A2(KEYINPUT74), .A3(new_n504), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT74), .B1(new_n516), .B2(new_n504), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n494), .B1(new_n488), .B2(new_n489), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n497), .B1(new_n530), .B2(new_n432), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n531), .B2(new_n503), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n534));
  NAND4_X1  g348(.A1(new_n496), .A2(new_n498), .A3(new_n503), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT72), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n531), .A2(new_n537), .A3(new_n503), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT32), .B(new_n526), .C1(new_n533), .C2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n516), .A2(new_n504), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT74), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT31), .B1(new_n499), .B2(new_n504), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n516), .A2(KEYINPUT74), .A3(new_n504), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n539), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(new_n547), .B2(new_n525), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n524), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G119), .B(G128), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT75), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT24), .B(G110), .Z(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT76), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n405), .B2(G128), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n557), .A2(KEYINPUT23), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(KEYINPUT23), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n559), .C1(G119), .C2(new_n335), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n255), .B1(G110), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(G110), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n551), .A2(new_n552), .ZN(new_n564));
  OAI221_X1 g378(.A(new_n288), .B1(new_n266), .B2(new_n267), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G137), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n562), .A2(new_n570), .A3(new_n565), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n224), .A3(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n217), .B1(G234), .B2(new_n224), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n572), .A2(new_n573), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n577), .A2(G902), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT81), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n398), .A2(new_n399), .A3(new_n465), .A4(new_n473), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT101), .B1(new_n586), .B2(new_n300), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n476), .A2(new_n549), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(new_n539), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n224), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n547), .A2(new_n525), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n584), .ZN(new_n597));
  INV_X1    g411(.A(new_n586), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n285), .B1(new_n295), .B2(new_n299), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n227), .ZN(new_n601));
  INV_X1    g415(.A(new_n222), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n602), .A2(KEYINPUT103), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(KEYINPUT103), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(KEYINPUT33), .A3(new_n220), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT102), .B(KEYINPUT33), .Z(new_n606));
  NAND3_X1  g420(.A1(new_n223), .A2(new_n225), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n224), .A2(G478), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n599), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n597), .A2(new_n598), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n293), .A2(new_n616), .A3(new_n294), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n297), .A2(new_n232), .A3(new_n224), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT104), .B1(new_n618), .B2(KEYINPUT20), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT105), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n298), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n292), .A2(G475), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT105), .A3(new_n294), .A4(new_n224), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n284), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n231), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n597), .A2(new_n598), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n571), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n566), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n581), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n578), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n533), .B2(new_n539), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n594), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT106), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n593), .A2(new_n640), .A3(new_n594), .A4(new_n635), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n639), .A2(new_n476), .A3(new_n641), .A4(new_n587), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G110), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AND3_X1   g459(.A1(new_n398), .A2(new_n399), .A3(new_n465), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n549), .A2(new_n635), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n616), .B1(new_n293), .B2(new_n294), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n618), .A2(KEYINPUT104), .A3(KEYINPUT20), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n622), .A4(new_n624), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n471), .B1(new_n468), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n627), .A2(new_n650), .A3(new_n285), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n335), .ZN(G30));
  AND2_X1   g472(.A1(new_n457), .A2(new_n464), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT109), .B(KEYINPUT38), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n403), .ZN(new_n663));
  INV_X1    g477(.A(new_n599), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n231), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n652), .B(KEYINPUT39), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n400), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT111), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n666), .B1(new_n670), .B2(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n594), .A2(KEYINPUT32), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n547), .A2(new_n541), .A3(new_n525), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n531), .A2(new_n504), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n224), .B1(new_n519), .B2(new_n503), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n635), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n671), .B(new_n680), .C1(KEYINPUT40), .C2(new_n670), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  NOR2_X1   g496(.A1(new_n611), .A2(new_n652), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n549), .A2(new_n635), .A3(new_n646), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT112), .B(G146), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G48));
  NAND2_X1  g500(.A1(new_n387), .A2(new_n224), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n399), .A3(new_n389), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n474), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n549), .A2(new_n585), .A3(new_n612), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n549), .A2(new_n585), .A3(new_n628), .A4(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND4_X1  g509(.A1(new_n549), .A2(new_n301), .A3(new_n635), .A4(new_n690), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AOI22_X1  g511(.A1(new_n536), .A2(new_n538), .B1(new_n521), .B2(new_n504), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n526), .B1(new_n698), .B2(new_n545), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT113), .B(G472), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n699), .B1(new_n592), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n583), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n689), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n703), .A2(new_n475), .A3(new_n665), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  INV_X1    g520(.A(new_n465), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n701), .A2(new_n635), .A3(new_n683), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n396), .A2(KEYINPUT114), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n713), .B(G469), .C1(new_n394), .C2(new_n395), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n389), .A3(new_n397), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n399), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n403), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n659), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n549), .A2(new_n585), .A3(new_n683), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n718), .A2(new_n611), .A3(new_n652), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n549), .A4(new_n702), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n711), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n722), .A2(new_n711), .A3(new_n724), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NAND3_X1  g543(.A1(new_n549), .A2(new_n585), .A3(new_n719), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(new_n656), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  INV_X1    g546(.A(new_n389), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n394), .A2(new_n395), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(KEYINPUT45), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n397), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n733), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(KEYINPUT46), .A3(new_n397), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n716), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n668), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n664), .A2(new_n610), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n744), .B2(KEYINPUT116), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(KEYINPUT116), .A3(KEYINPUT43), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT44), .A3(new_n596), .A4(new_n635), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n596), .A2(new_n635), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n748), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n457), .A2(new_n663), .A3(new_n464), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n743), .A2(new_n750), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(new_n549), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n584), .A2(new_n683), .A3(new_n754), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  AOI211_X1 g574(.A(new_n760), .B(new_n716), .C1(new_n740), .C2(new_n741), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  NOR2_X1   g577(.A1(new_n759), .A2(new_n761), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n688), .A2(new_n716), .A3(new_n389), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n703), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n748), .A3(new_n472), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n754), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n689), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n748), .A2(new_n472), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n662), .A2(new_n663), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n704), .A2(new_n754), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT120), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n584), .A2(new_n472), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(new_n679), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n599), .A2(new_n610), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n771), .A2(new_n776), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n701), .A2(new_n635), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n773), .A2(KEYINPUT50), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n769), .A2(new_n782), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n786), .A2(new_n774), .A3(new_n781), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(KEYINPUT51), .A3(new_n785), .A4(new_n769), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n757), .A2(new_n583), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT48), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT121), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(KEYINPUT121), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n792), .A2(new_n783), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n770), .A2(new_n771), .A3(new_n465), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(G952), .A3(new_n238), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n794), .B1(new_n783), .B2(new_n792), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n789), .A2(new_n791), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n684), .B(new_n709), .C1(new_n647), .C2(new_n656), .ZN(new_n802));
  INV_X1    g616(.A(new_n635), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n652), .A2(new_n716), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n715), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n664), .A2(new_n707), .A3(new_n231), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n678), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT52), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n803), .B1(new_n674), .B2(new_n524), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n654), .B(KEYINPUT108), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n812), .B(new_n646), .C1(new_n813), .C2(new_n683), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n678), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n709), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n705), .A2(new_n694), .A3(new_n691), .A4(new_n696), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n229), .A2(new_n230), .A3(new_n652), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n626), .A2(KEYINPUT117), .A3(new_n754), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n650), .A2(new_n754), .A3(new_n821), .A4(new_n285), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n549), .A3(new_n400), .A4(new_n635), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n611), .B1(new_n599), .B2(new_n231), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n595), .A2(new_n585), .A3(new_n598), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n642), .A3(new_n588), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n784), .A2(new_n683), .A3(new_n719), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n730), .B2(new_n656), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n722), .B2(new_n724), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n818), .A2(new_n820), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n811), .A3(new_n817), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n722), .A2(new_n711), .A3(new_n724), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n820), .B1(new_n838), .B2(new_n725), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n833), .A2(new_n811), .A3(new_n817), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n819), .B1(new_n726), .B2(new_n727), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT53), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n837), .A2(new_n839), .A3(new_n834), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT119), .B1(new_n847), .B2(new_n841), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(KEYINPUT54), .C1(new_n845), .C2(new_n846), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n801), .A2(new_n842), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n778), .A2(new_n612), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n851), .A2(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n688), .A2(new_n389), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n702), .A3(new_n717), .A4(new_n856), .ZN(new_n857));
  OR4_X1    g671(.A1(new_n678), .A2(new_n857), .A3(new_n662), .A4(new_n744), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n858), .ZN(G75));
  INV_X1    g673(.A(new_n835), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n837), .A2(new_n819), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n845), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n224), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n461), .B(new_n453), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n866), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n238), .A2(G952), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G51));
  XOR2_X1   g684(.A(new_n397), .B(KEYINPUT57), .Z(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n845), .B2(new_n861), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n842), .ZN(new_n874));
  INV_X1    g688(.A(new_n387), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT122), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OR3_X1    g690(.A1(new_n862), .A2(new_n224), .A3(new_n737), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n841), .B1(new_n836), .B2(new_n840), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n387), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n869), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(G54));
  NAND3_X1  g699(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n292), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n292), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n869), .ZN(G60));
  NAND3_X1  g703(.A1(new_n848), .A2(new_n842), .A3(new_n850), .ZN(new_n890));
  NAND2_X1  g704(.A1(G478), .A2(G902), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT59), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n890), .A2(new_n893), .B1(new_n605), .B2(new_n607), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n608), .B(new_n892), .C1(new_n873), .C2(new_n842), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n869), .A3(new_n895), .ZN(G63));
  NAND2_X1  g710(.A1(G217), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT60), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n862), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n579), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n869), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n862), .A2(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n633), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n901), .B(new_n903), .C1(new_n904), .C2(KEYINPUT61), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n904), .B(new_n884), .C1(new_n902), .C2(new_n579), .ZN(new_n907));
  INV_X1    g721(.A(new_n903), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n884), .B1(new_n902), .B2(new_n579), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(G66));
  INV_X1    g725(.A(G224), .ZN(new_n912));
  OAI21_X1  g726(.A(G953), .B1(new_n469), .B2(new_n912), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n588), .A2(new_n820), .A3(new_n642), .A4(new_n829), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n452), .B1(G898), .B2(new_n238), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(G69));
  XOR2_X1   g731(.A(KEYINPUT124), .B(KEYINPUT125), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n289), .B(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n530), .B(new_n919), .Z(new_n920));
  INV_X1    g734(.A(new_n802), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n681), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n754), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n670), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n926), .A2(new_n549), .A3(new_n585), .A4(new_n828), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n755), .A2(new_n762), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n920), .B1(new_n929), .B2(G953), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n931));
  INV_X1    g745(.A(new_n920), .ZN(new_n932));
  NAND2_X1  g746(.A1(G900), .A2(G953), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n743), .A2(new_n792), .A3(new_n809), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n731), .A2(new_n755), .A3(new_n762), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n728), .A3(new_n921), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n932), .B(new_n933), .C1(new_n936), .C2(G953), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n930), .A2(new_n931), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n238), .B1(G227), .B2(G900), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n930), .A2(new_n931), .A3(new_n941), .A4(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(G72));
  INV_X1    g757(.A(new_n675), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n924), .A2(new_n914), .A3(new_n927), .A4(new_n928), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n531), .B(new_n504), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n847), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n935), .A2(new_n728), .A3(new_n921), .A4(new_n914), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n499), .B(new_n503), .C1(new_n953), .C2(new_n947), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n954), .B2(new_n869), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n947), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n531), .A3(new_n504), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(KEYINPUT127), .A3(new_n884), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n948), .B(new_n951), .C1(new_n955), .C2(new_n958), .ZN(G57));
endmodule


