//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n467), .A3(G2104), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n475), .A2(new_n464), .A3(new_n466), .A4(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n475), .A2(G2105), .A3(new_n466), .A4(new_n477), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n464), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n478), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(G136), .B2(new_n487), .ZN(G162));
  AND4_X1   g063(.A1(G2105), .A2(new_n475), .A3(new_n466), .A4(new_n477), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n464), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n491), .A2(new_n492), .A3(new_n490), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n489), .A2(G126), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n464), .A2(G138), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n475), .A2(new_n466), .A3(new_n477), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n466), .A2(new_n468), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n469), .A2(new_n503), .A3(new_n499), .A4(new_n496), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n498), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n495), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n495), .B2(new_n505), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(G164));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n511), .A2(new_n510), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n519), .A2(G543), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(G651), .B1(new_n529), .B2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(new_n516), .A2(KEYINPUT73), .A3(new_n517), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n534), .B1(new_n511), .B2(new_n510), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n515), .A2(G89), .A3(new_n521), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n529), .A2(G51), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND3_X1  g118(.A1(new_n515), .A2(G90), .A3(new_n521), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n529), .A2(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n533), .A2(new_n535), .A3(G64), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(G171));
  NAND3_X1  g126(.A1(new_n515), .A2(G81), .A3(new_n521), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n529), .A2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n533), .A2(new_n535), .A3(G56), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n547), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(new_n553), .A4(new_n552), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND3_X1  g144(.A1(new_n515), .A2(G91), .A3(new_n521), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n515), .A2(KEYINPUT78), .A3(G91), .A4(new_n521), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n547), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  AND2_X1   g153(.A1(G53), .A2(G543), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n578), .B(new_n579), .C1(new_n512), .C2(new_n513), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n579), .B1(KEYINPUT75), .B2(new_n583), .C1(new_n512), .C2(new_n513), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n583), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n582), .A2(new_n584), .B1(new_n583), .B2(new_n580), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT77), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n574), .A2(new_n577), .A3(new_n589), .A4(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  NAND2_X1  g168(.A1(new_n522), .A2(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n529), .A2(G49), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n526), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n529), .A2(G48), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n522), .A2(KEYINPUT79), .A3(G86), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n515), .A2(G86), .A3(new_n521), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n603), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G305));
  NAND2_X1  g184(.A1(new_n536), .A2(G60), .ZN(new_n610));
  NAND2_X1  g185(.A1(G72), .A2(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n529), .A2(G47), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n522), .A2(G85), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n547), .B1(new_n610), .B2(new_n611), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n515), .A2(new_n521), .ZN(new_n619));
  INV_X1    g194(.A(G85), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT80), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(G290));
  NAND2_X1  g198(.A1(G301), .A2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(G79), .A2(G543), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n526), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G651), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n529), .A2(G54), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n515), .A2(G92), .A3(new_n521), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .A4(new_n521), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n624), .B1(G868), .B2(new_n635), .ZN(G284));
  XNOR2_X1  g211(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g212(.A1(G286), .A2(G868), .ZN(new_n638));
  INV_X1    g213(.A(G299), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(G868), .ZN(G297));
  OAI21_X1  g215(.A(new_n638), .B1(new_n639), .B2(G868), .ZN(G280));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n635), .B1(new_n642), .B2(G860), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT82), .Z(G148));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n642), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G868), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n564), .B2(G868), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n469), .A2(new_n473), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  OAI21_X1  g228(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n655));
  INV_X1    g230(.A(G111), .ZN(new_n656));
  AOI22_X1  g231(.A1(new_n654), .A2(new_n655), .B1(new_n656), .B2(G2105), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n655), .B2(new_n654), .ZN(new_n658));
  INV_X1    g233(.A(G135), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n478), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n489), .B2(G123), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n489), .A2(new_n661), .A3(G123), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(G2096), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(G2096), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n653), .A2(new_n667), .A3(new_n668), .ZN(G156));
  XNOR2_X1  g244(.A(G2427), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT14), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1341), .B(G1348), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2451), .B(G2454), .Z(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n683), .A2(G14), .A3(new_n684), .ZN(G401));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT17), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2084), .B(G2090), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n687), .B2(new_n689), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n688), .B2(new_n689), .ZN(new_n693));
  INV_X1    g268(.A(new_n689), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(new_n690), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT18), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n691), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G2100), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT88), .B(G2096), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G227));
  XNOR2_X1  g276(.A(G1971), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1961), .B(G1966), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT89), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1956), .B(G2474), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT20), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n706), .A2(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n713), .C1(new_n703), .C2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XOR2_X1   g290(.A(G1981), .B(G1986), .Z(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n715), .B(new_n720), .ZN(G229));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G28), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n723), .B2(G28), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n722), .B1(new_n724), .B2(new_n726), .C1(new_n666), .C2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(G168), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(G21), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n725), .A2(G33), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  INV_X1    g311(.A(G139), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n736), .B1(new_n737), .B2(new_n478), .C1(new_n738), .C2(new_n464), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2072), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n732), .A2(new_n733), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n728), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n728), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n727), .B(new_n743), .C1(G1961), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n725), .A2(G27), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT101), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n725), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n725), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n745), .A2(G1961), .B1(G2084), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G2084), .B2(new_n756), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n740), .A2(new_n741), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT97), .Z(new_n760));
  NAND4_X1  g335(.A1(new_n746), .A2(new_n751), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n725), .A2(G32), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n489), .A2(G129), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT99), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n473), .A2(G105), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n487), .A2(G141), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT98), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(new_n725), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT27), .ZN(new_n775));
  INV_X1    g350(.A(G1996), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n761), .A2(new_n777), .A3(KEYINPUT102), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n728), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n564), .B2(new_n728), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1341), .Z(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n635), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT94), .B(G1348), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G35), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G162), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT29), .B(G2090), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n781), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n725), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n487), .A2(G140), .ZN(new_n794));
  OR2_X1    g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n796));
  INV_X1    g371(.A(G128), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n482), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(new_n725), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  INV_X1    g377(.A(G2067), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n728), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1956), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n778), .A2(new_n790), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n728), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n728), .B2(G23), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT92), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n728), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n728), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(G1971), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(G1971), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n818), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n728), .A2(G6), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n608), .B2(new_n728), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT32), .B(G1981), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n824), .A2(KEYINPUT34), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT34), .B1(new_n824), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n728), .A2(G24), .ZN(new_n831));
  INV_X1    g406(.A(G290), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n728), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(G1986), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(G1986), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n725), .A2(G25), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n487), .A2(G131), .ZN(new_n837));
  INV_X1    g412(.A(G119), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n464), .A2(G107), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n482), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n836), .B1(new_n843), .B2(new_n725), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT35), .B(G1991), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT91), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n834), .A2(new_n835), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n829), .A2(new_n830), .A3(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT102), .B1(new_n761), .B2(new_n777), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n811), .A2(new_n851), .A3(new_n852), .ZN(G150));
  INV_X1    g428(.A(G150), .ZN(G311));
  NAND3_X1  g429(.A1(new_n515), .A2(G93), .A3(new_n521), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n529), .A2(G55), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n533), .A2(new_n535), .A3(G67), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n547), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G860), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n858), .A2(new_n859), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n856), .B(new_n855), .C1(new_n865), .C2(new_n547), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n563), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n560), .A2(new_n553), .A3(new_n552), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n635), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT104), .Z(new_n877));
  OAI21_X1  g452(.A(new_n862), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n864), .B1(new_n877), .B2(new_n878), .ZN(G145));
  XNOR2_X1  g454(.A(G162), .B(G160), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n666), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n495), .A2(new_n505), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n799), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n773), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n739), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n772), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n739), .A2(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(G106), .A2(G2105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n894));
  INV_X1    g469(.A(G142), .ZN(new_n895));
  INV_X1    g470(.A(G130), .ZN(new_n896));
  OAI221_X1 g471(.A(new_n894), .B1(new_n478), .B2(new_n895), .C1(new_n896), .C2(new_n482), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT106), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n651), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n843), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n884), .A2(new_n890), .A3(new_n888), .A4(new_n886), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n892), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n881), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  INV_X1    g481(.A(new_n881), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT107), .A4(new_n909), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT40), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(G395));
  XOR2_X1   g491(.A(new_n871), .B(new_n645), .Z(new_n917));
  AOI21_X1  g492(.A(new_n576), .B1(new_n572), .B2(new_n573), .ZN(new_n918));
  AOI221_X4 g493(.A(new_n588), .B1(new_n580), .B2(new_n583), .C1(new_n582), .C2(new_n584), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT77), .B1(new_n585), .B2(new_n586), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n918), .A2(new_n921), .A3(new_n635), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n635), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(new_n635), .ZN(new_n926));
  NAND2_X1  g501(.A1(G299), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n918), .A2(new_n921), .A3(new_n635), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n922), .A2(new_n923), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(KEYINPUT108), .A3(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n917), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n917), .A2(new_n932), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT42), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n524), .A2(KEYINPUT109), .A3(new_n530), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT109), .B1(new_n524), .B2(new_n530), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G290), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n617), .B(new_n622), .C1(new_n938), .C2(new_n939), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G305), .A2(new_n812), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n608), .A2(G288), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n941), .A2(new_n944), .A3(new_n945), .A4(new_n942), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT42), .B1(new_n935), .B2(new_n936), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n937), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n937), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g528(.A(G868), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G868), .B2(new_n861), .ZN(G295));
  OAI21_X1  g530(.A(new_n954), .B1(G868), .B2(new_n861), .ZN(G331));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n546), .B2(new_n550), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n548), .A2(new_n549), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G651), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT110), .A3(new_n545), .A4(new_n544), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G168), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(G286), .A3(new_n961), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n867), .A2(new_n963), .A3(new_n870), .A4(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n958), .A2(G286), .A3(new_n961), .ZN(new_n966));
  AOI21_X1  g541(.A(G286), .B1(new_n958), .B2(new_n961), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n861), .B1(new_n558), .B2(new_n562), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n966), .A2(new_n967), .B1(new_n968), .B2(new_n869), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n931), .A2(new_n933), .A3(new_n965), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n927), .A2(new_n929), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n965), .B2(new_n969), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n949), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n970), .A2(new_n949), .A3(new_n973), .A4(KEYINPUT111), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n970), .A2(new_n973), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n979), .B2(new_n950), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n924), .A2(new_n930), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n965), .A2(new_n969), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n972), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n909), .B1(new_n985), .B2(new_n949), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n982), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n992), .A3(KEYINPUT43), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n986), .B1(new_n976), .B2(new_n977), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT112), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n978), .A2(new_n995), .A3(new_n980), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n999), .A2(KEYINPUT44), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n997), .B2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n991), .B1(new_n1001), .B2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n882), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT114), .B(G40), .Z(new_n1007));
  NOR3_X1   g582(.A1(new_n472), .A2(new_n480), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n772), .A2(G1996), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n799), .B(new_n803), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n772), .B2(G1996), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1013), .B(new_n1014), .C1(new_n1010), .C2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n842), .B(new_n846), .Z(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(G290), .A2(G1986), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G290), .A2(G1986), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1009), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT45), .B(new_n1004), .C1(new_n507), .C2(new_n508), .ZN(new_n1025));
  OR3_X1    g600(.A1(new_n472), .A2(new_n480), .A3(new_n1007), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1028), .B2(G1966), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1008), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1004), .B1(new_n507), .B2(new_n508), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(KEYINPUT50), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1966), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT117), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1029), .A2(new_n1034), .A3(new_n1036), .A4(G168), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1033), .A2(new_n1032), .B1(new_n1035), .B2(KEYINPUT117), .ZN(new_n1039));
  AOI21_X1  g614(.A(G168), .B1(new_n1039), .B2(new_n1029), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT51), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT125), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1384), .B1(new_n495), .B2(new_n505), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1008), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G288), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n812), .A2(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(G8), .A4(new_n1047), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(new_n603), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(new_n605), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n608), .B2(new_n1056), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n1059), .B2(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1048), .B1(new_n1059), .B2(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1055), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT55), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1006), .B(G1384), .C1(new_n495), .C2(new_n505), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1031), .B2(new_n1006), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1971), .B1(new_n1072), .B2(new_n1008), .ZN(new_n1073));
  INV_X1    g648(.A(G2090), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1026), .B1(new_n1075), .B2(new_n1046), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n882), .A2(KEYINPUT70), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n495), .A2(new_n505), .A3(new_n506), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1384), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1074), .B(new_n1076), .C1(new_n1079), .C2(new_n1075), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(G8), .B(new_n1070), .C1(new_n1073), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1067), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1072), .A2(new_n1008), .ZN(new_n1084));
  INV_X1    g659(.A(G1971), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1075), .B(new_n1004), .C1(new_n507), .C2(new_n508), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1026), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1074), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1070), .B1(new_n1092), .B2(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1045), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1084), .A2(new_n1085), .B1(new_n1090), .B2(new_n1074), .ZN(new_n1095));
  INV_X1    g670(.A(G8), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1069), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT125), .A3(new_n1082), .A4(new_n1067), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1071), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n750), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n470), .A2(new_n471), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n464), .B1(new_n1101), .B2(KEYINPUT123), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n480), .B(new_n1100), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  XOR2_X1   g684(.A(G171), .B(KEYINPUT54), .Z(new_n1110));
  NOR3_X1   g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1084), .B2(G2078), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1076), .B1(new_n1079), .B2(new_n1075), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT122), .B(G1961), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1028), .A2(KEYINPUT53), .A3(new_n750), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1113), .A2(new_n1118), .A3(new_n1116), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1111), .A2(new_n1117), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1044), .A2(new_n1094), .A3(new_n1098), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1008), .A2(new_n776), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1124), .B(new_n1071), .C1(new_n1031), .C2(new_n1006), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  AND3_X1   g701(.A1(new_n1047), .A2(KEYINPUT119), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT119), .B1(new_n1047), .B2(new_n1126), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1123), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1031), .A2(new_n1006), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1131), .A2(new_n776), .A3(new_n1008), .A4(new_n1099), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1047), .A2(new_n1126), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1047), .A2(KEYINPUT119), .A3(new_n1126), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1132), .A2(new_n1137), .A3(KEYINPUT120), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1130), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1122), .B1(new_n1139), .B2(new_n564), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n563), .C1(new_n1130), .C2(new_n1138), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1131), .A2(new_n1008), .A3(new_n1099), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1956), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1089), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n918), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n590), .B1(new_n918), .B2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n639), .A2(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1146), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1140), .A2(new_n1141), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1125), .A2(new_n1129), .A3(new_n1123), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT120), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n564), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1139), .A2(new_n1122), .A3(new_n564), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT61), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(KEYINPUT121), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1047), .A2(G2067), .ZN(new_n1174));
  INV_X1    g749(.A(G1348), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1114), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(new_n635), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(KEYINPUT60), .B2(new_n1176), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1162), .A2(new_n1173), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1155), .B1(new_n926), .B2(new_n1176), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1157), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1121), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1119), .A2(G171), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1094), .A2(new_n1098), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1041), .A2(new_n1187), .A3(new_n1043), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1190));
  NOR2_X1   g765(.A1(G288), .A2(G1976), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1190), .A2(new_n1191), .B1(new_n1056), .B2(new_n608), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1067), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1192), .A2(new_n1048), .B1(new_n1193), .B2(new_n1082), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1039), .A2(new_n1029), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1195), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1070), .B1(new_n1197), .B2(G8), .ZN(new_n1198));
  OR3_X1    g773(.A1(new_n1196), .A2(new_n1083), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1097), .A2(new_n1082), .A3(new_n1067), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1195), .A2(G8), .A3(G168), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1194), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1189), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1023), .B1(new_n1183), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n842), .A2(new_n846), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1017), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n800), .A2(new_n803), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1009), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT46), .ZN(new_n1214));
  OAI211_X1 g789(.A(new_n773), .B(new_n1015), .C1(new_n1214), .C2(G1996), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1214), .B1(new_n1009), .B2(G1996), .ZN(new_n1217));
  AOI22_X1  g792(.A1(new_n1215), .A2(new_n1010), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT47), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1020), .A2(new_n1009), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT48), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1220), .B1(new_n1019), .B2(new_n1222), .ZN(new_n1223));
  NOR3_X1   g798(.A1(new_n1212), .A2(new_n1213), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1206), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g800(.A1(new_n462), .A2(G227), .A3(G229), .A4(G401), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n912), .B2(new_n913), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n1228), .A2(new_n989), .ZN(G225));
  INV_X1    g803(.A(G225), .ZN(G308));
endmodule


