

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n727), .A2(n726), .ZN(n522) );
  INV_X1 U556 ( .A(KEYINPUT101), .ZN(n714) );
  XNOR2_X1 U557 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n723) );
  XNOR2_X1 U558 ( .A(n724), .B(n723), .ZN(n735) );
  NAND2_X1 U559 ( .A1(n777), .A2(n682), .ZN(n729) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X1 U562 ( .A(KEYINPUT17), .B(n523), .Z(n881) );
  NAND2_X1 U563 ( .A1(n881), .A2(G138), .ZN(n532) );
  INV_X1 U564 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n526), .ZN(n877) );
  NAND2_X1 U566 ( .A1(G126), .A2(n877), .ZN(n525) );
  AND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U568 ( .A1(G114), .A2(n878), .ZN(n524) );
  NAND2_X1 U569 ( .A1(n525), .A2(n524), .ZN(n530) );
  NAND2_X1 U570 ( .A1(n526), .A2(G2104), .ZN(n527) );
  XNOR2_X2 U571 ( .A(n527), .B(KEYINPUT65), .ZN(n882) );
  NAND2_X1 U572 ( .A1(G102), .A2(n882), .ZN(n528) );
  XNOR2_X1 U573 ( .A(n528), .B(KEYINPUT83), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U575 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U576 ( .A(KEYINPUT84), .B(n533), .Z(G164) );
  INV_X1 U577 ( .A(G651), .ZN(n538) );
  NOR2_X1 U578 ( .A1(G543), .A2(n538), .ZN(n534) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n534), .Z(n643) );
  NAND2_X1 U580 ( .A1(n643), .A2(G64), .ZN(n537) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n644) );
  NOR2_X1 U582 ( .A1(G651), .A2(n644), .ZN(n535) );
  XNOR2_X1 U583 ( .A(KEYINPUT64), .B(n535), .ZN(n639) );
  NAND2_X1 U584 ( .A1(G52), .A2(n639), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n631) );
  NAND2_X1 U587 ( .A1(G90), .A2(n631), .ZN(n540) );
  NOR2_X1 U588 ( .A1(n644), .A2(n538), .ZN(n629) );
  NAND2_X1 U589 ( .A1(G77), .A2(n629), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U592 ( .A1(n543), .A2(n542), .ZN(G171) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G57), .ZN(G237) );
  INV_X1 U595 ( .A(G120), .ZN(G236) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  NAND2_X1 U598 ( .A1(n643), .A2(G62), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G50), .A2(n639), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G88), .A2(n631), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G75), .A2(n629), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT77), .B(n548), .Z(n549) );
  NOR2_X1 U605 ( .A1(n550), .A2(n549), .ZN(G166) );
  NAND2_X1 U606 ( .A1(n631), .A2(G89), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G76), .A2(n629), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U610 ( .A(n554), .B(KEYINPUT5), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G51), .A2(n639), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT70), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G63), .A2(n643), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n831) );
  NAND2_X1 U622 ( .A1(n831), .A2(G567), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U624 ( .A1(n631), .A2(G81), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G68), .A2(n629), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G43), .A2(n639), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n643), .A2(G56), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n953) );
  NAND2_X1 U634 ( .A1(G860), .A2(n953), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n573), .B(KEYINPUT66), .ZN(G153) );
  NAND2_X1 U636 ( .A1(G66), .A2(n643), .ZN(n580) );
  NAND2_X1 U637 ( .A1(G79), .A2(n629), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G54), .A2(n639), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G92), .A2(n631), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT67), .B(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT15), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT68), .B(n582), .ZN(n900) );
  NOR2_X1 U646 ( .A1(G868), .A2(n900), .ZN(n584) );
  INV_X1 U647 ( .A(G868), .ZN(n600) );
  NOR2_X1 U648 ( .A1(G171), .A2(n600), .ZN(n583) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(KEYINPUT69), .B(n585), .ZN(G284) );
  NAND2_X1 U651 ( .A1(n643), .A2(G65), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G53), .A2(n639), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G91), .A2(n631), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G78), .A2(n629), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n957) );
  INV_X1 U658 ( .A(n957), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G286), .A2(n600), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT71), .B(n592), .Z(n594) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n595), .ZN(G297) );
  INV_X1 U664 ( .A(G860), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n597), .A2(n900), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U668 ( .A1(G868), .A2(n900), .ZN(n599) );
  NOR2_X1 U669 ( .A1(G559), .A2(n599), .ZN(n602) );
  AND2_X1 U670 ( .A1(n600), .A2(n953), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G111), .A2(n878), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G99), .A2(n882), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n610) );
  NAND2_X1 U675 ( .A1(n877), .A2(G123), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G135), .A2(n881), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT73), .B(n608), .Z(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n928) );
  XNOR2_X1 U681 ( .A(n928), .B(G2096), .ZN(n612) );
  INV_X1 U682 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(G156) );
  XOR2_X1 U684 ( .A(n953), .B(KEYINPUT74), .Z(n614) );
  NAND2_X1 U685 ( .A1(G559), .A2(n900), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n614), .B(n613), .ZN(n654) );
  NOR2_X1 U687 ( .A1(G860), .A2(n654), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n643), .A2(G67), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G55), .A2(n639), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G93), .A2(n631), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G80), .A2(n629), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n657) );
  XNOR2_X1 U695 ( .A(n621), .B(n657), .ZN(G145) );
  AND2_X1 U696 ( .A1(G47), .A2(n639), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G85), .A2(n631), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G72), .A2(n629), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n643), .A2(G60), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U703 ( .A1(n643), .A2(G61), .ZN(n628) );
  XNOR2_X1 U704 ( .A(KEYINPUT75), .B(n628), .ZN(n635) );
  NAND2_X1 U705 ( .A1(G73), .A2(n629), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n630), .B(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n631), .A2(G86), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT76), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G48), .A2(n639), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G651), .A2(G74), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G49), .A2(n639), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n644), .A2(G87), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n646), .A2(n645), .ZN(G288) );
  XNOR2_X1 U719 ( .A(n957), .B(G290), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n647), .B(G305), .ZN(n651) );
  XNOR2_X1 U721 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n649) );
  XNOR2_X1 U722 ( .A(G288), .B(KEYINPUT78), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U724 ( .A(n651), .B(n650), .Z(n653) );
  XNOR2_X1 U725 ( .A(G166), .B(n657), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n903) );
  XNOR2_X1 U727 ( .A(n903), .B(n654), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n655), .A2(G868), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(KEYINPUT80), .ZN(n659) );
  OR2_X1 U730 ( .A1(n657), .A2(G868), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U738 ( .A1(G220), .A2(G219), .ZN(n664) );
  XOR2_X1 U739 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U740 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U741 ( .A1(G96), .A2(n666), .ZN(n836) );
  AND2_X1 U742 ( .A1(G2106), .A2(n836), .ZN(n672) );
  NOR2_X1 U743 ( .A1(G236), .A2(G237), .ZN(n667) );
  NAND2_X1 U744 ( .A1(G69), .A2(n667), .ZN(n668) );
  XNOR2_X1 U745 ( .A(KEYINPUT81), .B(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n669), .A2(G108), .ZN(n835) );
  NAND2_X1 U747 ( .A1(G567), .A2(n835), .ZN(n670) );
  XOR2_X1 U748 ( .A(KEYINPUT82), .B(n670), .Z(n671) );
  NOR2_X1 U749 ( .A1(n672), .A2(n671), .ZN(G319) );
  INV_X1 U750 ( .A(G319), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n834) );
  NAND2_X1 U753 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G125), .A2(n877), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G113), .A2(n878), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n681) );
  NAND2_X1 U757 ( .A1(G101), .A2(n882), .ZN(n677) );
  XOR2_X1 U758 ( .A(KEYINPUT23), .B(n677), .Z(n679) );
  NAND2_X1 U759 ( .A1(n881), .A2(G137), .ZN(n678) );
  NAND2_X1 U760 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U761 ( .A1(n681), .A2(n680), .ZN(G160) );
  INV_X1 U762 ( .A(G166), .ZN(G303) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n776) );
  INV_X1 U764 ( .A(n776), .ZN(n682) );
  INV_X1 U765 ( .A(n729), .ZN(n698) );
  BUF_X1 U766 ( .A(n698), .Z(n688) );
  XNOR2_X1 U767 ( .A(G1961), .B(KEYINPUT96), .ZN(n985) );
  NOR2_X1 U768 ( .A1(n688), .A2(n985), .ZN(n683) );
  XNOR2_X1 U769 ( .A(n683), .B(KEYINPUT97), .ZN(n685) );
  XNOR2_X1 U770 ( .A(G2078), .B(KEYINPUT25), .ZN(n1010) );
  NAND2_X1 U771 ( .A1(n688), .A2(n1010), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n720), .A2(G171), .ZN(n713) );
  NAND2_X1 U774 ( .A1(G2072), .A2(n698), .ZN(n686) );
  XNOR2_X1 U775 ( .A(n686), .B(KEYINPUT98), .ZN(n687) );
  XNOR2_X1 U776 ( .A(KEYINPUT27), .B(n687), .ZN(n690) );
  INV_X1 U777 ( .A(G1956), .ZN(n956) );
  NOR2_X1 U778 ( .A1(n688), .A2(n956), .ZN(n689) );
  NOR2_X1 U779 ( .A1(n690), .A2(n689), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n692), .A2(n957), .ZN(n691) );
  XOR2_X1 U781 ( .A(n691), .B(KEYINPUT28), .Z(n710) );
  NAND2_X1 U782 ( .A1(n957), .A2(n692), .ZN(n708) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n698), .ZN(n693) );
  XNOR2_X1 U784 ( .A(KEYINPUT26), .B(n693), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n694), .A2(n953), .ZN(n697) );
  NAND2_X1 U786 ( .A1(G1341), .A2(n729), .ZN(n695) );
  XNOR2_X1 U787 ( .A(KEYINPUT99), .B(n695), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n900), .A2(n704), .ZN(n703) );
  AND2_X1 U790 ( .A1(n698), .A2(G2067), .ZN(n699) );
  XOR2_X1 U791 ( .A(n699), .B(KEYINPUT100), .Z(n701) );
  NAND2_X1 U792 ( .A1(n729), .A2(G1348), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n706) );
  OR2_X1 U795 ( .A1(n900), .A2(n704), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U799 ( .A(KEYINPUT29), .B(n711), .Z(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n733) );
  NAND2_X1 U801 ( .A1(G8), .A2(n729), .ZN(n769) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n769), .ZN(n727) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n729), .ZN(n725) );
  NOR2_X1 U804 ( .A1(n727), .A2(n725), .ZN(n715) );
  XNOR2_X1 U805 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n716), .A2(G8), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n717), .B(KEYINPUT30), .ZN(n718) );
  NOR2_X1 U808 ( .A1(G168), .A2(n718), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n719), .B(KEYINPUT102), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n720), .A2(G171), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n733), .A2(n735), .ZN(n728) );
  AND2_X1 U813 ( .A1(G8), .A2(n725), .ZN(n726) );
  AND2_X1 U814 ( .A1(n728), .A2(n522), .ZN(n744) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n769), .ZN(n731) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n732), .A2(G303), .ZN(n736) );
  AND2_X1 U819 ( .A1(n733), .A2(n736), .ZN(n734) );
  NAND2_X1 U820 ( .A1(n735), .A2(n734), .ZN(n740) );
  INV_X1 U821 ( .A(n736), .ZN(n737) );
  OR2_X1 U822 ( .A1(n737), .A2(G286), .ZN(n738) );
  AND2_X1 U823 ( .A1(G8), .A2(n738), .ZN(n739) );
  NAND2_X1 U824 ( .A1(n740), .A2(n739), .ZN(n742) );
  XOR2_X1 U825 ( .A(KEYINPUT104), .B(KEYINPUT32), .Z(n741) );
  XNOR2_X1 U826 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U827 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U828 ( .A(n745), .B(KEYINPUT105), .ZN(n762) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n746) );
  XNOR2_X1 U831 ( .A(KEYINPUT106), .B(n746), .ZN(n747) );
  NOR2_X1 U832 ( .A1(n959), .A2(n747), .ZN(n750) );
  NOR2_X1 U833 ( .A1(G1981), .A2(G305), .ZN(n748) );
  XNOR2_X1 U834 ( .A(KEYINPUT24), .B(n748), .ZN(n758) );
  INV_X1 U835 ( .A(n758), .ZN(n749) );
  AND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n762), .A2(n751), .ZN(n760) );
  NAND2_X1 U838 ( .A1(G288), .A2(G1976), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT107), .ZN(n961) );
  INV_X1 U840 ( .A(n961), .ZN(n756) );
  XNOR2_X1 U841 ( .A(KEYINPUT108), .B(G1981), .ZN(n753) );
  XNOR2_X1 U842 ( .A(n753), .B(G305), .ZN(n951) );
  NAND2_X1 U843 ( .A1(n959), .A2(KEYINPUT33), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n769), .A2(n754), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n951), .A2(n755), .ZN(n764) );
  AND2_X1 U846 ( .A1(n756), .A2(n764), .ZN(n757) );
  OR2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  OR2_X1 U849 ( .A1(n761), .A2(n769), .ZN(n775) );
  INV_X1 U850 ( .A(n762), .ZN(n768) );
  NAND2_X1 U851 ( .A1(G8), .A2(G166), .ZN(n763) );
  NOR2_X1 U852 ( .A1(G2090), .A2(n763), .ZN(n766) );
  NAND2_X1 U853 ( .A1(KEYINPUT33), .A2(n764), .ZN(n771) );
  INV_X1 U854 ( .A(n771), .ZN(n765) );
  OR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n773) );
  INV_X1 U857 ( .A(n769), .ZN(n770) );
  AND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  OR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n816) );
  NOR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n826) );
  NAND2_X1 U862 ( .A1(G140), .A2(n881), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G104), .A2(n882), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n780), .ZN(n786) );
  NAND2_X1 U866 ( .A1(n877), .A2(G128), .ZN(n781) );
  XOR2_X1 U867 ( .A(KEYINPUT85), .B(n781), .Z(n783) );
  NAND2_X1 U868 ( .A1(n878), .A2(G116), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U870 ( .A(n784), .B(KEYINPUT35), .Z(n785) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U872 ( .A(KEYINPUT36), .B(n787), .Z(n788) );
  XOR2_X1 U873 ( .A(KEYINPUT86), .B(n788), .Z(n898) );
  XNOR2_X1 U874 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NOR2_X1 U875 ( .A1(n898), .A2(n824), .ZN(n940) );
  NAND2_X1 U876 ( .A1(n826), .A2(n940), .ZN(n822) );
  NAND2_X1 U877 ( .A1(G119), .A2(n877), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G107), .A2(n878), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U880 ( .A(KEYINPUT87), .B(n791), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G131), .A2(n881), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT89), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G95), .A2(n882), .ZN(n793) );
  XOR2_X1 U884 ( .A(KEYINPUT88), .B(n793), .Z(n794) );
  NOR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U887 ( .A(KEYINPUT90), .B(n798), .ZN(n888) );
  AND2_X1 U888 ( .A1(n888), .A2(G1991), .ZN(n810) );
  NAND2_X1 U889 ( .A1(G141), .A2(n881), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(KEYINPUT92), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G105), .A2(n882), .ZN(n800) );
  XNOR2_X1 U892 ( .A(n800), .B(KEYINPUT38), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n877), .A2(G129), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G117), .A2(n878), .ZN(n803) );
  XNOR2_X1 U896 ( .A(KEYINPUT91), .B(n803), .ZN(n804) );
  NOR2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U899 ( .A(KEYINPUT93), .B(n808), .ZN(n868) );
  INV_X1 U900 ( .A(G1996), .ZN(n1008) );
  NOR2_X1 U901 ( .A1(n868), .A2(n1008), .ZN(n809) );
  NOR2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n938) );
  XOR2_X1 U903 ( .A(n826), .B(KEYINPUT94), .Z(n811) );
  NOR2_X1 U904 ( .A1(n938), .A2(n811), .ZN(n819) );
  XNOR2_X1 U905 ( .A(KEYINPUT95), .B(n819), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n822), .A2(n812), .ZN(n814) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n965) );
  AND2_X1 U908 ( .A1(n965), .A2(n826), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n829) );
  AND2_X1 U911 ( .A1(n1008), .A2(n868), .ZN(n933) );
  NOR2_X1 U912 ( .A1(n888), .A2(G1991), .ZN(n929) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n929), .A2(n817), .ZN(n818) );
  NOR2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n933), .A2(n820), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n898), .A2(n824), .ZN(n942) );
  NAND2_X1 U920 ( .A1(n825), .A2(n942), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U926 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(G2096), .B(G2072), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2090), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U937 ( .A(KEYINPUT112), .B(G2678), .Z(n840) );
  XNOR2_X1 U938 ( .A(G2100), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT111), .B(KEYINPUT113), .Z(n842) );
  XNOR2_X1 U941 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U947 ( .A(KEYINPUT116), .B(G1976), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1956), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n851), .B(KEYINPUT41), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U953 ( .A(G1981), .B(G1966), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1971), .B(G1961), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2474), .B(KEYINPUT115), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n877), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT44), .B(n860), .Z(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT117), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G112), .A2(n878), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G136), .A2(n881), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G100), .A2(n882), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U968 ( .A(G160), .B(n868), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G139), .A2(n881), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G103), .A2(n882), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G127), .A2(n877), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G115), .A2(n878), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n924) );
  XNOR2_X1 U977 ( .A(n876), .B(n924), .ZN(n894) );
  NAND2_X1 U978 ( .A1(G130), .A2(n877), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G142), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G106), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n889) );
  XOR2_X1 U986 ( .A(n889), .B(n888), .Z(n890) );
  XOR2_X1 U987 ( .A(n890), .B(KEYINPUT48), .Z(n892) );
  XNOR2_X1 U988 ( .A(G162), .B(KEYINPUT46), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n896) );
  XNOR2_X1 U991 ( .A(G164), .B(n928), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U993 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U994 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U995 ( .A(KEYINPUT118), .B(n953), .Z(n902) );
  INV_X1 U996 ( .A(n900), .ZN(n969) );
  XNOR2_X1 U997 ( .A(G171), .B(n969), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n903), .B(G286), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(G397) );
  XNOR2_X1 U1002 ( .A(G2451), .B(G2435), .ZN(n916) );
  XOR2_X1 U1003 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G2454), .B(G2430), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2438), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2427), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G171), .ZN(G301) );
  INV_X1 U1022 ( .A(G69), .ZN(G235) );
  INV_X1 U1023 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1024 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(KEYINPUT50), .B(n927), .ZN(n946) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT51), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT119), .B(n941), .Z(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(n944), .Z(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G29), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(G11), .A2(n949), .ZN(n1028) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n975) );
  XOR2_X1 U1045 ( .A(G1966), .B(G168), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(KEYINPUT57), .B(n952), .Z(n973) );
  XOR2_X1 U1048 ( .A(n953), .B(G1341), .Z(n955) );
  XOR2_X1 U1049 ( .A(G171), .B(G1961), .Z(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n968) );
  XNOR2_X1 U1051 ( .A(n957), .B(n956), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n963) );
  XOR2_X1 U1053 ( .A(G1971), .B(G166), .Z(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n966), .B(KEYINPUT124), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(G1348), .B(n969), .ZN(n970) );
  NOR2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1061 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1062 ( .A1(n975), .A2(n974), .ZN(n1001) );
  INV_X1 U1063 ( .A(G16), .ZN(n999) );
  XNOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(n976), .B(G4), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(G1956), .B(G20), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G19), .B(G1341), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1070 ( .A(KEYINPUT125), .B(G1981), .Z(n981) );
  XNOR2_X1 U1071 ( .A(G6), .B(n981), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(KEYINPUT60), .B(n984), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(n985), .B(G5), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G21), .B(G1966), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n996) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G23), .B(G1976), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(n994), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(KEYINPUT61), .B(n997), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(KEYINPUT126), .B(n1002), .Z(n1026) );
  XOR2_X1 U1089 ( .A(G2090), .B(G35), .Z(n1005) );
  XOR2_X1 U1090 ( .A(G34), .B(KEYINPUT54), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(n1003), .B(G2084), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1021) );
  XNOR2_X1 U1093 ( .A(G1991), .B(G25), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G33), .B(G2072), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(G32), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(G28), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G27), .B(n1010), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT121), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G26), .B(G2067), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT122), .B(n1018), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT53), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT123), .B(n1022), .Z(n1023) );
  NOR2_X1 U1108 ( .A1(G29), .A2(n1023), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(KEYINPUT55), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

