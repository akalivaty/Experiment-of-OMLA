

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585;

  XNOR2_X1 U320 ( .A(n430), .B(n429), .ZN(n448) );
  XNOR2_X1 U321 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n429) );
  XOR2_X1 U322 ( .A(G92GAT), .B(G85GAT), .Z(n374) );
  XNOR2_X1 U323 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U324 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U325 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U326 ( .A(n347), .B(n346), .ZN(n577) );
  XNOR2_X1 U327 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U328 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n294) );
  XOR2_X1 U330 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n289) );
  NAND2_X1 U331 ( .A1(G227GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U332 ( .A(n289), .B(n288), .ZN(n292) );
  XOR2_X1 U333 ( .A(G127GAT), .B(KEYINPUT82), .Z(n291) );
  XNOR2_X1 U334 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n439) );
  XNOR2_X1 U336 ( .A(n292), .B(n439), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n296) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n295), .B(G120GAT), .ZN(n342) );
  XOR2_X1 U340 ( .A(n296), .B(n342), .Z(n304) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(G15GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n297), .B(G113GAT), .ZN(n358) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n299) );
  XNOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n300), .B(G183GAT), .Z(n302) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n428) );
  XNOR2_X1 U349 ( .A(n358), .B(n428), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n533) );
  XOR2_X1 U351 ( .A(KEYINPUT90), .B(G218GAT), .Z(n306) );
  XNOR2_X1 U352 ( .A(G211GAT), .B(G204GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U354 ( .A(KEYINPUT21), .B(n307), .Z(n417) );
  XOR2_X1 U355 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT88), .B(KEYINPUT93), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n314) );
  XNOR2_X1 U358 ( .A(KEYINPUT2), .B(KEYINPUT91), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n310), .B(KEYINPUT92), .ZN(n311) );
  XOR2_X1 U360 ( .A(n311), .B(KEYINPUT3), .Z(n313) );
  XNOR2_X1 U361 ( .A(G155GAT), .B(G162GAT), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n443) );
  XOR2_X1 U363 ( .A(n314), .B(n443), .Z(n326) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n315), .B(G148GAT), .ZN(n343) );
  XOR2_X1 U366 ( .A(KEYINPUT24), .B(n343), .Z(n317) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n319) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(KEYINPUT22), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U372 ( .A(n320), .B(KEYINPUT87), .Z(n322) );
  XOR2_X1 U373 ( .A(G141GAT), .B(G22GAT), .Z(n352) );
  XNOR2_X1 U374 ( .A(G50GAT), .B(n352), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n417), .B(n327), .ZN(n468) );
  INV_X1 U379 ( .A(G64GAT), .ZN(n328) );
  NAND2_X1 U380 ( .A1(KEYINPUT75), .A2(n328), .ZN(n331) );
  INV_X1 U381 ( .A(KEYINPUT75), .ZN(n329) );
  NAND2_X1 U382 ( .A1(n329), .A2(G64GAT), .ZN(n330) );
  NAND2_X1 U383 ( .A1(n331), .A2(n330), .ZN(n421) );
  XNOR2_X1 U384 ( .A(n374), .B(n421), .ZN(n333) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT31), .B(KEYINPUT77), .Z(n335) );
  XNOR2_X1 U388 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n337) );
  AND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(KEYINPUT76), .B(n340), .ZN(n347) );
  XNOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n341), .B(KEYINPUT73), .ZN(n394) );
  XOR2_X1 U394 ( .A(n342), .B(n394), .Z(n345) );
  XOR2_X1 U395 ( .A(n343), .B(KEYINPUT33), .Z(n344) );
  XNOR2_X1 U396 ( .A(n577), .B(KEYINPUT41), .ZN(n507) );
  INV_X1 U397 ( .A(n507), .ZN(n452) );
  XOR2_X1 U398 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n349) );
  XNOR2_X1 U399 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n365) );
  XOR2_X1 U401 ( .A(KEYINPUT70), .B(G1GAT), .Z(n390) );
  XOR2_X1 U402 ( .A(KEYINPUT71), .B(n390), .Z(n351) );
  XOR2_X1 U403 ( .A(G197GAT), .B(G8GAT), .Z(n418) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(n418), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U406 ( .A(n353), .B(n352), .Z(n363) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(KEYINPUT69), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n354), .B(G29GAT), .ZN(n355) );
  XOR2_X1 U409 ( .A(n355), .B(KEYINPUT8), .Z(n357) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n384) );
  XOR2_X1 U412 ( .A(n358), .B(KEYINPUT68), .Z(n360) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n384), .B(n361), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n365), .B(n364), .ZN(n571) );
  NAND2_X1 U418 ( .A1(n452), .A2(n571), .ZN(n368) );
  INV_X1 U419 ( .A(n368), .ZN(n367) );
  INV_X1 U420 ( .A(KEYINPUT46), .ZN(n366) );
  NAND2_X1 U421 ( .A1(n367), .A2(n366), .ZN(n370) );
  NAND2_X1 U422 ( .A1(KEYINPUT46), .A2(n368), .ZN(n369) );
  NAND2_X1 U423 ( .A1(n370), .A2(n369), .ZN(n407) );
  XOR2_X1 U424 ( .A(G162GAT), .B(G218GAT), .Z(n372) );
  XNOR2_X1 U425 ( .A(G43GAT), .B(G99GAT), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U427 ( .A(n374), .B(n373), .Z(n376) );
  NAND2_X1 U428 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U430 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n378) );
  XNOR2_X1 U431 ( .A(G190GAT), .B(G106GAT), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U433 ( .A(n380), .B(n379), .Z(n386) );
  XOR2_X1 U434 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n382) );
  XNOR2_X1 U435 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n541) );
  XOR2_X1 U439 ( .A(G155GAT), .B(G78GAT), .Z(n388) );
  XNOR2_X1 U440 ( .A(G22GAT), .B(G211GAT), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U442 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U445 ( .A(n393), .B(KEYINPUT12), .Z(n396) );
  XNOR2_X1 U446 ( .A(n394), .B(KEYINPUT14), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n396), .B(n395), .ZN(n404) );
  XOR2_X1 U448 ( .A(G127GAT), .B(G71GAT), .Z(n398) );
  XNOR2_X1 U449 ( .A(G15GAT), .B(G183GAT), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U451 ( .A(KEYINPUT15), .B(G64GAT), .Z(n400) );
  XNOR2_X1 U452 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U454 ( .A(n402), .B(n401), .Z(n403) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n580) );
  INV_X1 U456 ( .A(n580), .ZN(n405) );
  AND2_X1 U457 ( .A1(n541), .A2(n405), .ZN(n406) );
  AND2_X1 U458 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U459 ( .A(n408), .B(KEYINPUT47), .ZN(n415) );
  XOR2_X1 U460 ( .A(KEYINPUT114), .B(KEYINPUT45), .Z(n409) );
  XNOR2_X1 U461 ( .A(KEYINPUT64), .B(n409), .ZN(n411) );
  XOR2_X1 U462 ( .A(KEYINPUT36), .B(n541), .Z(n582) );
  NAND2_X1 U463 ( .A1(n580), .A2(n582), .ZN(n410) );
  XOR2_X1 U464 ( .A(n411), .B(n410), .Z(n412) );
  NOR2_X1 U465 ( .A1(n577), .A2(n412), .ZN(n413) );
  XNOR2_X1 U466 ( .A(KEYINPUT72), .B(n571), .ZN(n560) );
  INV_X1 U467 ( .A(n560), .ZN(n475) );
  NAND2_X1 U468 ( .A1(n413), .A2(n475), .ZN(n414) );
  NAND2_X1 U469 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(KEYINPUT48), .B(n416), .ZN(n548) );
  XOR2_X1 U471 ( .A(G92GAT), .B(n417), .Z(n420) );
  XNOR2_X1 U472 ( .A(G36GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n426) );
  XOR2_X1 U474 ( .A(KEYINPUT97), .B(n421), .Z(n423) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT81), .B(n424), .Z(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n480) );
  NAND2_X1 U480 ( .A1(n548), .A2(n480), .ZN(n430) );
  XOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n432) );
  XNOR2_X1 U482 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n447) );
  XOR2_X1 U484 ( .A(G85GAT), .B(G148GAT), .Z(n434) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(G141GAT), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U487 ( .A(G57GAT), .B(G120GAT), .Z(n436) );
  XNOR2_X1 U488 ( .A(G113GAT), .B(G1GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U490 ( .A(n438), .B(n437), .Z(n445) );
  XOR2_X1 U491 ( .A(n439), .B(KEYINPUT96), .Z(n441) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U496 ( .A(n447), .B(n446), .Z(n520) );
  NAND2_X1 U497 ( .A1(n448), .A2(n520), .ZN(n569) );
  NOR2_X1 U498 ( .A1(n468), .A2(n569), .ZN(n449) );
  XNOR2_X1 U499 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NOR2_X1 U500 ( .A1(n533), .A2(n450), .ZN(n451) );
  XNOR2_X1 U501 ( .A(KEYINPUT122), .B(n451), .ZN(n566) );
  NAND2_X1 U502 ( .A1(n566), .A2(n452), .ZN(n456) );
  XOR2_X1 U503 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n454) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT56), .Z(n453) );
  INV_X1 U505 ( .A(n533), .ZN(n457) );
  NAND2_X1 U506 ( .A1(n480), .A2(n457), .ZN(n458) );
  XNOR2_X1 U507 ( .A(KEYINPUT99), .B(n458), .ZN(n459) );
  NOR2_X1 U508 ( .A1(n468), .A2(n459), .ZN(n460) );
  XNOR2_X1 U509 ( .A(n460), .B(KEYINPUT25), .ZN(n463) );
  XOR2_X1 U510 ( .A(n480), .B(KEYINPUT27), .Z(n465) );
  NAND2_X1 U511 ( .A1(n468), .A2(n533), .ZN(n461) );
  XOR2_X1 U512 ( .A(KEYINPUT26), .B(n461), .Z(n547) );
  INV_X1 U513 ( .A(n547), .ZN(n570) );
  OR2_X1 U514 ( .A1(n465), .A2(n570), .ZN(n462) );
  NAND2_X1 U515 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U516 ( .A1(n464), .A2(n520), .ZN(n471) );
  XNOR2_X1 U517 ( .A(n533), .B(KEYINPUT86), .ZN(n469) );
  NOR2_X1 U518 ( .A1(n520), .A2(n465), .ZN(n466) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(n466), .Z(n550) );
  XOR2_X1 U520 ( .A(KEYINPUT28), .B(KEYINPUT65), .Z(n467) );
  XNOR2_X1 U521 ( .A(n468), .B(n467), .ZN(n485) );
  NOR2_X1 U522 ( .A1(n550), .A2(n485), .ZN(n531) );
  NAND2_X1 U523 ( .A1(n469), .A2(n531), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U525 ( .A(n472), .B(KEYINPUT100), .ZN(n489) );
  NAND2_X1 U526 ( .A1(n541), .A2(n580), .ZN(n473) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U528 ( .A1(n489), .A2(n474), .ZN(n508) );
  NOR2_X1 U529 ( .A1(n577), .A2(n475), .ZN(n476) );
  XNOR2_X1 U530 ( .A(n476), .B(KEYINPUT78), .ZN(n492) );
  NAND2_X1 U531 ( .A1(n508), .A2(n492), .ZN(n477) );
  XOR2_X1 U532 ( .A(KEYINPUT101), .B(n477), .Z(n486) );
  NOR2_X1 U533 ( .A1(n520), .A2(n486), .ZN(n478) );
  XOR2_X1 U534 ( .A(G1GAT), .B(n478), .Z(n479) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n479), .ZN(G1324GAT) );
  INV_X1 U536 ( .A(n480), .ZN(n523) );
  NOR2_X1 U537 ( .A1(n523), .A2(n486), .ZN(n481) );
  XOR2_X1 U538 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n533), .A2(n486), .ZN(n484) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n485), .ZN(n528) );
  NOR2_X1 U544 ( .A1(n528), .A2(n486), .ZN(n488) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  NAND2_X1 U547 ( .A1(n582), .A2(n489), .ZN(n490) );
  NOR2_X1 U548 ( .A1(n580), .A2(n490), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n491), .Z(n519) );
  NAND2_X1 U550 ( .A1(n492), .A2(n519), .ZN(n495) );
  XOR2_X1 U551 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT104), .B(n493), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n505) );
  NOR2_X1 U554 ( .A1(n505), .A2(n520), .ZN(n499) );
  XOR2_X1 U555 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT106), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n523), .A2(n505), .ZN(n500) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n502) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(KEYINPUT108), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n504) );
  NOR2_X1 U564 ( .A1(n533), .A2(n505), .ZN(n503) );
  XOR2_X1 U565 ( .A(n504), .B(n503), .Z(G1330GAT) );
  NOR2_X1 U566 ( .A1(n528), .A2(n505), .ZN(n506) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  NOR2_X1 U568 ( .A1(n507), .A2(n571), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n518), .A2(n508), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n509), .B(KEYINPUT110), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n520), .A2(n515), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(KEYINPUT111), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n515), .A2(n523), .ZN(n513) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n533), .A2(n515), .ZN(n514) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n528), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n520), .A2(n527), .ZN(n521) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n521), .Z(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT112), .B(n522), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n533), .A2(n527), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1338GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT115), .Z(n535) );
  NAND2_X1 U595 ( .A1(n548), .A2(n531), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n542), .A2(n560), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U600 ( .A1(n542), .A2(n452), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U603 ( .A1(n542), .A2(n580), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n544) );
  INV_X1 U607 ( .A(n541), .ZN(n565) );
  NAND2_X1 U608 ( .A1(n542), .A2(n565), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT117), .Z(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  XOR2_X1 U612 ( .A(G141GAT), .B(KEYINPUT119), .Z(n552) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n558), .A2(n571), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U619 ( .A1(n558), .A2(n452), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n580), .A2(n558), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n566), .A2(n580), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT124), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT125), .B(n564), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n583), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(n574), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U643 ( .A1(n583), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n583), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

