//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(KEYINPUT1), .C1(new_n192), .C2(G146), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n188), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n194), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT73), .B(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(new_n188), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n200), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n191), .B(new_n193), .C1(new_n206), .C2(new_n188), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G224), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G953), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G110), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT8), .ZN(new_n220));
  INV_X1    g034(.A(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT2), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G116), .B(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n221), .B1(new_n226), .B2(KEYINPUT5), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n229), .A2(KEYINPUT5), .A3(G119), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n230), .A2(KEYINPUT84), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(KEYINPUT84), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n235), .A2(KEYINPUT77), .A3(G107), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT76), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G107), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G104), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n235), .A2(G107), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(G104), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT76), .B(KEYINPUT3), .C1(new_n244), .C2(KEYINPUT77), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n238), .A2(new_n242), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G104), .B(G107), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT78), .B1(new_n247), .B2(new_n243), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT78), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(G101), .C1(new_n240), .C2(new_n241), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AND4_X1   g065(.A1(new_n227), .A2(new_n233), .A3(new_n246), .A4(new_n251), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n227), .A2(new_n233), .B1(new_n246), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n220), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n210), .B1(new_n202), .B2(new_n203), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n215), .A2(KEYINPUT7), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n216), .A2(new_n254), .A3(new_n255), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n246), .A2(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT80), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(new_n251), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n261), .A2(new_n227), .A3(new_n233), .A4(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n229), .A2(G119), .ZN(new_n265));
  INV_X1    g079(.A(G119), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G116), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n222), .B(new_n224), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n227), .A3(KEYINPUT66), .ZN(new_n269));
  OR3_X1    g083(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n242), .A2(new_n245), .ZN(new_n274));
  INV_X1    g088(.A(new_n238), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n273), .B(G101), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n235), .A2(G107), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n244), .B2(KEYINPUT76), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n237), .B1(new_n241), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n278), .B1(new_n280), .B2(KEYINPUT3), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n243), .B1(new_n281), .B2(new_n238), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n246), .A2(KEYINPUT4), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n272), .B(new_n276), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n264), .A2(new_n284), .A3(new_n219), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n259), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n214), .B1(new_n204), .B2(new_n211), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n287), .A2(KEYINPUT7), .B1(new_n256), .B2(new_n257), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n255), .B1(new_n288), .B2(new_n254), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT88), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n285), .A2(KEYINPUT6), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n219), .B1(new_n264), .B2(new_n284), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT86), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n264), .A2(new_n284), .ZN(new_n296));
  INV_X1    g110(.A(new_n219), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(KEYINPUT6), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n256), .B(new_n214), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT86), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n298), .A2(new_n301), .A3(KEYINPUT6), .A4(new_n285), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n299), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT88), .B(new_n187), .C1(new_n286), .C2(new_n289), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n292), .A2(new_n303), .A3(new_n306), .A4(new_n304), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT81), .B(G469), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n261), .A2(KEYINPUT10), .A3(new_n202), .A4(new_n263), .ZN(new_n315));
  INV_X1    g129(.A(G137), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G134), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT11), .B1(new_n318), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT11), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n316), .A3(G134), .ZN(new_n321));
  AOI211_X1 g135(.A(G131), .B(new_n317), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n321), .ZN(new_n324));
  INV_X1    g138(.A(new_n317), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n194), .A2(KEYINPUT79), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n194), .A2(KEYINPUT79), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n195), .A2(G128), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n329), .A2(new_n330), .B1(new_n200), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n332), .B2(new_n260), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n208), .A2(new_n209), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n334), .B(new_n276), .C1(new_n282), .C2(new_n283), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n315), .A2(new_n327), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G140), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n338), .A2(G227), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n337), .B(new_n339), .Z(new_n340));
  NAND2_X1  g154(.A1(new_n331), .A2(new_n200), .ZN(new_n341));
  INV_X1    g155(.A(new_n330), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n194), .A2(KEYINPUT79), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n251), .A3(new_n246), .ZN(new_n345));
  INV_X1    g159(.A(new_n194), .ZN(new_n346));
  INV_X1    g160(.A(new_n198), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n197), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n348));
  OAI21_X1  g162(.A(G128), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(new_n200), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n260), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n327), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT12), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT12), .ZN(new_n355));
  AOI211_X1 g169(.A(new_n355), .B(new_n327), .C1(new_n345), .C2(new_n351), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n336), .B(new_n340), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n335), .A2(new_n333), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n202), .A2(KEYINPUT10), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n246), .A2(new_n251), .A3(new_n262), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n262), .B1(new_n246), .B2(new_n251), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n340), .B1(new_n363), .B2(new_n336), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n357), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT82), .B(new_n340), .C1(new_n363), .C2(new_n336), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n187), .B(new_n314), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n336), .A2(new_n340), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n336), .B1(new_n354), .B2(new_n356), .ZN(new_n370));
  INV_X1    g184(.A(new_n340), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n369), .A2(new_n363), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G469), .B1(new_n372), .B2(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n313), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n376), .ZN(new_n378));
  AOI211_X1 g192(.A(KEYINPUT83), .B(new_n378), .C1(new_n368), .C2(new_n373), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n312), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(G234), .B2(new_n187), .ZN(new_n382));
  INV_X1    g196(.A(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G125), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n203), .A2(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n190), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(G146), .A3(new_n388), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(G119), .B(G128), .Z(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT24), .B(G110), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n266), .B2(G128), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n397), .B(new_n398), .C1(G119), .C2(new_n188), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(G110), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G125), .B(G140), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(new_n190), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n399), .A2(G110), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n394), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n391), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT74), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT22), .B(G137), .Z(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n400), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(new_n390), .B2(new_n391), .ZN(new_n415));
  INV_X1    g229(.A(new_n407), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n417), .A3(new_n187), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT25), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n382), .B1(new_n420), .B2(KEYINPUT75), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n418), .A2(new_n419), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT75), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n413), .A2(new_n417), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n382), .A2(G902), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n422), .A2(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n334), .B1(new_n322), .B2(new_n326), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n324), .A2(new_n323), .A3(new_n325), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n316), .B2(G134), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n318), .A2(KEYINPUT64), .A3(G137), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n433), .A2(new_n434), .B1(G134), .B2(new_n316), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n323), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n430), .B1(new_n350), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n272), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n430), .B(new_n271), .C1(new_n350), .C2(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT28), .ZN(new_n441));
  INV_X1    g255(.A(new_n439), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n442), .A2(KEYINPUT28), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT26), .B(G101), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n338), .A3(G210), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n445), .B(KEYINPUT68), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n455), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n444), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n437), .A2(KEYINPUT30), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n430), .B(new_n462), .C1(new_n350), .C2(new_n436), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n442), .B1(new_n464), .B2(new_n272), .ZN(new_n465));
  INV_X1    g279(.A(new_n459), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT31), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n271), .B1(new_n461), .B2(new_n463), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT31), .ZN(new_n469));
  NOR4_X1   g283(.A1(new_n468), .A2(new_n469), .A3(new_n459), .A4(new_n442), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n460), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G472), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n187), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT32), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(KEYINPUT32), .A3(new_n472), .A4(new_n187), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n439), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n433), .A2(new_n434), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n316), .A2(G134), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n323), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n322), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n202), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(KEYINPUT69), .A3(new_n271), .A4(new_n430), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n438), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT28), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n459), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n443), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n459), .B1(new_n468), .B2(new_n442), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n487), .B(new_n491), .C1(new_n444), .C2(new_n459), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n486), .A2(new_n493), .A3(new_n443), .A4(new_n488), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n490), .A2(new_n492), .A3(new_n187), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G472), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n475), .A2(new_n476), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT71), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT71), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n475), .A2(new_n496), .A3(new_n499), .A4(new_n476), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n429), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n338), .A2(G952), .ZN(new_n502));
  NAND2_X1  g316(.A1(G234), .A2(G237), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(G902), .A3(G953), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n448), .A2(new_n338), .A3(G214), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(G143), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n323), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT17), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n511), .B(new_n192), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G131), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n323), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n390), .A2(new_n391), .A3(new_n514), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G113), .B(G122), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n235), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(KEYINPUT18), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n512), .B1(new_n524), .B2(new_n323), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n385), .A2(new_n386), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n190), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n523), .B(new_n525), .C1(new_n527), .C2(new_n403), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n520), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n516), .A2(new_n517), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n402), .A2(KEYINPUT19), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n526), .B2(KEYINPUT19), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n391), .B(new_n530), .C1(new_n532), .C2(G146), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n522), .B1(new_n533), .B2(new_n528), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n510), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT20), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(new_n510), .C1(new_n529), .C2(new_n534), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n522), .B1(new_n520), .B2(new_n528), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n187), .B1(new_n529), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n536), .A2(new_n538), .B1(G475), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n375), .A2(new_n381), .A3(G953), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT92), .ZN(new_n547));
  INV_X1    g361(.A(G122), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G116), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n229), .A2(G122), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G107), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n550), .A3(new_n239), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n192), .A2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n188), .A2(G143), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n318), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n192), .A2(G128), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT89), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT13), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n555), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n568));
  OAI211_X1 g382(.A(KEYINPUT90), .B(new_n555), .C1(new_n568), .C2(new_n560), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n564), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n558), .B1(new_n572), .B2(G134), .ZN(new_n573));
  OAI21_X1  g387(.A(G134), .B1(new_n566), .B2(new_n560), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n557), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n553), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT91), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT14), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n229), .B2(G122), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n581), .B2(new_n550), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n578), .B1(new_n582), .B2(new_n577), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n576), .B1(G107), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n547), .B1(new_n573), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n569), .A2(new_n571), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n570), .A2(new_n556), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT90), .B1(new_n587), .B2(new_n555), .ZN(new_n588));
  OAI21_X1  g402(.A(G134), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n558), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n546), .B(KEYINPUT92), .Z(new_n592));
  AND2_X1   g406(.A1(new_n575), .A2(new_n553), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n583), .A2(G107), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n596), .A3(new_n187), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n585), .A2(new_n596), .A3(KEYINPUT93), .A4(new_n187), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n545), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n597), .A2(new_n545), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT94), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n601), .A2(KEYINPUT94), .A3(new_n602), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n509), .B(new_n542), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n380), .A2(new_n501), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT95), .B(G101), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  AOI21_X1  g422(.A(KEYINPUT33), .B1(new_n585), .B2(new_n596), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n589), .A2(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n547), .B1(new_n610), .B2(KEYINPUT96), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(new_n592), .C1(new_n573), .C2(new_n584), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n609), .B1(new_n614), .B2(KEYINPUT33), .ZN(new_n615));
  OAI21_X1  g429(.A(G478), .B1(new_n615), .B2(G902), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n599), .A2(new_n600), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n543), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n617), .B1(new_n616), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n542), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n312), .A2(new_n509), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n377), .A2(new_n379), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n471), .A2(new_n187), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n473), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n429), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  INV_X1    g445(.A(new_n311), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n308), .B2(new_n309), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n604), .A2(new_n603), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n542), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n509), .B(KEYINPUT98), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n624), .A3(new_n628), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NAND2_X1  g454(.A1(new_n401), .A2(new_n407), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n422), .A2(new_n424), .B1(new_n427), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n627), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n624), .A2(new_n605), .A3(new_n633), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT99), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n646), .B(new_n648), .ZN(G12));
  NAND2_X1  g463(.A1(new_n498), .A2(new_n500), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n380), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n506), .A2(G900), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n504), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n634), .A2(new_n542), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n644), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XNOR2_X1  g473(.A(new_n653), .B(KEYINPUT39), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT102), .B1(new_n624), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT40), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n624), .A2(new_n660), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n661), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n310), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n536), .A2(new_n538), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n540), .A2(G475), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n632), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n603), .A3(new_n604), .ZN(new_n675));
  INV_X1    g489(.A(new_n463), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n462), .B1(new_n483), .B2(new_n430), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n272), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n466), .A3(new_n439), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n485), .A2(new_n459), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(KEYINPUT101), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n187), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT101), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n475), .A2(new_n476), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n644), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n671), .A2(new_n675), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n664), .A2(new_n669), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  NOR3_X1   g503(.A1(new_n622), .A2(new_n644), .A3(new_n654), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n651), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OAI21_X1  g506(.A(new_n187), .B1(new_n366), .B2(new_n367), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n368), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n378), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n623), .A2(new_n501), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND3_X1  g513(.A1(new_n501), .A2(new_n637), .A3(new_n696), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n696), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n312), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n650), .A3(new_n605), .A4(new_n656), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  NOR2_X1   g520(.A1(G472), .A2(G902), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n486), .A2(new_n443), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n486), .A2(new_n710), .A3(new_n443), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n466), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n679), .A2(new_n469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n465), .A2(KEYINPUT31), .A3(new_n466), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n706), .B(new_n707), .C1(new_n712), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n626), .ZN(new_n718));
  INV_X1    g532(.A(new_n711), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n710), .B1(new_n486), .B2(new_n443), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n459), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n715), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n706), .B1(new_n722), .B2(new_n707), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n428), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n636), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n702), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n675), .B1(new_n308), .B2(new_n309), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NAND2_X1  g545(.A1(new_n616), .A2(new_n619), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT97), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n541), .B(new_n654), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n696), .A2(new_n735), .A3(new_n633), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n724), .B2(new_n656), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n718), .A2(new_n723), .A3(new_n644), .A4(KEYINPUT105), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  AND3_X1   g555(.A1(new_n308), .A2(new_n311), .A3(new_n309), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n378), .B1(new_n368), .B2(new_n373), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n735), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n476), .A2(KEYINPUT106), .ZN(new_n745));
  AOI21_X1  g559(.A(G902), .B1(new_n715), .B2(new_n460), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT32), .A4(new_n472), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n748), .A3(new_n475), .A4(new_n496), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT42), .A3(new_n428), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n308), .A2(new_n311), .A3(new_n309), .ZN(new_n752));
  INV_X1    g566(.A(new_n743), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n650), .A2(new_n428), .A3(new_n735), .A4(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n323), .ZN(G33));
  NAND3_X1  g572(.A1(new_n501), .A2(new_n655), .A3(new_n754), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  NOR2_X1   g574(.A1(new_n620), .A2(new_n621), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT43), .B1(new_n761), .B2(new_n542), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n644), .B1(new_n473), .B2(new_n626), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n733), .A2(new_n734), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n541), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n752), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT44), .A4(new_n766), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(G469), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n187), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n369), .A2(new_n363), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n370), .A2(new_n371), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT45), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n372), .A2(KEYINPUT107), .A3(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n372), .B2(KEYINPUT45), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n774), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT108), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n774), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n784), .A2(KEYINPUT46), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n785), .A2(new_n368), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n791), .A2(new_n376), .A3(new_n660), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n772), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT110), .B(G137), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G39));
  NAND3_X1  g611(.A1(new_n742), .A2(new_n735), .A3(new_n429), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n650), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n791), .A2(KEYINPUT47), .A3(new_n376), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT47), .B1(new_n791), .B2(new_n376), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND2_X1  g618(.A1(new_n428), .A2(new_n505), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n702), .A2(new_n685), .A3(new_n752), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n542), .A3(new_n764), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n762), .A2(new_n505), .A3(new_n766), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n725), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n703), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n502), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n808), .A2(new_n702), .A3(new_n752), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n749), .A2(new_n428), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n813), .A2(KEYINPUT48), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT48), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n811), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n671), .A2(new_n632), .A3(new_n696), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n818), .A2(KEYINPUT50), .A3(new_n809), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT50), .B1(new_n818), .B2(new_n809), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n812), .B1(new_n739), .B2(new_n738), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n806), .A2(new_n541), .A3(new_n761), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n809), .A2(new_n742), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT116), .ZN(new_n828));
  INV_X1    g642(.A(new_n802), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(new_n800), .C1(new_n376), .C2(new_n695), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n817), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(KEYINPUT117), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n821), .A3(new_n825), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n753), .A2(new_n654), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n729), .A3(new_n644), .A4(new_n685), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n380), .B(new_n650), .C1(new_n657), .C2(new_n690), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n740), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT113), .A4(new_n740), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n740), .A3(new_n842), .ZN(new_n850));
  XNOR2_X1  g664(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n601), .A2(new_n602), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n541), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n727), .B1(new_n622), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n624), .A2(new_n633), .A3(new_n628), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n650), .A2(new_n428), .ZN(new_n858));
  INV_X1    g672(.A(new_n377), .ZN(new_n859));
  INV_X1    g673(.A(new_n379), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n605), .A4(new_n633), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n646), .B(new_n857), .C1(new_n858), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n606), .A2(KEYINPUT112), .A3(new_n646), .A4(new_n857), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n697), .A2(new_n704), .A3(new_n730), .A4(new_n700), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n742), .A2(new_n735), .A3(new_n743), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n738), .B2(new_n739), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n541), .A2(new_n653), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n752), .A2(new_n854), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n650), .A2(new_n871), .A3(new_n624), .A4(new_n656), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n759), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n757), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n853), .A2(new_n875), .A3(KEYINPUT53), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n850), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n845), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n840), .B1(new_n884), .B2(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n876), .A2(new_n883), .A3(KEYINPUT115), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n880), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n847), .A2(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n877), .B1(new_n889), .B2(new_n882), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n839), .A2(new_n885), .A3(new_n887), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n428), .A2(new_n311), .A3(new_n376), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT111), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n896), .A2(new_n542), .A3(new_n761), .A4(new_n685), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n695), .B(KEYINPUT49), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n671), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G75));
  AOI21_X1  g714(.A(KEYINPUT53), .B1(new_n875), .B2(new_n880), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n889), .A2(new_n882), .A3(new_n877), .ZN(new_n902));
  OAI211_X1 g716(.A(G210), .B(G902), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n295), .A2(new_n299), .A3(new_n302), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n300), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n338), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT118), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n903), .A2(new_n904), .ZN(new_n914));
  INV_X1    g728(.A(new_n907), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n908), .A4(new_n910), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n913), .A2(new_n918), .ZN(G51));
  XNOR2_X1  g733(.A(new_n884), .B(new_n886), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n774), .B(KEYINPUT57), .Z(new_n921));
  OAI22_X1  g735(.A1(new_n920), .A2(new_n921), .B1(new_n367), .B2(new_n366), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n187), .B1(new_n876), .B2(new_n883), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n788), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n909), .B1(new_n922), .B2(new_n924), .ZN(G54));
  OR2_X1    g739(.A1(new_n529), .A2(new_n534), .ZN(new_n926));
  AND2_X1   g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n923), .B2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n909), .ZN(G60));
  INV_X1    g744(.A(new_n615), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n885), .A2(new_n887), .A3(new_n892), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT59), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n910), .B1(new_n920), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(G63));
  XNOR2_X1  g752(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n381), .A2(new_n187), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n884), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n643), .B(KEYINPUT120), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n909), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(KEYINPUT61), .C1(new_n426), .C2(new_n942), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n942), .A2(new_n426), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n884), .A2(new_n941), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n910), .B1(new_n949), .B2(new_n943), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n947), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G66));
  AND2_X1   g766(.A1(new_n866), .A2(new_n867), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n338), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n508), .B2(new_n213), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n905), .B1(G898), .B2(new_n338), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n956), .B2(new_n338), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G69));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n729), .A2(new_n428), .A3(new_n749), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n791), .A2(new_n968), .A3(new_n376), .A4(new_n660), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n759), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n755), .A2(new_n756), .ZN(new_n971));
  INV_X1    g785(.A(new_n751), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n844), .A2(new_n740), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n803), .A2(new_n970), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n967), .B1(new_n976), .B2(new_n795), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n829), .A2(new_n800), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n974), .B1(new_n978), .B2(new_n799), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n973), .A2(new_n759), .A3(new_n969), .ZN(new_n980));
  INV_X1    g794(.A(new_n794), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n772), .A3(new_n792), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT123), .A4(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n977), .A2(new_n983), .A3(new_n338), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n464), .B(new_n532), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(G900), .B2(G953), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n622), .A2(new_n855), .ZN(new_n988));
  OR4_X1    g802(.A1(new_n858), .A2(new_n665), .A3(new_n988), .A4(new_n752), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n803), .B(new_n989), .C1(new_n793), .C2(new_n794), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n688), .A2(new_n975), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n688), .A2(KEYINPUT62), .A3(new_n975), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n985), .B1(new_n995), .B2(G953), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n987), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n338), .B1(G227), .B2(G900), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n966), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  AOI211_X1 g816(.A(KEYINPUT125), .B(new_n1000), .C1(new_n987), .C2(new_n996), .ZN(new_n1003));
  INV_X1    g817(.A(new_n998), .ZN(new_n1004));
  OAI22_X1  g818(.A1(new_n1002), .A2(new_n1003), .B1(KEYINPUT124), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n990), .ZN(new_n1006));
  INV_X1    g820(.A(new_n994), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT62), .B1(new_n688), .B2(new_n975), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n338), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n1010), .A2(new_n985), .B1(new_n984), .B2(new_n986), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT125), .B1(new_n1011), .B2(new_n1000), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1004), .A2(KEYINPUT124), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n997), .A2(new_n966), .A3(new_n1001), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1005), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT126), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n956), .B2(new_n1009), .ZN(new_n1021));
  INV_X1    g835(.A(new_n465), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1021), .A2(KEYINPUT127), .A3(new_n466), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n953), .B(KEYINPUT121), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1019), .B1(new_n1025), .B2(new_n995), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1022), .A2(new_n466), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n465), .A2(new_n459), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n977), .B(new_n983), .C1(new_n954), .C2(new_n955), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n1020), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n491), .A2(new_n679), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n891), .A2(new_n1018), .A3(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1032), .A2(new_n1034), .A3(new_n909), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n1029), .A2(new_n1035), .ZN(G57));
endmodule


