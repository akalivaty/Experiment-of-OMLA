//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT34), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G15gat), .B(G43gat), .Z(new_n206));
  XNOR2_X1  g005(.A(G71gat), .B(G99gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G227gat), .ZN(new_n209));
  INV_X1    g008(.A(G233gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(new_n214), .B2(new_n215), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n220), .A2(KEYINPUT28), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  OAI221_X1 g022(.A(new_n213), .B1(new_n218), .B2(new_n219), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n225), .A2(G169gat), .A3(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT23), .B1(new_n214), .B2(new_n215), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(new_n216), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(new_n221), .A3(KEYINPUT67), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(new_n232), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n236), .A3(KEYINPUT25), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n221), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n230), .A4(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n238), .B1(new_n228), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n237), .B1(new_n244), .B2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  AOI211_X1 g045(.A(new_n246), .B(new_n238), .C1(new_n228), .C2(new_n243), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n224), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249));
  INV_X1    g048(.A(G127gat), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(G134gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(G134gat), .ZN(new_n252));
  OAI22_X1  g051(.A1(new_n249), .A2(KEYINPUT1), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G113gat), .ZN(new_n255));
  INV_X1    g054(.A(G113gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G127gat), .B(G134gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n248), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n224), .C1(new_n245), .C2(new_n247), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n212), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n208), .B1(new_n266), .B2(KEYINPUT33), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT32), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n263), .A2(new_n265), .ZN(new_n271));
  AOI221_X4 g070(.A(new_n268), .B1(KEYINPUT33), .B2(new_n208), .C1(new_n271), .C2(new_n211), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n205), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n267), .A2(new_n269), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n275), .A2(new_n272), .A3(new_n204), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n263), .A2(new_n212), .A3(new_n265), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n202), .A2(new_n203), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n274), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n273), .A3(new_n205), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n204), .B1(new_n275), .B2(new_n272), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286));
  XNOR2_X1  g085(.A(G1gat), .B(G29gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT0), .ZN(new_n288));
  XNOR2_X1  g087(.A(G57gat), .B(G85gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  XNOR2_X1  g089(.A(G141gat), .B(G148gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(KEYINPUT2), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n292), .A3(KEYINPUT2), .ZN(new_n296));
  AND2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT74), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n293), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n295), .A2(new_n296), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n297), .A2(new_n298), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n293), .A2(KEYINPUT2), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n306), .A2(new_n308), .A3(new_n291), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT3), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n311));
  AND2_X1   g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n296), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n304), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n306), .A2(new_n291), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n307), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n310), .A2(new_n321), .A3(new_n262), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n319), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n262), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n316), .A2(new_n315), .B1(new_n318), .B2(new_n307), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n264), .A3(KEYINPUT4), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n322), .A2(new_n325), .A3(new_n327), .A4(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n324), .A2(new_n323), .A3(new_n262), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT4), .B1(new_n326), .B2(new_n264), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(KEYINPUT78), .A3(new_n322), .A4(new_n331), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n305), .A2(new_n262), .A3(new_n309), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n317), .A2(new_n319), .B1(new_n261), .B2(new_n253), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n330), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n322), .A2(new_n325), .A3(new_n327), .A4(new_n329), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n345), .B(new_n330), .C1(new_n340), .C2(new_n341), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n343), .A2(new_n344), .A3(new_n328), .A4(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n290), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT6), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n339), .A2(new_n290), .A3(new_n347), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n348), .B1(new_n353), .B2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n358));
  NAND2_X1  g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G211gat), .B(G218gat), .Z(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G211gat), .B(G218gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT71), .ZN(new_n366));
  INV_X1    g165(.A(G197gat), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(G204gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n359), .A2(new_n358), .A3(new_n360), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(G204gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT71), .B(new_n365), .C1(new_n371), .C2(new_n361), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n228), .A2(new_n243), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n246), .B1(new_n376), .B2(new_n238), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n237), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n381), .B(KEYINPUT72), .Z(new_n382));
  AOI22_X1  g181(.A1(new_n379), .A2(new_n224), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n382), .B(new_n224), .C1(new_n245), .C2(new_n247), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n375), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n382), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n248), .B1(KEYINPUT29), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n375), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n384), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND3_X1  g192(.A1(new_n386), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT73), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n386), .A2(new_n390), .A3(KEYINPUT73), .A4(new_n393), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n386), .B2(new_n390), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n383), .A2(new_n385), .A3(new_n375), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n389), .B1(new_n388), .B2(new_n384), .ZN(new_n402));
  INV_X1    g201(.A(new_n393), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n404), .B2(KEYINPUT30), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n286), .B1(new_n357), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n399), .A2(new_n405), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n351), .A2(new_n355), .A3(new_n352), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n355), .B1(new_n351), .B2(new_n352), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n409), .A2(new_n410), .A3(new_n348), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT80), .B(new_n408), .C1(new_n411), .C2(new_n350), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n413), .B(KEYINPUT82), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n321), .A2(new_n380), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n415), .A2(new_n375), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n373), .A2(new_n374), .A3(new_n380), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n326), .B1(new_n417), .B2(new_n320), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n375), .ZN(new_n420));
  INV_X1    g219(.A(new_n413), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n420), .B(new_n421), .C1(new_n418), .C2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n418), .A2(new_n422), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G22gat), .ZN(new_n426));
  INV_X1    g225(.A(G22gat), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n419), .B(new_n427), .C1(new_n423), .C2(new_n424), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(KEYINPUT85), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(KEYINPUT85), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(new_n428), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n431), .B(KEYINPUT81), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT84), .B(new_n437), .C1(new_n426), .C2(new_n428), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n433), .A2(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n285), .A2(new_n407), .A3(new_n412), .A4(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n280), .B1(new_n274), .B2(new_n276), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n282), .A2(new_n283), .A3(new_n279), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n348), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n352), .A3(new_n351), .ZN(new_n448));
  AOI211_X1 g247(.A(KEYINPUT35), .B(new_n406), .C1(new_n349), .C2(new_n448), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n442), .A2(KEYINPUT35), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n322), .A2(new_n325), .A3(new_n327), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n330), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n329), .B1(new_n337), .B2(new_n322), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n340), .A2(new_n341), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT39), .B1(new_n455), .B2(new_n330), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n453), .B(new_n290), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT87), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT86), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n406), .A3(new_n447), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n386), .A2(new_n467), .A3(new_n390), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n386), .A2(new_n390), .A3(KEYINPUT89), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n467), .B1(new_n402), .B2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n386), .A2(new_n474), .A3(new_n390), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n393), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n467), .B1(new_n386), .B2(new_n390), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n479), .A2(new_n478), .A3(new_n393), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n477), .A2(new_n478), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n448), .A2(new_n349), .A3(new_n396), .A4(new_n398), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n441), .B(new_n466), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT69), .B(KEYINPUT36), .Z(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n281), .B2(new_n284), .ZN(new_n485));
  NOR2_X1   g284(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n443), .A2(new_n444), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n441), .B1(new_n407), .B2(new_n412), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n450), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G43gat), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n492), .A2(G50gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT15), .B1(new_n492), .B2(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OR3_X1    g297(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT15), .B1(new_n493), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT91), .B1(new_n492), .B2(G50gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n493), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n496), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n495), .A2(new_n502), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT16), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(G1gat), .B2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n518), .B(G8gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT92), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n503), .A2(KEYINPUT17), .A3(new_n510), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n513), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n526), .A2(KEYINPUT93), .B1(new_n511), .B2(new_n523), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT95), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT95), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n511), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n520), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n511), .A2(new_n523), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(KEYINPUT94), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(KEYINPUT94), .B2(new_n538), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n529), .B(KEYINPUT13), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT18), .A4(new_n529), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G197gat), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT11), .B(G169gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT12), .Z(new_n549));
  NOR2_X1   g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n531), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n542), .A3(new_n543), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n535), .A2(new_n550), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n556), .B2(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n561), .B2(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n555), .B(KEYINPUT98), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n559), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n570));
  AND2_X1   g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G127gat), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n523), .B1(new_n569), .B2(KEYINPUT21), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT99), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n300), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n513), .A2(new_n525), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n511), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n597), .A2(new_n598), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n599), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n583), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n569), .A2(new_n592), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n564), .A2(new_n568), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n569), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n611), .ZN(new_n618));
  INV_X1    g417(.A(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n617), .A2(new_n620), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR4_X1   g429(.A1(new_n491), .A2(new_n553), .A3(new_n608), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n357), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G1gat), .ZN(G1324gat));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n406), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n631), .A2(KEYINPUT42), .A3(new_n406), .A4(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(G8gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n631), .A2(new_n642), .A3(new_n285), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n443), .A2(new_n444), .A3(new_n486), .ZN(new_n644));
  INV_X1    g443(.A(new_n484), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n443), .B2(new_n444), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n643), .B1(new_n650), .B2(new_n642), .ZN(G1326gat));
  INV_X1    g450(.A(new_n441), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n407), .A2(new_n412), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT35), .B1(new_n657), .B2(new_n445), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n446), .A2(new_n449), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n652), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n647), .A3(new_n483), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n607), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n583), .A2(new_n553), .A3(new_n630), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n357), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n665), .A2(G29gat), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT45), .Z(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(KEYINPUT44), .C1(new_n491), .C2(new_n607), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n647), .B(new_n483), .C1(new_n489), .C2(KEYINPUT104), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n489), .A2(KEYINPUT104), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n660), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n669), .A3(new_n606), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n664), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n666), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n668), .A2(new_n679), .ZN(G1328gat));
  OAI21_X1  g479(.A(G36gat), .B1(new_n678), .B2(new_n408), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n665), .A2(G36gat), .A3(new_n408), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT46), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1329gat));
  NAND4_X1  g483(.A1(new_n677), .A2(G43gat), .A3(new_n648), .A4(new_n664), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n443), .A2(new_n444), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n492), .B1(new_n665), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT106), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(KEYINPUT106), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(G1330gat));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n652), .A3(new_n664), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G50gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n441), .A2(G50gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n663), .A2(new_n664), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(KEYINPUT48), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n663), .A2(new_n701), .A3(new_n664), .A4(new_n697), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n695), .B2(G50gat), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT48), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n699), .B1(new_n707), .B2(new_n710), .ZN(G1331gat));
  INV_X1    g510(.A(new_n675), .ZN(new_n712));
  INV_X1    g511(.A(new_n534), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n550), .A2(new_n532), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n552), .A2(new_n549), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n630), .ZN(new_n717));
  NOR4_X1   g516(.A1(new_n712), .A2(new_n716), .A3(new_n608), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n357), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n406), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  NAND2_X1  g523(.A1(new_n718), .A2(new_n648), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n686), .A2(G71gat), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n725), .A2(G71gat), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n718), .A2(new_n652), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n583), .A2(new_n716), .A3(new_n717), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n677), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n666), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n583), .A2(new_n716), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n675), .A2(new_n606), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n357), .A2(new_n587), .A3(new_n630), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(G1336gat));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n408), .A2(G92gat), .A3(new_n717), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G92gat), .B1(new_n733), .B2(new_n408), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n733), .B2(new_n647), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n686), .A2(G99gat), .A3(new_n717), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n739), .B2(new_n749), .ZN(G1338gat));
  OAI21_X1  g549(.A(G106gat), .B1(new_n733), .B2(new_n441), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n441), .A2(G106gat), .A3(new_n717), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n738), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n540), .A2(new_n541), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n529), .B1(new_n527), .B2(new_n528), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n548), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n714), .A2(new_n630), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n617), .A2(KEYINPUT54), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n619), .B1(new_n613), .B2(new_n614), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n628), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(KEYINPUT55), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n629), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT55), .B1(new_n762), .B2(new_n765), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n760), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n768), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(KEYINPUT111), .A3(new_n629), .A4(new_n766), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n759), .B1(new_n772), .B2(new_n553), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n607), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT112), .B1(new_n714), .B2(new_n758), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n771), .A3(new_n606), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n714), .A2(KEYINPUT112), .A3(new_n758), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n583), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n583), .A2(new_n553), .A3(new_n607), .A4(new_n717), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n357), .B(new_n446), .C1(new_n781), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n406), .B1(new_n784), .B2(KEYINPUT113), .ZN(new_n785));
  INV_X1    g584(.A(new_n583), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n716), .A2(new_n769), .A3(new_n771), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n606), .B1(new_n787), .B2(new_n759), .ZN(new_n788));
  INV_X1    g587(.A(new_n779), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(new_n775), .A3(new_n777), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n445), .B1(new_n791), .B2(new_n782), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n357), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n785), .A2(new_n716), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n784), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n408), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n716), .A2(G113gat), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n795), .A2(G113gat), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT114), .ZN(G1340gat));
  OAI21_X1  g599(.A(G120gat), .B1(new_n797), .B2(new_n717), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n630), .A2(new_n254), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT115), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n794), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1341gat));
  NAND4_X1  g604(.A1(new_n796), .A2(G127gat), .A3(new_n408), .A4(new_n583), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n583), .A3(new_n794), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n250), .B2(new_n808), .ZN(G1342gat));
  NOR2_X1   g608(.A1(new_n607), .A2(G134gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n794), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n785), .A2(KEYINPUT117), .A3(new_n794), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT56), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n813), .A2(new_n819), .A3(new_n814), .ZN(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n797), .B2(new_n607), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n815), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  NOR3_X1   g623(.A1(new_n648), .A2(new_n666), .A3(new_n406), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n441), .B1(new_n791), .B2(new_n782), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n652), .A2(KEYINPUT57), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n767), .A2(new_n768), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n716), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n606), .B1(new_n829), .B2(new_n759), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n786), .B1(new_n790), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n827), .B1(new_n831), .B2(new_n782), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n826), .A2(KEYINPUT57), .B1(new_n832), .B2(KEYINPUT119), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n832), .A2(KEYINPUT119), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n825), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n716), .A2(G141gat), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(G141gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n652), .B1(new_n781), .B2(new_n783), .ZN(new_n839));
  INV_X1    g638(.A(new_n825), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n553), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n837), .A2(KEYINPUT58), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1344gat));
  INV_X1    g647(.A(G148gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n841), .A2(new_n849), .A3(new_n630), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(KEYINPUT59), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n835), .B2(new_n717), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n441), .A2(KEYINPUT57), .ZN(new_n855));
  INV_X1    g654(.A(new_n830), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n828), .A2(new_n606), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT121), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(KEYINPUT121), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n776), .A3(new_n779), .A4(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n583), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n855), .B1(new_n861), .B2(new_n783), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n630), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G148gat), .B1(new_n863), .B2(new_n840), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT59), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n853), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n850), .B1(new_n866), .B2(new_n867), .ZN(G1345gat));
  OAI21_X1  g667(.A(G155gat), .B1(new_n835), .B2(new_n786), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n300), .A3(new_n583), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n835), .B2(new_n607), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n841), .A2(new_n301), .A3(new_n606), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(KEYINPUT122), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n357), .A2(new_n408), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n792), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n553), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(new_n214), .ZN(G1348gat));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n717), .ZN(new_n883));
  XOR2_X1   g682(.A(KEYINPUT123), .B(G176gat), .Z(new_n884));
  XNOR2_X1  g683(.A(new_n883), .B(new_n884), .ZN(G1349gat));
  NAND3_X1  g684(.A1(new_n792), .A2(new_n583), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n231), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n220), .B2(new_n886), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g688(.A1(new_n792), .A2(new_n606), .A3(new_n879), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(G190gat), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT124), .Z(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(G190gat), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT61), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(KEYINPUT61), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(G1351gat));
  NAND2_X1  g696(.A1(new_n647), .A2(new_n879), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n826), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n367), .B1(new_n900), .B2(new_n553), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n854), .A2(new_n862), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n716), .A2(G197gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT125), .ZN(G1352gat));
  NOR3_X1   g705(.A1(new_n900), .A2(G204gat), .A3(new_n717), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT62), .ZN(new_n908));
  OAI21_X1  g707(.A(G204gat), .B1(new_n863), .B2(new_n898), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1353gat));
  OR3_X1    g709(.A1(new_n900), .A2(G211gat), .A3(new_n786), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n583), .A3(new_n899), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT63), .B1(new_n912), .B2(G211gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(G1354gat));
  NAND2_X1  g715(.A1(new_n606), .A2(G218gat), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT126), .Z(new_n918));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n607), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n903), .A2(new_n918), .B1(G218gat), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(G1355gat));
endmodule


