

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n561), .B(n560), .ZN(n677) );
  AND2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n915) );
  BUF_X4 U557 ( .A(n764), .Z(n521) );
  XNOR2_X1 U558 ( .A(n714), .B(KEYINPUT64), .ZN(n764) );
  AND2_X1 U559 ( .A1(n713), .A2(n712), .ZN(n801) );
  XNOR2_X1 U560 ( .A(n585), .B(n584), .ZN(n709) );
  XNOR2_X1 U561 ( .A(n550), .B(n549), .ZN(n598) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n550) );
  XNOR2_X1 U563 ( .A(n535), .B(KEYINPUT102), .ZN(n534) );
  INV_X1 U564 ( .A(n543), .ZN(n538) );
  OR2_X1 U565 ( .A1(n544), .A2(n762), .ZN(n542) );
  OR2_X1 U566 ( .A1(n758), .A2(n745), .ZN(n748) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n532) );
  NOR2_X1 U568 ( .A1(n524), .A2(n761), .ZN(n543) );
  NOR2_X1 U569 ( .A1(G1966), .A2(n800), .ZN(n758) );
  NAND2_X1 U570 ( .A1(n539), .A2(n536), .ZN(n780) );
  AND2_X1 U571 ( .A1(n542), .A2(n540), .ZN(n539) );
  XNOR2_X1 U572 ( .A(n553), .B(KEYINPUT66), .ZN(n596) );
  NOR2_X1 U573 ( .A1(n554), .A2(G2104), .ZN(n553) );
  NOR2_X2 U574 ( .A1(G651), .A2(G543), .ZN(n672) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n559), .Z(n673) );
  NAND2_X1 U576 ( .A1(n599), .A2(G101), .ZN(n585) );
  XOR2_X1 U577 ( .A(KEYINPUT7), .B(n573), .Z(n522) );
  XOR2_X1 U578 ( .A(n722), .B(n721), .Z(n523) );
  NAND2_X1 U579 ( .A1(n756), .A2(n755), .ZN(n763) );
  AND2_X1 U580 ( .A1(n758), .A2(n547), .ZN(n524) );
  INV_X1 U581 ( .A(G2105), .ZN(n554) );
  AND2_X1 U582 ( .A1(n546), .A2(n537), .ZN(n525) );
  NOR2_X1 U583 ( .A1(n758), .A2(n547), .ZN(n526) );
  OR2_X1 U584 ( .A1(n800), .A2(n799), .ZN(n527) );
  AND2_X1 U585 ( .A1(n845), .A2(n835), .ZN(n528) );
  XNOR2_X1 U586 ( .A(n529), .B(KEYINPUT113), .ZN(n837) );
  NAND2_X1 U587 ( .A1(n530), .A2(n528), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n531), .A2(n527), .ZN(n530) );
  XNOR2_X1 U589 ( .A(n797), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n533), .B(n532), .ZN(n743) );
  NAND2_X1 U591 ( .A1(n534), .A2(n523), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n736), .A2(n737), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n544), .A2(n525), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n538), .A2(KEYINPUT108), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n541), .A2(KEYINPUT108), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n546), .A2(n543), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n545), .A2(n526), .ZN(n544) );
  INV_X1 U598 ( .A(n759), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n759), .A2(n547), .ZN(n546) );
  INV_X1 U600 ( .A(KEYINPUT107), .ZN(n547) );
  BUF_X1 U601 ( .A(n598), .Z(n912) );
  XOR2_X1 U602 ( .A(KEYINPUT74), .B(n622), .Z(n548) );
  NOR2_X1 U603 ( .A1(n521), .A2(n972), .ZN(n717) );
  XNOR2_X1 U604 ( .A(n746), .B(KEYINPUT104), .ZN(n747) );
  NOR2_X1 U605 ( .A1(n749), .A2(G168), .ZN(n750) );
  INV_X1 U606 ( .A(KEYINPUT106), .ZN(n757) );
  NAND2_X1 U607 ( .A1(n803), .A2(n801), .ZN(n714) );
  NAND2_X1 U608 ( .A1(n521), .A2(G8), .ZN(n800) );
  AND2_X1 U609 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U610 ( .A1(n677), .A2(G51), .ZN(n562) );
  INV_X1 U611 ( .A(KEYINPUT17), .ZN(n549) );
  INV_X1 U612 ( .A(KEYINPUT65), .ZN(n560) );
  XNOR2_X1 U613 ( .A(n626), .B(KEYINPUT15), .ZN(n998) );
  INV_X1 U614 ( .A(KEYINPUT23), .ZN(n584) );
  XNOR2_X1 U615 ( .A(KEYINPUT76), .B(n522), .ZN(G168) );
  NAND2_X1 U616 ( .A1(G138), .A2(n598), .ZN(n552) );
  AND2_X4 U617 ( .A1(n554), .A2(G2104), .ZN(n599) );
  NAND2_X1 U618 ( .A1(G102), .A2(n599), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n596), .A2(G126), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n915), .A2(G114), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(G164) );
  INV_X1 U624 ( .A(G651), .ZN(n567) );
  NOR2_X1 U625 ( .A1(G543), .A2(n567), .ZN(n559) );
  NAND2_X1 U626 ( .A1(G63), .A2(n673), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT0), .B(G543), .Z(n653) );
  NOR2_X1 U628 ( .A1(G651), .A2(n653), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT6), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G89), .A2(n672), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT75), .B(n565), .Z(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT4), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n653), .A2(n567), .ZN(n676) );
  NAND2_X1 U635 ( .A1(G76), .A2(n676), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(n570), .B(KEYINPUT5), .Z(n571) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n677), .A2(G52), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT70), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G64), .A2(n673), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n672), .A2(G90), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT71), .B(n577), .Z(n579) );
  NAND2_X1 U645 ( .A1(n676), .A2(G77), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(n580), .Z(n581) );
  NOR2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(KEYINPUT72), .B(n583), .ZN(G171) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(n598), .A2(G137), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G113), .A2(n915), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n588), .B(KEYINPUT67), .ZN(n712) );
  NAND2_X1 U655 ( .A1(G125), .A2(n596), .ZN(n711) );
  AND2_X1 U656 ( .A1(n712), .A2(n711), .ZN(n589) );
  AND2_X1 U657 ( .A1(n709), .A2(n589), .ZN(G160) );
  NAND2_X1 U658 ( .A1(G91), .A2(n672), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G65), .A2(n673), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G78), .A2(n676), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G53), .A2(n677), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  OR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G299) );
  BUF_X1 U665 ( .A(n596), .Z(n916) );
  NAND2_X1 U666 ( .A1(n916), .A2(G123), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U668 ( .A1(G135), .A2(n912), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G99), .A2(n599), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n915), .A2(G111), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT78), .B(n602), .Z(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n954) );
  XNOR2_X1 U675 ( .A(G2096), .B(n954), .ZN(n607) );
  OR2_X1 U676 ( .A1(G2100), .A2(n607), .ZN(G156) );
  INV_X1 U677 ( .A(G120), .ZN(G236) );
  NAND2_X1 U678 ( .A1(G94), .A2(G452), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U680 ( .A1(G7), .A2(G661), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U682 ( .A(G223), .ZN(n853) );
  NAND2_X1 U683 ( .A1(n853), .A2(G567), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT11), .B(n610), .Z(G234) );
  NAND2_X1 U685 ( .A1(G56), .A2(n673), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT14), .B(n611), .Z(n617) );
  NAND2_X1 U687 ( .A1(n672), .A2(G81), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G68), .A2(n676), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U691 ( .A(KEYINPUT13), .B(n615), .Z(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n677), .A2(G43), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n999) );
  INV_X1 U695 ( .A(G860), .ZN(n631) );
  OR2_X1 U696 ( .A1(n999), .A2(n631), .ZN(G153) );
  NAND2_X1 U697 ( .A1(G301), .A2(G868), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G54), .A2(n677), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G79), .A2(n676), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G66), .A2(n673), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n672), .A2(G92), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n623), .A2(n548), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U705 ( .A1(n998), .A2(G868), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(G284) );
  XOR2_X1 U707 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U708 ( .A1(G868), .A2(G286), .ZN(n630) );
  INV_X1 U709 ( .A(G868), .ZN(n691) );
  NAND2_X1 U710 ( .A1(G299), .A2(n691), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(G297) );
  NAND2_X1 U712 ( .A1(n631), .A2(G559), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n632), .A2(n998), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n633), .B(KEYINPUT16), .ZN(n634) );
  XOR2_X1 U715 ( .A(KEYINPUT77), .B(n634), .Z(G148) );
  NOR2_X1 U716 ( .A1(G868), .A2(n999), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G868), .A2(n998), .ZN(n635) );
  NOR2_X1 U718 ( .A1(G559), .A2(n635), .ZN(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G282) );
  NAND2_X1 U720 ( .A1(G85), .A2(n672), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(KEYINPUT68), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n673), .A2(G60), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G72), .A2(n676), .ZN(n641) );
  XNOR2_X1 U725 ( .A(KEYINPUT69), .B(n641), .ZN(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n677), .A2(G47), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G75), .A2(n676), .ZN(n646) );
  XNOR2_X1 U730 ( .A(n646), .B(KEYINPUT86), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n672), .A2(G88), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G62), .A2(n673), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G50), .A2(n677), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U736 ( .A1(n652), .A2(n651), .ZN(G166) );
  INV_X1 U737 ( .A(G166), .ZN(G303) );
  NAND2_X1 U738 ( .A1(n653), .A2(G87), .ZN(n654) );
  XNOR2_X1 U739 ( .A(KEYINPUT82), .B(n654), .ZN(n660) );
  NAND2_X1 U740 ( .A1(G49), .A2(n677), .ZN(n656) );
  NAND2_X1 U741 ( .A1(G74), .A2(G651), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U743 ( .A1(n673), .A2(n657), .ZN(n658) );
  XOR2_X1 U744 ( .A(KEYINPUT81), .B(n658), .Z(n659) );
  NAND2_X1 U745 ( .A1(n660), .A2(n659), .ZN(G288) );
  XOR2_X1 U746 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n662) );
  NAND2_X1 U747 ( .A1(G73), .A2(n676), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n662), .B(n661), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n673), .A2(G61), .ZN(n663) );
  XNOR2_X1 U750 ( .A(KEYINPUT83), .B(n663), .ZN(n664) );
  NOR2_X1 U751 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n672), .A2(G86), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(KEYINPUT85), .ZN(n670) );
  NAND2_X1 U755 ( .A1(G48), .A2(n677), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n670), .A2(n669), .ZN(G305) );
  NAND2_X1 U757 ( .A1(G559), .A2(n998), .ZN(n671) );
  XOR2_X1 U758 ( .A(n999), .B(n671), .Z(n857) );
  XOR2_X1 U759 ( .A(KEYINPUT88), .B(KEYINPUT19), .Z(n684) );
  NAND2_X1 U760 ( .A1(G93), .A2(n672), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G67), .A2(n673), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G80), .A2(n676), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G55), .A2(n677), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U766 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U767 ( .A(KEYINPUT80), .B(n682), .Z(n860) );
  XNOR2_X1 U768 ( .A(n860), .B(KEYINPUT87), .ZN(n683) );
  XNOR2_X1 U769 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(G299), .ZN(n688) );
  XNOR2_X1 U771 ( .A(G290), .B(G303), .ZN(n686) );
  XNOR2_X1 U772 ( .A(n686), .B(G288), .ZN(n687) );
  XNOR2_X1 U773 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U774 ( .A(n689), .B(G305), .ZN(n926) );
  XNOR2_X1 U775 ( .A(n857), .B(n926), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n690), .A2(G868), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n691), .A2(n860), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n693), .A2(n692), .ZN(G295) );
  NAND2_X1 U779 ( .A1(G2084), .A2(G2078), .ZN(n694) );
  XOR2_X1 U780 ( .A(KEYINPUT20), .B(n694), .Z(n695) );
  NAND2_X1 U781 ( .A1(G2090), .A2(n695), .ZN(n696) );
  XNOR2_X1 U782 ( .A(KEYINPUT21), .B(n696), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n697), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U784 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U785 ( .A1(G69), .A2(G57), .ZN(n698) );
  NOR2_X1 U786 ( .A1(G236), .A2(n698), .ZN(n699) );
  XNOR2_X1 U787 ( .A(KEYINPUT90), .B(n699), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n700), .A2(G108), .ZN(n861) );
  NAND2_X1 U789 ( .A1(n861), .A2(G567), .ZN(n706) );
  XOR2_X1 U790 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n702) );
  NAND2_X1 U791 ( .A1(G132), .A2(G82), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U793 ( .A1(n703), .A2(G218), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G96), .A2(n704), .ZN(n862) );
  NAND2_X1 U795 ( .A1(n862), .A2(G2106), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n863) );
  NAND2_X1 U797 ( .A1(G483), .A2(G661), .ZN(n707) );
  NOR2_X1 U798 ( .A1(n863), .A2(n707), .ZN(n856) );
  NAND2_X1 U799 ( .A1(n856), .A2(G36), .ZN(G176) );
  NOR2_X1 U800 ( .A1(G164), .A2(G1384), .ZN(n803) );
  AND2_X1 U801 ( .A1(G40), .A2(n709), .ZN(n710) );
  INV_X1 U802 ( .A(n800), .ZN(n788) );
  INV_X1 U803 ( .A(G2072), .ZN(n972) );
  XOR2_X1 U804 ( .A(KEYINPUT99), .B(KEYINPUT27), .Z(n715) );
  XNOR2_X1 U805 ( .A(KEYINPUT98), .B(n715), .ZN(n716) );
  XNOR2_X1 U806 ( .A(n717), .B(n716), .ZN(n720) );
  BUF_X1 U807 ( .A(n521), .Z(n718) );
  NAND2_X1 U808 ( .A1(n718), .A2(G1956), .ZN(n719) );
  NAND2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n733) );
  NAND2_X1 U810 ( .A1(G299), .A2(n733), .ZN(n722) );
  XOR2_X1 U811 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n721) );
  INV_X1 U812 ( .A(n521), .ZN(n738) );
  NAND2_X1 U813 ( .A1(G2067), .A2(n738), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n521), .A2(G1348), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U816 ( .A(n725), .B(KEYINPUT101), .ZN(n732) );
  OR2_X1 U817 ( .A1(n998), .A2(n732), .ZN(n731) );
  NAND2_X1 U818 ( .A1(n738), .A2(G1996), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n726), .B(KEYINPUT26), .ZN(n728) );
  NAND2_X1 U820 ( .A1(n521), .A2(G1341), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n999), .A2(n729), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n737) );
  AND2_X1 U824 ( .A1(n732), .A2(n998), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G299), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U827 ( .A(G2078), .B(KEYINPUT25), .Z(n971) );
  NOR2_X1 U828 ( .A1(n718), .A2(n971), .ZN(n740) );
  NOR2_X1 U829 ( .A1(G1961), .A2(n738), .ZN(n739) );
  NOR2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n751) );
  NOR2_X1 U831 ( .A1(G301), .A2(n751), .ZN(n741) );
  XNOR2_X1 U832 ( .A(KEYINPUT97), .B(n741), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n756) );
  NOR2_X1 U834 ( .A1(n521), .A2(G2084), .ZN(n760) );
  INV_X1 U835 ( .A(n760), .ZN(n744) );
  NAND2_X1 U836 ( .A1(n744), .A2(G8), .ZN(n745) );
  XOR2_X1 U837 ( .A(KEYINPUT30), .B(KEYINPUT103), .Z(n746) );
  XNOR2_X1 U838 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U839 ( .A(n750), .B(KEYINPUT105), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n751), .A2(G301), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U842 ( .A(n754), .B(KEYINPUT31), .ZN(n755) );
  XNOR2_X1 U843 ( .A(n763), .B(n757), .ZN(n759) );
  AND2_X1 U844 ( .A1(G8), .A2(n760), .ZN(n761) );
  INV_X1 U845 ( .A(KEYINPUT108), .ZN(n762) );
  NAND2_X1 U846 ( .A1(G286), .A2(n763), .ZN(n770) );
  NOR2_X1 U847 ( .A1(n521), .A2(G2090), .ZN(n765) );
  XOR2_X1 U848 ( .A(KEYINPUT109), .B(n765), .Z(n767) );
  NOR2_X1 U849 ( .A1(G1971), .A2(n800), .ZN(n766) );
  NOR2_X1 U850 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U851 ( .A1(n768), .A2(G303), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U853 ( .A1(G8), .A2(n771), .ZN(n772) );
  XNOR2_X1 U854 ( .A(KEYINPUT32), .B(n772), .ZN(n778) );
  AND2_X1 U855 ( .A1(n780), .A2(n778), .ZN(n775) );
  NAND2_X1 U856 ( .A1(G8), .A2(G166), .ZN(n773) );
  NOR2_X1 U857 ( .A1(G2090), .A2(n773), .ZN(n774) );
  NOR2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U859 ( .A1(n788), .A2(n776), .ZN(n796) );
  XNOR2_X1 U860 ( .A(G1981), .B(G305), .ZN(n996) );
  NAND2_X1 U861 ( .A1(G288), .A2(G1976), .ZN(n777) );
  XOR2_X1 U862 ( .A(KEYINPUT110), .B(n777), .Z(n1009) );
  NOR2_X1 U863 ( .A1(n800), .A2(n1009), .ZN(n781) );
  AND2_X1 U864 ( .A1(n778), .A2(n781), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n786) );
  INV_X1 U866 ( .A(KEYINPUT33), .ZN(n790) );
  INV_X1 U867 ( .A(n781), .ZN(n783) );
  NOR2_X1 U868 ( .A1(G1976), .A2(G288), .ZN(n787) );
  NOR2_X1 U869 ( .A1(G1971), .A2(G303), .ZN(n782) );
  NOR2_X1 U870 ( .A1(n787), .A2(n782), .ZN(n1007) );
  OR2_X1 U871 ( .A1(n783), .A2(n1007), .ZN(n784) );
  AND2_X1 U872 ( .A1(n790), .A2(n784), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n793) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U876 ( .A(n791), .B(KEYINPUT111), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U878 ( .A1(n996), .A2(n794), .ZN(n795) );
  NOR2_X1 U879 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XOR2_X1 U881 ( .A(n798), .B(KEYINPUT24), .Z(n799) );
  INV_X1 U882 ( .A(n801), .ZN(n802) );
  NOR2_X1 U883 ( .A1(n803), .A2(n802), .ZN(n848) );
  NAND2_X1 U884 ( .A1(n912), .A2(G140), .ZN(n804) );
  XOR2_X1 U885 ( .A(KEYINPUT91), .B(n804), .Z(n806) );
  NAND2_X1 U886 ( .A1(n599), .A2(G104), .ZN(n805) );
  NAND2_X1 U887 ( .A1(n806), .A2(n805), .ZN(n808) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n807) );
  XNOR2_X1 U889 ( .A(n808), .B(n807), .ZN(n813) );
  NAND2_X1 U890 ( .A1(n915), .A2(G116), .ZN(n810) );
  NAND2_X1 U891 ( .A1(G128), .A2(n916), .ZN(n809) );
  NAND2_X1 U892 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n811), .Z(n812) );
  NOR2_X1 U894 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n814), .ZN(n909) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n838) );
  NOR2_X1 U897 ( .A1(n909), .A2(n838), .ZN(n957) );
  NAND2_X1 U898 ( .A1(n848), .A2(n957), .ZN(n845) );
  NAND2_X1 U899 ( .A1(G131), .A2(n912), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G95), .A2(n599), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U902 ( .A(KEYINPUT93), .B(n817), .ZN(n821) );
  NAND2_X1 U903 ( .A1(n916), .A2(G119), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n915), .A2(G107), .ZN(n818) );
  AND2_X1 U905 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n821), .A2(n820), .ZN(n895) );
  NAND2_X1 U907 ( .A1(G1991), .A2(n895), .ZN(n822) );
  XOR2_X1 U908 ( .A(KEYINPUT94), .B(n822), .Z(n833) );
  NAND2_X1 U909 ( .A1(n915), .A2(G117), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G129), .A2(n916), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n824), .A2(n823), .ZN(n827) );
  NAND2_X1 U912 ( .A1(n599), .A2(G105), .ZN(n825) );
  XOR2_X1 U913 ( .A(KEYINPUT38), .B(n825), .Z(n826) );
  NOR2_X1 U914 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U915 ( .A(KEYINPUT95), .B(n828), .Z(n830) );
  NAND2_X1 U916 ( .A1(n912), .A2(G141), .ZN(n829) );
  NAND2_X1 U917 ( .A1(n830), .A2(n829), .ZN(n906) );
  NAND2_X1 U918 ( .A1(G1996), .A2(n906), .ZN(n831) );
  XOR2_X1 U919 ( .A(KEYINPUT96), .B(n831), .Z(n832) );
  NOR2_X1 U920 ( .A1(n833), .A2(n832), .ZN(n962) );
  INV_X1 U921 ( .A(n848), .ZN(n834) );
  NOR2_X1 U922 ( .A1(n962), .A2(n834), .ZN(n841) );
  INV_X1 U923 ( .A(n841), .ZN(n835) );
  XNOR2_X1 U924 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U925 ( .A1(n1005), .A2(n848), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(n851) );
  NAND2_X1 U927 ( .A1(n909), .A2(n838), .ZN(n950) );
  NOR2_X1 U928 ( .A1(G1996), .A2(n906), .ZN(n964) );
  NOR2_X1 U929 ( .A1(G1991), .A2(n895), .ZN(n953) );
  NOR2_X1 U930 ( .A1(G1986), .A2(G290), .ZN(n839) );
  NOR2_X1 U931 ( .A1(n953), .A2(n839), .ZN(n840) );
  NOR2_X1 U932 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U933 ( .A1(n964), .A2(n842), .ZN(n843) );
  XNOR2_X1 U934 ( .A(KEYINPUT39), .B(n843), .ZN(n844) );
  XNOR2_X1 U935 ( .A(n844), .B(KEYINPUT114), .ZN(n846) );
  NAND2_X1 U936 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U937 ( .A1(n950), .A2(n847), .ZN(n849) );
  NAND2_X1 U938 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U939 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U940 ( .A(n852), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U943 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U945 ( .A1(n856), .A2(n855), .ZN(G188) );
  XOR2_X1 U946 ( .A(G69), .B(KEYINPUT116), .Z(G235) );
  XNOR2_X1 U948 ( .A(KEYINPUT79), .B(n857), .ZN(n858) );
  NOR2_X1 U949 ( .A1(G860), .A2(n858), .ZN(n859) );
  XOR2_X1 U950 ( .A(n860), .B(n859), .Z(G145) );
  INV_X1 U951 ( .A(G132), .ZN(G219) );
  INV_X1 U952 ( .A(G108), .ZN(G238) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  INV_X1 U954 ( .A(G82), .ZN(G220) );
  INV_X1 U955 ( .A(G57), .ZN(G237) );
  NOR2_X1 U956 ( .A1(n862), .A2(n861), .ZN(G325) );
  INV_X1 U957 ( .A(G325), .ZN(G261) );
  INV_X1 U958 ( .A(n863), .ZN(G319) );
  XOR2_X1 U959 ( .A(G2096), .B(G2072), .Z(n865) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2090), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n875) );
  XOR2_X1 U962 ( .A(KEYINPUT120), .B(G2678), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U965 ( .A(G2100), .B(KEYINPUT43), .Z(n869) );
  XNOR2_X1 U966 ( .A(KEYINPUT42), .B(KEYINPUT119), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U969 ( .A(G2084), .B(G2078), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U971 ( .A(n875), .B(n874), .Z(G227) );
  XOR2_X1 U972 ( .A(G1956), .B(G1966), .Z(n877) );
  XNOR2_X1 U973 ( .A(G1986), .B(G1981), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n878), .B(KEYINPUT41), .Z(n880) );
  XNOR2_X1 U976 ( .A(G1996), .B(G1991), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U978 ( .A(G2474), .B(G1976), .Z(n882) );
  XNOR2_X1 U979 ( .A(G1961), .B(G1971), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(G229) );
  NAND2_X1 U982 ( .A1(G100), .A2(n599), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G112), .A2(n915), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(KEYINPUT121), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G136), .A2(n912), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n916), .A2(G124), .ZN(n890) );
  XOR2_X1 U989 ( .A(KEYINPUT44), .B(n890), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(G162) );
  XOR2_X1 U991 ( .A(KEYINPUT48), .B(KEYINPUT122), .Z(n894) );
  XNOR2_X1 U992 ( .A(G164), .B(KEYINPUT46), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n898) );
  XNOR2_X1 U994 ( .A(G162), .B(n895), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(n954), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n911) );
  NAND2_X1 U997 ( .A1(n915), .A2(G118), .ZN(n900) );
  NAND2_X1 U998 ( .A1(G130), .A2(n916), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n912), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n599), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(n903), .B(KEYINPUT45), .Z(n904) );
  NOR2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n923) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n912), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(G103), .A2(n599), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n921) );
  NAND2_X1 U1011 ( .A1(n915), .A2(G115), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(G127), .A2(n916), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1014 ( .A(KEYINPUT47), .B(n919), .Z(n920) );
  NOR2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n946) );
  XNOR2_X1 U1016 ( .A(n946), .B(G160), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n924), .ZN(G395) );
  XNOR2_X1 U1019 ( .A(n998), .B(n999), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n925), .B(G286), .ZN(n928) );
  XOR2_X1 U1021 ( .A(G301), .B(n926), .Z(n927) );
  XNOR2_X1 U1022 ( .A(n928), .B(n927), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n929), .ZN(G397) );
  XOR2_X1 U1024 ( .A(G2430), .B(G2451), .Z(n931) );
  XNOR2_X1 U1025 ( .A(G2446), .B(G2427), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n931), .B(n930), .ZN(n938) );
  XOR2_X1 U1027 ( .A(G2438), .B(G2435), .Z(n933) );
  XNOR2_X1 U1028 ( .A(G2443), .B(KEYINPUT115), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n933), .B(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(n934), .B(G2454), .Z(n936) );
  XNOR2_X1 U1031 ( .A(G1341), .B(G1348), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(G14), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(G319), .A2(n945), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(G227), .A2(G229), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT49), .B(n940), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(G395), .A2(G397), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(G225) );
  INV_X1 U1041 ( .A(G225), .ZN(G308) );
  INV_X1 U1042 ( .A(n945), .ZN(G401) );
  XOR2_X1 U1043 ( .A(G164), .B(G2078), .Z(n948) );
  XNOR2_X1 U1044 ( .A(n972), .B(n946), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n949), .B(KEYINPUT50), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n960) );
  XOR2_X1 U1048 ( .A(G160), .B(G2084), .Z(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT123), .B(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n967) );
  XOR2_X1 U1055 ( .A(G2090), .B(G162), .Z(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n965), .B(KEYINPUT51), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(KEYINPUT52), .B(n968), .ZN(n969) );
  INV_X1 U1060 ( .A(KEYINPUT55), .ZN(n991) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n991), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n970), .A2(G29), .ZN(n1047) );
  XOR2_X1 U1063 ( .A(KEYINPUT125), .B(KEYINPUT53), .Z(n984) );
  XOR2_X1 U1064 ( .A(n971), .B(G27), .Z(n974) );
  XNOR2_X1 U1065 ( .A(n972), .B(G33), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n978) );
  XOR2_X1 U1067 ( .A(G1991), .B(G25), .Z(n975) );
  NAND2_X1 U1068 ( .A1(n975), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT124), .B(n976), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(G2067), .B(G26), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G32), .B(G1996), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n984), .B(n983), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G2084), .B(G34), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n985), .B(KEYINPUT54), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(G35), .B(G2090), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n991), .B(n990), .ZN(n993) );
  INV_X1 U1082 ( .A(G29), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(G11), .A2(n994), .ZN(n1045) );
  XNOR2_X1 U1085 ( .A(G16), .B(KEYINPUT56), .ZN(n1018) );
  XOR2_X1 U1086 ( .A(G168), .B(G1966), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT57), .B(n997), .Z(n1016) );
  XNOR2_X1 U1089 ( .A(n998), .B(G1348), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G299), .B(G1956), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n999), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  NAND2_X1 U1095 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT126), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G301), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1043) );
  INV_X1 U1104 ( .A(G16), .ZN(n1041) );
  XOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .Z(n1019) );
  XNOR2_X1 U1106 ( .A(G4), .B(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(G20), .B(G1956), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(G1981), .B(G6), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(G19), .B(G1341), .ZN(n1022) );
  NOR2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(n1026), .B(KEYINPUT127), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(KEYINPUT60), .B(n1027), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(G1966), .B(G21), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G1961), .B(G5), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1038) );
  XNOR2_X1 U1119 ( .A(G1971), .B(G22), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(G23), .B(G1976), .ZN(n1032) );
  NOR2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1035) );
  XOR2_X1 U1122 ( .A(G1986), .B(G24), .Z(n1034) );
  NAND2_X1 U1123 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1124 ( .A(KEYINPUT58), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1125 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1126 ( .A(KEYINPUT61), .B(n1039), .ZN(n1040) );
  NAND2_X1 U1127 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1128 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NOR2_X1 U1129 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1130 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XOR2_X1 U1131 ( .A(KEYINPUT62), .B(n1048), .Z(G311) );
  INV_X1 U1132 ( .A(G311), .ZN(G150) );
endmodule

