//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G116), .B(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n194), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(KEYINPUT69), .A3(new_n204), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n210), .B(new_n211), .C1(new_n213), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(G146), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT0), .A4(G128), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT68), .B1(new_n216), .B2(new_n219), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT11), .B1(new_n223), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G134), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(new_n226), .B2(G134), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n223), .A3(G137), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n227), .ZN(new_n234));
  INV_X1    g048(.A(G131), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n229), .A4(new_n231), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n212), .C2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G128), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT66), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n217), .A3(new_n218), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n226), .A2(G134), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n223), .A2(G137), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n236), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n222), .A2(new_n237), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n209), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n216), .A2(new_n219), .ZN(new_n260));
  INV_X1    g074(.A(new_n236), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n229), .A2(new_n231), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n235), .B1(new_n262), .B2(new_n234), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n264), .A2(KEYINPUT65), .B1(new_n247), .B2(new_n251), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n216), .A2(new_n219), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n233), .B2(new_n236), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT30), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n219), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n237), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n251), .A2(new_n247), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(KEYINPUT30), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n205), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n253), .B(new_n259), .C1(new_n270), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n205), .B1(new_n252), .B2(KEYINPUT30), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n243), .A2(new_n246), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n236), .A2(new_n250), .ZN(new_n285));
  OAI22_X1  g099(.A1(new_n267), .A2(new_n268), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT65), .B(new_n266), .C1(new_n236), .C2(new_n233), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n253), .A4(new_n259), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n253), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n275), .A3(new_n269), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n277), .B1(new_n209), .B2(new_n252), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n295), .B2(new_n291), .ZN(new_n296));
  INV_X1    g110(.A(new_n259), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n281), .A2(new_n290), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n187), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n281), .A2(new_n290), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT32), .A3(new_n299), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n274), .A2(new_n275), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n207), .A2(new_n208), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n282), .B2(new_n288), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT71), .B1(new_n310), .B2(new_n259), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n253), .B1(new_n270), .B2(new_n278), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n297), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n259), .B(new_n292), .C1(new_n295), .C2(new_n291), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n311), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n309), .A2(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n307), .A2(new_n308), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n253), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(KEYINPUT28), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n297), .A2(new_n315), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n306), .B1(new_n324), .B2(G472), .ZN(new_n325));
  INV_X1    g139(.A(G472), .ZN(new_n326));
  AOI211_X1 g140(.A(KEYINPUT72), .B(new_n326), .C1(new_n317), .C2(new_n323), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n301), .B(new_n305), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G217), .ZN(new_n329));
  INV_X1    g143(.A(G902), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(G234), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT76), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G137), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT23), .B1(new_n244), .B2(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT73), .B1(new_n188), .B2(G128), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  XOR2_X1   g156(.A(G119), .B(G128), .Z(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n346));
  INV_X1    g160(.A(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G125), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G140), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT16), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT16), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n347), .A3(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G146), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n346), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n349), .A2(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n214), .B1(new_n356), .B2(new_n347), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT16), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(KEYINPUT74), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(G146), .B1(new_n358), .B2(new_n353), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n355), .A2(new_n359), .B1(new_n360), .B2(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n353), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n214), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n345), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n358), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n348), .A2(new_n350), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n341), .A2(new_n342), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n343), .A2(new_n344), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n338), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n343), .A2(new_n344), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n188), .B2(G128), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(new_n340), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n378), .B2(G110), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n214), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n351), .A2(new_n346), .A3(new_n354), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT74), .B1(new_n357), .B2(new_n358), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n373), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n337), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n374), .A2(new_n387), .A3(new_n330), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n374), .A2(new_n387), .A3(KEYINPUT25), .A4(new_n330), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n332), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n374), .A2(new_n387), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n331), .A2(G902), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G113), .B(G122), .ZN(new_n398));
  INV_X1    g212(.A(G104), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(G143), .B1(new_n255), .B2(G214), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n235), .ZN(new_n405));
  INV_X1    g219(.A(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n401), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G131), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n368), .B(KEYINPUT19), .Z(new_n410));
  OAI211_X1 g224(.A(new_n409), .B(new_n367), .C1(new_n410), .C2(G146), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n404), .B1(new_n412), .B2(new_n235), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n368), .B(new_n214), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(KEYINPUT18), .A3(G131), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n400), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n405), .A2(new_n408), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n355), .A2(new_n359), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n407), .A2(KEYINPUT17), .A3(G131), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n365), .A3(new_n380), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n423), .B2(KEYINPUT87), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n361), .A2(new_n425), .A3(new_n365), .A4(new_n422), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n418), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n417), .B1(new_n427), .B2(new_n400), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(KEYINPUT87), .ZN(new_n432));
  INV_X1    g246(.A(new_n420), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n400), .A3(new_n416), .ZN(new_n435));
  INV_X1    g249(.A(new_n417), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n429), .ZN(new_n439));
  INV_X1    g253(.A(new_n400), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n440), .B(new_n418), .C1(new_n424), .C2(new_n426), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n400), .B1(new_n434), .B2(new_n416), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n330), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n431), .A2(new_n439), .B1(new_n443), .B2(G475), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT9), .B(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n445), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n233), .A2(new_n449), .A3(new_n236), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n233), .B2(new_n236), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n399), .A2(G107), .ZN(new_n453));
  INV_X1    g267(.A(G101), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n456));
  INV_X1    g270(.A(G107), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G104), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT3), .A4(G104), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n399), .A2(G107), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n454), .B1(new_n464), .B2(new_n453), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT10), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n455), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT3), .B1(new_n463), .B2(new_n456), .ZN(new_n469));
  INV_X1    g283(.A(new_n461), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n244), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n246), .B1(new_n472), .B2(new_n238), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n457), .A2(G104), .ZN(new_n474));
  OAI21_X1  g288(.A(G101), .B1(new_n463), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n247), .A2(new_n467), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n460), .B2(new_n461), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n471), .B(KEYINPUT4), .C1(new_n478), .C2(new_n454), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n460), .A2(new_n461), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n453), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n454), .A2(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n479), .A2(new_n271), .A3(new_n273), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n452), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n462), .A2(new_n465), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n476), .B1(new_n247), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n237), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G140), .ZN(new_n491));
  INV_X1    g305(.A(G227), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n487), .A2(new_n237), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n485), .A2(new_n490), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n483), .A2(new_n273), .A3(new_n271), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n471), .A2(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n454), .B1(new_n480), .B2(new_n453), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n467), .A2(new_n247), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n476), .A2(new_n466), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n237), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n495), .B1(new_n507), .B2(new_n485), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n498), .B1(new_n508), .B2(KEYINPUT80), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n510));
  AOI211_X1 g324(.A(new_n510), .B(new_n495), .C1(new_n507), .C2(new_n485), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n448), .B(new_n330), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n471), .A2(new_n475), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n246), .A3(new_n243), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n514), .A2(new_n476), .B1(new_n236), .B2(new_n233), .ZN(new_n515));
  INV_X1    g329(.A(new_n489), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n497), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n452), .A2(new_n477), .A3(new_n484), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n494), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n507), .A2(new_n495), .A3(new_n485), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(G469), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(G469), .A2(G902), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n447), .B1(new_n512), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n525));
  INV_X1    g339(.A(G122), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G116), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n190), .A2(G122), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n457), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n212), .A2(G128), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n244), .A2(G143), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n223), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G134), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT88), .B1(new_n528), .B2(KEYINPUT14), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT14), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n190), .A4(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(KEYINPUT14), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n538), .A2(new_n527), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G107), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n527), .A2(new_n528), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G107), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n547), .A2(new_n529), .B1(new_n533), .B2(new_n223), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n531), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n532), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n531), .A2(new_n549), .ZN(new_n552));
  OAI21_X1  g366(.A(G134), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n445), .A2(new_n329), .A3(G953), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n545), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n545), .B2(new_n554), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n525), .B(new_n330), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(G478), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n545), .A2(new_n554), .ZN(new_n561));
  INV_X1    g375(.A(new_n555), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n537), .A2(new_n544), .B1(new_n548), .B2(new_n553), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n555), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(G478), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n525), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT90), .B(G952), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G953), .ZN(new_n571));
  NAND2_X1  g385(.A1(G234), .A2(G237), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT21), .B(G898), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(G902), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n574), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G214), .B1(G237), .B2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n582));
  OAI21_X1  g396(.A(G113), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n201), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n486), .ZN(new_n586));
  INV_X1    g400(.A(new_n482), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n203), .B(new_n204), .C1(new_n478), .C2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n502), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(G110), .B(G122), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n586), .B(new_n590), .C1(new_n502), .C2(new_n588), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(KEYINPUT6), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT6), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n589), .A2(new_n595), .A3(new_n591), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n243), .A2(new_n349), .A3(new_n246), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n266), .A2(G125), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n333), .A2(G224), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT81), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n599), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n594), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n583), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n200), .A2(KEYINPUT5), .ZN(new_n606));
  OAI211_X1 g420(.A(KEYINPUT82), .B(G113), .C1(new_n189), .C2(KEYINPUT5), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n513), .B1(new_n201), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n590), .B(KEYINPUT8), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n486), .B2(new_n584), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT83), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n201), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n486), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n585), .A2(new_n513), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .A4(new_n610), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n597), .A2(KEYINPUT84), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n598), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n597), .A2(KEYINPUT84), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT85), .B(KEYINPUT7), .ZN(new_n622));
  OAI22_X1  g436(.A1(new_n620), .A2(new_n621), .B1(new_n601), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT7), .B1(new_n601), .B2(KEYINPUT86), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(KEYINPUT86), .B2(new_n601), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n598), .A3(new_n597), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n618), .A2(new_n593), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n603), .A2(new_n330), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G210), .B1(G237), .B2(G902), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n603), .A2(new_n330), .A3(new_n627), .A4(new_n629), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n581), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n444), .A2(new_n524), .A3(new_n579), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n328), .A2(new_n397), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  INV_X1    g450(.A(new_n524), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n304), .A2(new_n299), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n397), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n438), .B1(new_n437), .B2(new_n429), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT20), .B(new_n430), .C1(new_n435), .C2(new_n436), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n434), .A2(new_n416), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n440), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n646), .B2(new_n435), .ZN(new_n647));
  INV_X1    g461(.A(G475), .ZN(new_n648));
  OAI22_X1  g462(.A1(new_n643), .A2(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR3_X1    g463(.A1(new_n566), .A2(KEYINPUT93), .A3(G478), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT93), .B1(new_n566), .B2(G478), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n563), .A2(new_n565), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT33), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n562), .B1(new_n564), .B2(KEYINPUT91), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n545), .A2(KEYINPUT91), .A3(new_n554), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT92), .ZN(new_n657));
  OAI22_X1  g471(.A1(new_n655), .A2(new_n656), .B1(new_n556), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT91), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n555), .B1(new_n561), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n564), .A2(KEYINPUT91), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(KEYINPUT92), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n654), .B1(new_n663), .B2(KEYINPUT33), .ZN(new_n664));
  INV_X1    g478(.A(G478), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(G902), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n652), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n578), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n627), .A2(new_n330), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n629), .B1(new_n671), .B2(new_n603), .ZN(new_n672));
  INV_X1    g486(.A(new_n632), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n670), .B(new_n580), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n642), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  INV_X1    g492(.A(KEYINPUT94), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n439), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n437), .A2(KEYINPUT94), .A3(new_n438), .A4(new_n429), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n431), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n560), .A2(new_n568), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(G475), .B2(new_n443), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n674), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n642), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  INV_X1    g503(.A(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n390), .A2(new_n391), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n331), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n361), .A2(new_n365), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n373), .B1(new_n693), .B2(new_n379), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n338), .A2(KEYINPUT36), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n394), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n692), .A2(KEYINPUT95), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT95), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n392), .B2(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n690), .B1(new_n640), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT95), .B1(new_n692), .B2(new_n699), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n392), .A2(new_n698), .A3(new_n701), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(KEYINPUT96), .A3(new_n639), .A4(new_n638), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n634), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT37), .B(G110), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G12));
  NAND2_X1  g525(.A1(new_n512), .A2(new_n523), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n446), .A3(new_n702), .A4(new_n700), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n574), .B1(new_n715), .B2(new_n577), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n682), .A2(new_n684), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n631), .A2(new_n632), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n580), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n328), .A2(new_n714), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G128), .ZN(G30));
  XNOR2_X1  g537(.A(new_n719), .B(KEYINPUT38), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n259), .B1(new_n253), .B2(new_n319), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n726), .A2(new_n279), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n728), .B2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n301), .A3(new_n305), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n692), .A2(new_n699), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n444), .A2(new_n731), .A3(new_n683), .A4(new_n581), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n724), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT98), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n716), .B(KEYINPUT39), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n637), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(KEYINPUT40), .Z(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n212), .ZN(G45));
  INV_X1    g553(.A(KEYINPUT99), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n649), .A2(new_n668), .A3(new_n717), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(new_n720), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n660), .A2(new_n661), .B1(KEYINPUT92), .B2(new_n565), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT33), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n654), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n747), .A2(new_n666), .B1(new_n651), .B2(new_n650), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n444), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT99), .A3(new_n633), .A4(new_n717), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n328), .A2(new_n714), .A3(new_n742), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  OAI21_X1  g566(.A(new_n330), .B1(new_n509), .B2(new_n511), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n512), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n755), .A2(new_n641), .A3(new_n447), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n328), .A2(new_n675), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NOR2_X1   g573(.A1(new_n325), .A2(new_n327), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n305), .A2(new_n301), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n686), .B(new_n756), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G116), .ZN(G18));
  NAND4_X1  g577(.A1(new_n633), .A2(new_n446), .A3(new_n512), .A4(new_n754), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n444), .A2(new_n700), .A3(new_n579), .A4(new_n702), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n328), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  INV_X1    g582(.A(new_n764), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n302), .B1(new_n259), .B2(new_n321), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n299), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n638), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT100), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n397), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n649), .A2(new_n569), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n578), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n769), .A2(new_n773), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  NAND3_X1  g595(.A1(new_n771), .A2(new_n638), .A3(new_n731), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n741), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n769), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT101), .B(G125), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G27));
  INV_X1    g600(.A(new_n777), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n305), .A2(KEYINPUT104), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT104), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n304), .A2(new_n789), .A3(KEYINPUT32), .A4(new_n299), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n788), .A2(new_n790), .A3(new_n301), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n292), .A3(new_n322), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n330), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n310), .A2(KEYINPUT71), .A3(new_n259), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n313), .B1(new_n312), .B2(new_n297), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n316), .A2(new_n315), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT72), .B1(new_n799), .B2(new_n326), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n324), .A2(new_n306), .A3(G472), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n787), .B1(new_n791), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n631), .A2(new_n446), .A3(new_n580), .A4(new_n632), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n520), .A2(KEYINPUT103), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT103), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n507), .A2(new_n807), .A3(new_n485), .A4(new_n495), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(G469), .A3(new_n519), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n522), .B(KEYINPUT102), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n512), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT42), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n813), .A3(new_n741), .ZN(new_n814));
  INV_X1    g628(.A(new_n741), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n512), .A2(new_n809), .A3(new_n810), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n641), .A3(new_n804), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n815), .B(new_n817), .C1(new_n760), .C2(new_n761), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n803), .A2(new_n814), .B1(new_n818), .B2(new_n813), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n235), .ZN(G33));
  INV_X1    g634(.A(new_n718), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n328), .A2(new_n821), .A3(new_n817), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G134), .ZN(G36));
  NAND2_X1  g637(.A1(new_n444), .A2(new_n668), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT43), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n640), .A3(new_n731), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT44), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n631), .A2(new_n580), .A3(new_n632), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n735), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n806), .A2(KEYINPUT45), .A3(new_n519), .A4(new_n808), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n519), .A2(new_n520), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n833), .B(G469), .C1(KEYINPUT45), .C2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n810), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT46), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n512), .B1(new_n836), .B2(KEYINPUT46), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n446), .B(new_n832), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n828), .B2(new_n827), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n831), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(KEYINPUT105), .B(G137), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(G39));
  OAI21_X1  g657(.A(new_n446), .B1(new_n837), .B2(new_n838), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT47), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n328), .A2(new_n397), .A3(new_n741), .A4(new_n830), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT106), .B(G140), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(G42));
  NAND3_X1  g664(.A1(new_n788), .A2(new_n790), .A3(new_n301), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n777), .B1(new_n851), .B2(new_n760), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n755), .A2(new_n573), .A3(new_n804), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n826), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT48), .Z(new_n856));
  INV_X1    g670(.A(new_n730), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n853), .A3(new_n397), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n749), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n787), .A2(new_n772), .A3(new_n573), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n826), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n769), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n571), .A3(new_n860), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n444), .A3(new_n748), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n782), .B2(new_n854), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n724), .A2(new_n580), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n862), .A2(new_n868), .A3(new_n447), .A4(new_n755), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT50), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n830), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n755), .A2(new_n446), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n873), .B(new_n863), .C1(new_n846), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n865), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n778), .A2(new_n720), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n731), .A2(new_n447), .A3(new_n716), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n730), .A3(new_n811), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n751), .A2(new_n722), .A3(new_n784), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n784), .A2(new_n883), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n751), .A3(KEYINPUT52), .A4(new_n722), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n783), .A2(new_n811), .A3(new_n805), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n822), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n761), .B1(new_n800), .B2(new_n801), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n683), .B(new_n717), .C1(new_n647), .C2(new_n648), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n830), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n707), .A3(new_n524), .A4(new_n682), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n672), .A2(new_n673), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n716), .B(new_n569), .C1(new_n443), .C2(G475), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n682), .A3(new_n900), .A4(new_n580), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n713), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n328), .A2(new_n902), .A3(KEYINPUT110), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n892), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n803), .A2(new_n814), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n818), .A2(new_n813), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n757), .A2(new_n762), .A3(new_n780), .A4(new_n767), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT108), .B1(new_n444), .B2(new_n748), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n578), .B(new_n581), .C1(new_n631), .C2(new_n632), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT108), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n649), .A2(new_n911), .A3(new_n668), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT109), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n431), .A2(new_n439), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n684), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n684), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT109), .B1(new_n674), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n913), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n642), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n921), .A2(new_n635), .A3(new_n709), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n904), .A2(new_n907), .A3(new_n908), .A4(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n880), .B1(new_n890), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(new_n722), .A3(new_n751), .A4(new_n784), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n886), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n894), .A2(new_n893), .A3(new_n897), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT110), .B1(new_n328), .B2(new_n902), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n822), .B(new_n891), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n921), .A2(new_n635), .A3(new_n709), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT113), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n757), .A2(new_n762), .A3(new_n780), .A4(new_n767), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n819), .A2(new_n933), .A3(new_n880), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT113), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n898), .A2(new_n903), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n812), .A2(new_n782), .A3(new_n741), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n805), .A2(new_n397), .A3(new_n811), .ZN(new_n938));
  INV_X1    g752(.A(new_n761), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n802), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n940), .B2(new_n821), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n922), .A2(new_n935), .A3(new_n936), .A4(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n927), .A2(new_n932), .A3(new_n934), .A4(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n924), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n751), .A2(new_n722), .A3(new_n784), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n947), .A2(new_n925), .B1(new_n884), .B2(new_n885), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n880), .B1(new_n923), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT111), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(KEYINPUT111), .B(new_n880), .C1(new_n923), .C2(new_n948), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n930), .A2(new_n931), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n819), .A2(new_n933), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n889), .A2(new_n953), .A3(KEYINPUT53), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT112), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n907), .A2(new_n908), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n635), .A2(new_n709), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(new_n936), .A3(new_n941), .A4(new_n921), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT112), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT53), .A4(new_n889), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n951), .A2(new_n952), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT54), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n945), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI22_X1  g779(.A1(new_n879), .A2(new_n965), .B1(G952), .B2(G953), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n755), .A2(KEYINPUT49), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT107), .Z(new_n968));
  NOR3_X1   g782(.A1(new_n724), .A2(new_n447), .A3(new_n581), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n824), .B1(new_n755), .B2(KEYINPUT49), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n969), .A2(new_n857), .A3(new_n777), .A4(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n966), .B1(new_n968), .B2(new_n971), .ZN(G75));
  NOR2_X1   g786(.A1(new_n333), .A2(G952), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n330), .B1(new_n924), .B2(new_n943), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT56), .B1(new_n974), .B2(G210), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n594), .A2(new_n596), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n602), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT55), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT115), .ZN(new_n981));
  OR3_X1    g795(.A1(new_n975), .A2(new_n981), .A3(new_n979), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n975), .B2(new_n979), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n973), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(G51));
  INV_X1    g798(.A(new_n944), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT53), .B1(new_n960), .B2(new_n889), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n927), .A2(new_n932), .A3(new_n934), .A4(new_n942), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT116), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n989), .A3(new_n945), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n924), .A2(new_n943), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(KEYINPUT116), .A3(new_n985), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n810), .B(KEYINPUT57), .Z(new_n993));
  NAND3_X1  g807(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n511), .B2(new_n509), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n835), .B(KEYINPUT117), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n974), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n973), .B1(new_n995), .B2(new_n997), .ZN(G54));
  NAND3_X1  g812(.A1(new_n974), .A2(KEYINPUT58), .A3(G475), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n999), .A2(new_n428), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n428), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n973), .ZN(G60));
  INV_X1    g816(.A(new_n945), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n956), .A2(new_n962), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n960), .A2(new_n927), .ZN(new_n1005));
  AOI21_X1  g819(.A(KEYINPUT111), .B1(new_n1005), .B2(new_n880), .ZN(new_n1006));
  INV_X1    g820(.A(new_n952), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1003), .B1(new_n1008), .B2(KEYINPUT54), .ZN(new_n1009));
  XNOR2_X1  g823(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n665), .A2(new_n330), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1010), .B(new_n1011), .Z(new_n1012));
  OAI21_X1  g826(.A(new_n664), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT119), .ZN(new_n1014));
  INV_X1    g828(.A(new_n973), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n664), .A2(new_n1012), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n990), .A2(new_n992), .A3(new_n1016), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1012), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n747), .B1(new_n965), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1017), .A2(new_n1015), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT119), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1018), .A2(new_n1022), .ZN(G63));
  INV_X1    g837(.A(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G217), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT120), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT60), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n991), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1028), .A2(new_n393), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1024), .B1(new_n1029), .B2(KEYINPUT122), .ZN(new_n1030));
  INV_X1    g844(.A(new_n696), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n991), .A2(new_n1031), .A3(new_n1027), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT122), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n1028), .B2(new_n393), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1030), .A2(new_n1015), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1032), .A2(new_n1015), .ZN(new_n1036));
  OAI211_X1 g850(.A(KEYINPUT121), .B(new_n1024), .C1(new_n1029), .C2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1024), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT121), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1035), .A2(new_n1037), .A3(new_n1040), .ZN(G66));
  INV_X1    g855(.A(G224), .ZN(new_n1042));
  OAI21_X1  g856(.A(G953), .B1(new_n575), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n933), .A2(new_n931), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1043), .B1(new_n1044), .B2(G953), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n976), .B1(G898), .B2(new_n333), .ZN(new_n1046));
  XNOR2_X1  g860(.A(new_n1045), .B(new_n1046), .ZN(G69));
  AOI22_X1  g861(.A1(new_n846), .A2(new_n847), .B1(new_n831), .B2(new_n840), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n819), .B1(new_n821), .B2(new_n940), .ZN(new_n1049));
  NOR4_X1   g863(.A1(new_n839), .A2(new_n852), .A3(new_n720), .A4(new_n778), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1050), .A2(new_n946), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n1048), .A2(new_n333), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1052), .B1(new_n715), .B2(new_n333), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n288), .A2(new_n276), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1054), .B(new_n410), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  OR3_X1    g870(.A1(new_n738), .A2(KEYINPUT62), .A3(new_n946), .ZN(new_n1057));
  OAI21_X1  g871(.A(KEYINPUT62), .B1(new_n738), .B2(new_n946), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n328), .A2(new_n397), .A3(new_n736), .A4(new_n873), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n916), .B1(new_n909), .B2(new_n912), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g875(.A(new_n1061), .B(KEYINPUT123), .Z(new_n1062));
  NAND4_X1  g876(.A1(new_n1057), .A2(new_n1048), .A3(new_n1058), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n1055), .A2(G953), .ZN(new_n1064));
  OAI21_X1  g878(.A(G953), .B1(new_n492), .B2(new_n715), .ZN(new_n1065));
  AOI22_X1  g879(.A1(new_n1063), .A2(new_n1064), .B1(KEYINPUT124), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1056), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n1065), .A2(KEYINPUT124), .ZN(new_n1068));
  XNOR2_X1  g882(.A(new_n1068), .B(KEYINPUT125), .ZN(new_n1069));
  XOR2_X1   g883(.A(new_n1067), .B(new_n1069), .Z(G72));
  NAND2_X1  g884(.A1(new_n310), .A2(new_n297), .ZN(new_n1071));
  NAND4_X1  g885(.A1(new_n1048), .A2(new_n1044), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1072));
  NAND2_X1  g886(.A1(G472), .A2(G902), .ZN(new_n1073));
  XOR2_X1   g887(.A(new_n1073), .B(KEYINPUT63), .Z(new_n1074));
  AOI21_X1  g888(.A(new_n1071), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g889(.A(KEYINPUT126), .ZN(new_n1076));
  OR3_X1    g890(.A1(new_n1075), .A2(new_n1076), .A3(new_n973), .ZN(new_n1077));
  OAI21_X1  g891(.A(new_n1076), .B1(new_n1075), .B2(new_n973), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g893(.A1(new_n797), .A2(new_n279), .ZN(new_n1080));
  NAND3_X1  g894(.A1(new_n1008), .A2(new_n1074), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g895(.A(new_n1044), .ZN(new_n1082));
  OAI21_X1  g896(.A(new_n1074), .B1(new_n1063), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g897(.A1(new_n1083), .A2(new_n312), .A3(new_n259), .ZN(new_n1084));
  NAND3_X1  g898(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1085), .A2(KEYINPUT127), .ZN(new_n1086));
  INV_X1    g900(.A(KEYINPUT127), .ZN(new_n1087));
  NAND4_X1  g901(.A1(new_n1079), .A2(new_n1087), .A3(new_n1081), .A4(new_n1084), .ZN(new_n1088));
  NAND2_X1  g902(.A1(new_n1086), .A2(new_n1088), .ZN(G57));
endmodule


