

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n725), .A2(n724), .ZN(n772) );
  XOR2_X1 U555 ( .A(KEYINPUT14), .B(n574), .Z(n521) );
  XNOR2_X2 U556 ( .A(n784), .B(KEYINPUT32), .ZN(n803) );
  NOR2_X1 U557 ( .A1(n772), .A2(n961), .ZN(n727) );
  NAND2_X1 U558 ( .A1(n890), .A2(G138), .ZN(n535) );
  AND2_X1 U559 ( .A1(n893), .A2(G114), .ZN(n522) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n726) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n749) );
  INV_X1 U562 ( .A(KEYINPUT109), .ZN(n799) );
  INV_X1 U563 ( .A(KEYINPUT17), .ZN(n529) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n541), .Z(n658) );
  OR2_X1 U565 ( .A1(n538), .A2(n522), .ZN(n539) );
  XOR2_X1 U566 ( .A(KEYINPUT23), .B(KEYINPUT68), .Z(n524) );
  XOR2_X1 U567 ( .A(KEYINPUT66), .B(G2104), .Z(n525) );
  NOR2_X1 U568 ( .A1(n525), .A2(G2105), .ZN(n611) );
  NAND2_X1 U569 ( .A1(G101), .A2(n611), .ZN(n523) );
  XNOR2_X1 U570 ( .A(n524), .B(n523), .ZN(n528) );
  AND2_X2 U571 ( .A1(n525), .A2(G2105), .ZN(n894) );
  NAND2_X1 U572 ( .A1(G125), .A2(n894), .ZN(n526) );
  XOR2_X1 U573 ( .A(KEYINPUT67), .B(n526), .Z(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n534) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XNOR2_X2 U576 ( .A(n530), .B(n529), .ZN(n890) );
  NAND2_X1 U577 ( .A1(G137), .A2(n890), .ZN(n532) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U579 ( .A1(G113), .A2(n893), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U581 ( .A1(n534), .A2(n533), .ZN(G160) );
  XNOR2_X1 U582 ( .A(KEYINPUT97), .B(n535), .ZN(n540) );
  NAND2_X1 U583 ( .A1(G102), .A2(n611), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G126), .A2(n894), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U586 ( .A1(n540), .A2(n539), .ZN(G164) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n654) );
  NOR2_X1 U588 ( .A1(G651), .A2(n654), .ZN(n653) );
  NAND2_X1 U589 ( .A1(G52), .A2(n653), .ZN(n543) );
  INV_X1 U590 ( .A(G651), .ZN(n545) );
  NOR2_X1 U591 ( .A1(G543), .A2(n545), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G64), .A2(n658), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U594 ( .A(KEYINPUT71), .B(n544), .Z(n550) );
  NOR2_X1 U595 ( .A1(n654), .A2(n545), .ZN(n646) );
  NAND2_X1 U596 ( .A1(G77), .A2(n646), .ZN(n547) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n643) );
  NAND2_X1 U598 ( .A1(G90), .A2(n643), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U601 ( .A1(n550), .A2(n549), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  XOR2_X1 U605 ( .A(KEYINPUT4), .B(KEYINPUT80), .Z(n552) );
  NAND2_X1 U606 ( .A1(G89), .A2(n643), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U608 ( .A(KEYINPUT79), .B(n553), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n646), .A2(G76), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n556), .ZN(n562) );
  NAND2_X1 U612 ( .A1(n658), .A2(G63), .ZN(n557) );
  XOR2_X1 U613 ( .A(KEYINPUT81), .B(n557), .Z(n559) );
  NAND2_X1 U614 ( .A1(n653), .A2(G51), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(n563), .ZN(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(n564) );
  XNOR2_X1 U620 ( .A(KEYINPUT82), .B(n564), .ZN(G286) );
  XOR2_X1 U621 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n566) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U623 ( .A(n566), .B(n565), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n838) );
  NAND2_X1 U625 ( .A1(n838), .A2(G567), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  XOR2_X1 U627 ( .A(G860), .B(KEYINPUT77), .Z(n601) );
  NAND2_X1 U628 ( .A1(n643), .A2(G81), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G68), .A2(n646), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT13), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G43), .A2(n653), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n658), .A2(G56), .ZN(n574) );
  NOR2_X1 U636 ( .A1(n575), .A2(n521), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT76), .B(n576), .Z(n983) );
  INV_X1 U638 ( .A(n983), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n601), .A2(n577), .ZN(G153) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G79), .A2(n646), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G92), .A2(n643), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G54), .A2(n653), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G66), .A2(n658), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT15), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(KEYINPUT78), .B(n585), .ZN(n737) );
  INV_X1 U650 ( .A(n737), .ZN(n984) );
  NOR2_X1 U651 ( .A1(n984), .A2(G868), .ZN(n587) );
  INV_X1 U652 ( .A(G868), .ZN(n672) );
  NOR2_X1 U653 ( .A1(n672), .A2(G301), .ZN(n586) );
  NOR2_X1 U654 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G91), .A2(n643), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT72), .B(n588), .Z(n593) );
  NAND2_X1 U657 ( .A1(G53), .A2(n653), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G65), .A2(n658), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U660 ( .A(KEYINPUT73), .B(n591), .Z(n592) );
  NOR2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n646), .A2(G78), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G299) );
  XNOR2_X1 U664 ( .A(KEYINPUT83), .B(G868), .ZN(n596) );
  NOR2_X1 U665 ( .A1(G286), .A2(n596), .ZN(n599) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT84), .ZN(n598) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(G297) );
  INV_X1 U669 ( .A(G559), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U671 ( .A1(n984), .A2(n602), .ZN(n603) );
  XOR2_X1 U672 ( .A(KEYINPUT16), .B(n603), .Z(G148) );
  NOR2_X1 U673 ( .A1(n983), .A2(G868), .ZN(n604) );
  XOR2_X1 U674 ( .A(KEYINPUT85), .B(n604), .Z(n607) );
  NAND2_X1 U675 ( .A1(G868), .A2(n737), .ZN(n605) );
  NOR2_X1 U676 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G135), .A2(n890), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G111), .A2(n893), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G123), .A2(n894), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT18), .ZN(n613) );
  BUF_X1 U683 ( .A(n611), .Z(n878) );
  NAND2_X1 U684 ( .A1(n878), .A2(G99), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n942) );
  XOR2_X1 U687 ( .A(G2096), .B(n942), .Z(n616) );
  NOR2_X1 U688 ( .A1(G2100), .A2(n616), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT86), .B(n617), .Z(G156) );
  NAND2_X1 U690 ( .A1(G80), .A2(n646), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G93), .A2(n643), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U693 ( .A(KEYINPUT88), .B(n620), .Z(n622) );
  NAND2_X1 U694 ( .A1(n653), .A2(G55), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G67), .A2(n658), .ZN(n623) );
  XNOR2_X1 U697 ( .A(KEYINPUT89), .B(n623), .ZN(n624) );
  OR2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n671) );
  NAND2_X1 U699 ( .A1(n737), .A2(G559), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(n983), .ZN(n668) );
  NOR2_X1 U701 ( .A1(n668), .A2(G860), .ZN(n627) );
  XOR2_X1 U702 ( .A(KEYINPUT87), .B(n627), .Z(n628) );
  XOR2_X1 U703 ( .A(n671), .B(n628), .Z(G145) );
  NAND2_X1 U704 ( .A1(n653), .A2(G47), .ZN(n635) );
  NAND2_X1 U705 ( .A1(G72), .A2(n646), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G85), .A2(n643), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G60), .A2(n658), .ZN(n631) );
  XNOR2_X1 U709 ( .A(KEYINPUT69), .B(n631), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT70), .ZN(G290) );
  NAND2_X1 U713 ( .A1(G75), .A2(n646), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G88), .A2(n643), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G50), .A2(n653), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G62), .A2(n658), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(G166) );
  NAND2_X1 U720 ( .A1(G86), .A2(n643), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G48), .A2(n653), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G73), .A2(n646), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n647), .B(KEYINPUT91), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(KEYINPUT2), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n658), .A2(G61), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n660) );
  NAND2_X1 U730 ( .A1(G49), .A2(n653), .ZN(n656) );
  NAND2_X1 U731 ( .A1(G87), .A2(n654), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(KEYINPUT90), .ZN(G288) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(KEYINPUT92), .Z(n663) );
  INV_X1 U737 ( .A(G299), .ZN(n990) );
  XNOR2_X1 U738 ( .A(n990), .B(G166), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U740 ( .A(n671), .B(n664), .Z(n666) );
  XNOR2_X1 U741 ( .A(G305), .B(G288), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U743 ( .A(G290), .B(n667), .ZN(n905) );
  XNOR2_X1 U744 ( .A(n668), .B(n905), .ZN(n669) );
  XNOR2_X1 U745 ( .A(KEYINPUT93), .B(n669), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U748 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(KEYINPUT94), .Z(n675) );
  XNOR2_X1 U751 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U754 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XOR2_X1 U755 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n681) );
  XNOR2_X1 U758 ( .A(KEYINPUT22), .B(KEYINPUT95), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U760 ( .A1(n682), .A2(G218), .ZN(n683) );
  NAND2_X1 U761 ( .A1(G96), .A2(n683), .ZN(n844) );
  NAND2_X1 U762 ( .A1(n844), .A2(G2106), .ZN(n688) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U765 ( .A1(G108), .A2(n685), .ZN(n843) );
  NAND2_X1 U766 ( .A1(G567), .A2(n843), .ZN(n686) );
  XNOR2_X1 U767 ( .A(KEYINPUT96), .B(n686), .ZN(n687) );
  NAND2_X1 U768 ( .A1(n688), .A2(n687), .ZN(n845) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U770 ( .A1(n845), .A2(n689), .ZN(n842) );
  NAND2_X1 U771 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G166), .ZN(G303) );
  NAND2_X1 U773 ( .A1(G119), .A2(n894), .ZN(n696) );
  NAND2_X1 U774 ( .A1(G131), .A2(n890), .ZN(n691) );
  NAND2_X1 U775 ( .A1(G95), .A2(n878), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U777 ( .A1(G107), .A2(n893), .ZN(n692) );
  XNOR2_X1 U778 ( .A(KEYINPUT101), .B(n692), .ZN(n693) );
  NOR2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U780 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U781 ( .A(n697), .B(KEYINPUT102), .ZN(n872) );
  AND2_X1 U782 ( .A1(G1991), .A2(n872), .ZN(n706) );
  NAND2_X1 U783 ( .A1(G141), .A2(n890), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G117), .A2(n893), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U786 ( .A1(n878), .A2(G105), .ZN(n700) );
  XOR2_X1 U787 ( .A(KEYINPUT38), .B(n700), .Z(n701) );
  NOR2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n894), .A2(G129), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n704), .A2(n703), .ZN(n873) );
  AND2_X1 U791 ( .A1(G1996), .A2(n873), .ZN(n705) );
  NOR2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n932) );
  NOR2_X1 U793 ( .A1(G164), .A2(G1384), .ZN(n708) );
  INV_X1 U794 ( .A(KEYINPUT65), .ZN(n707) );
  XNOR2_X1 U795 ( .A(n708), .B(n707), .ZN(n724) );
  NAND2_X1 U796 ( .A1(G160), .A2(G40), .ZN(n723) );
  NOR2_X1 U797 ( .A1(n724), .A2(n723), .ZN(n709) );
  XNOR2_X1 U798 ( .A(KEYINPUT98), .B(n709), .ZN(n831) );
  XNOR2_X1 U799 ( .A(KEYINPUT103), .B(n831), .ZN(n710) );
  NOR2_X1 U800 ( .A1(n932), .A2(n710), .ZN(n823) );
  XOR2_X1 U801 ( .A(KEYINPUT104), .B(n823), .Z(n722) );
  XNOR2_X1 U802 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n715) );
  NAND2_X1 U803 ( .A1(G116), .A2(n893), .ZN(n712) );
  NAND2_X1 U804 ( .A1(G128), .A2(n894), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT35), .ZN(n714) );
  XNOR2_X1 U807 ( .A(n715), .B(n714), .ZN(n720) );
  NAND2_X1 U808 ( .A1(G140), .A2(n890), .ZN(n717) );
  NAND2_X1 U809 ( .A1(G104), .A2(n878), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U811 ( .A(KEYINPUT34), .B(n718), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U813 ( .A(KEYINPUT36), .B(n721), .ZN(n902) );
  XNOR2_X1 U814 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NOR2_X1 U815 ( .A1(n902), .A2(n828), .ZN(n938) );
  NAND2_X1 U816 ( .A1(n938), .A2(n831), .ZN(n826) );
  NAND2_X1 U817 ( .A1(n722), .A2(n826), .ZN(n818) );
  XNOR2_X1 U818 ( .A(KEYINPUT105), .B(n723), .ZN(n725) );
  INV_X1 U819 ( .A(G1996), .ZN(n961) );
  XNOR2_X1 U820 ( .A(n727), .B(n726), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n772), .A2(G1341), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n983), .A2(n730), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n736), .A2(n737), .ZN(n734) );
  INV_X1 U825 ( .A(n772), .ZN(n752) );
  NOR2_X1 U826 ( .A1(n752), .A2(G1348), .ZN(n732) );
  NOR2_X1 U827 ( .A1(G2067), .A2(n772), .ZN(n731) );
  NOR2_X1 U828 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U830 ( .A(n735), .B(KEYINPUT108), .ZN(n739) );
  OR2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n752), .A2(G2072), .ZN(n740) );
  XNOR2_X1 U834 ( .A(n740), .B(KEYINPUT27), .ZN(n742) );
  INV_X1 U835 ( .A(G1956), .ZN(n1006) );
  NOR2_X1 U836 ( .A1(n1006), .A2(n752), .ZN(n741) );
  NOR2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n745) );
  NAND2_X1 U838 ( .A1(n990), .A2(n745), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n748) );
  NOR2_X1 U840 ( .A1(n990), .A2(n745), .ZN(n746) );
  XOR2_X1 U841 ( .A(n746), .B(KEYINPUT28), .Z(n747) );
  NAND2_X1 U842 ( .A1(n748), .A2(n747), .ZN(n750) );
  XNOR2_X1 U843 ( .A(n750), .B(n749), .ZN(n770) );
  NOR2_X1 U844 ( .A1(n752), .A2(G1961), .ZN(n751) );
  XNOR2_X1 U845 ( .A(KEYINPUT107), .B(n751), .ZN(n754) );
  XNOR2_X1 U846 ( .A(KEYINPUT25), .B(G2078), .ZN(n967) );
  NAND2_X1 U847 ( .A1(n967), .A2(n752), .ZN(n753) );
  NAND2_X1 U848 ( .A1(n754), .A2(n753), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n763), .A2(G171), .ZN(n771) );
  NOR2_X1 U850 ( .A1(G2084), .A2(n772), .ZN(n758) );
  AND2_X1 U851 ( .A1(G8), .A2(n758), .ZN(n755) );
  NAND2_X1 U852 ( .A1(G8), .A2(n772), .ZN(n814) );
  NOR2_X1 U853 ( .A1(G1966), .A2(n814), .ZN(n759) );
  OR2_X1 U854 ( .A1(n755), .A2(n759), .ZN(n767) );
  INV_X1 U855 ( .A(n767), .ZN(n756) );
  AND2_X1 U856 ( .A1(n771), .A2(n756), .ZN(n757) );
  NAND2_X1 U857 ( .A1(n770), .A2(n757), .ZN(n769) );
  NOR2_X1 U858 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U859 ( .A1(G8), .A2(n760), .ZN(n761) );
  XNOR2_X1 U860 ( .A(KEYINPUT30), .B(n761), .ZN(n762) );
  NOR2_X1 U861 ( .A1(G168), .A2(n762), .ZN(n765) );
  NOR2_X1 U862 ( .A1(G171), .A2(n763), .ZN(n764) );
  NOR2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U864 ( .A(KEYINPUT31), .B(n766), .Z(n776) );
  OR2_X1 U865 ( .A1(n767), .A2(n776), .ZN(n768) );
  AND2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n804) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n989) );
  AND2_X1 U868 ( .A1(n804), .A2(n989), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n771), .A2(n770), .ZN(n778) );
  NOR2_X1 U870 ( .A1(G1971), .A2(n814), .ZN(n774) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n772), .ZN(n773) );
  NOR2_X1 U872 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U873 ( .A1(n775), .A2(G303), .ZN(n779) );
  AND2_X1 U874 ( .A1(n776), .A2(n779), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n783) );
  INV_X1 U876 ( .A(n779), .ZN(n780) );
  OR2_X1 U877 ( .A1(n780), .A2(G286), .ZN(n781) );
  AND2_X1 U878 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n803), .ZN(n790) );
  INV_X1 U881 ( .A(n989), .ZN(n787) );
  NOR2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n795) );
  NOR2_X1 U883 ( .A1(G1971), .A2(G303), .ZN(n786) );
  NOR2_X1 U884 ( .A1(n795), .A2(n786), .ZN(n991) );
  OR2_X1 U885 ( .A1(n787), .A2(n991), .ZN(n788) );
  OR2_X1 U886 ( .A1(n814), .A2(n788), .ZN(n789) );
  NAND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U888 ( .A(n791), .B(KEYINPUT64), .ZN(n793) );
  INV_X1 U889 ( .A(KEYINPUT33), .ZN(n792) );
  NAND2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n798) );
  INV_X1 U891 ( .A(n814), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n796), .A2(KEYINPUT33), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n800) );
  XNOR2_X1 U895 ( .A(n800), .B(n799), .ZN(n802) );
  XOR2_X1 U896 ( .A(G1981), .B(KEYINPUT110), .Z(n801) );
  XNOR2_X1 U897 ( .A(G305), .B(n801), .ZN(n980) );
  NAND2_X1 U898 ( .A1(n802), .A2(n980), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n807) );
  NOR2_X1 U900 ( .A1(G2090), .A2(G303), .ZN(n805) );
  NAND2_X1 U901 ( .A1(G8), .A2(n805), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n808), .A2(n814), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n816) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XOR2_X1 U906 ( .A(n811), .B(KEYINPUT106), .Z(n812) );
  XNOR2_X1 U907 ( .A(KEYINPUT24), .B(n812), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n820) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U912 ( .A1(n998), .A2(n831), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n834) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n873), .ZN(n935) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n872), .ZN(n941) );
  NOR2_X1 U917 ( .A1(n821), .A2(n941), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n935), .A2(n824), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n902), .A2(n828), .ZN(n940) );
  NAND2_X1 U923 ( .A1(n829), .A2(n940), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT111), .B(n830), .Z(n832) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n837) );
  XOR2_X1 U927 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n835) );
  XNOR2_X1 U928 ( .A(KEYINPUT40), .B(n835), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n837), .B(n836), .ZN(G329) );
  NAND2_X1 U930 ( .A1(n838), .A2(G2106), .ZN(n839) );
  XOR2_X1 U931 ( .A(KEYINPUT117), .B(n839), .Z(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U933 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  INV_X1 U942 ( .A(n845), .ZN(G319) );
  XOR2_X1 U943 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U952 ( .A(G1976), .B(G1971), .Z(n855) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1961), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n856), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(G2474), .B(G1981), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1966), .B(G1956), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G124), .A2(n894), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n863), .B(KEYINPUT118), .ZN(n864) );
  XNOR2_X1 U964 ( .A(KEYINPUT44), .B(n864), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G112), .A2(n893), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT119), .B(n865), .Z(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G136), .A2(n890), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G100), .A2(n878), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U972 ( .A(n942), .B(G162), .Z(n875) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n889) );
  NAND2_X1 U975 ( .A1(G118), .A2(n893), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G130), .A2(n894), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G142), .A2(n890), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G106), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(n884), .Z(n885) );
  XOR2_X1 U984 ( .A(n885), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U985 ( .A(G164), .B(KEYINPUT120), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(n889), .B(n888), .Z(n901) );
  NAND2_X1 U988 ( .A1(G139), .A2(n890), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G103), .A2(n878), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U991 ( .A1(G115), .A2(n893), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G127), .A2(n894), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n928) );
  XNOR2_X1 U996 ( .A(G160), .B(n928), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U998 ( .A(n903), .B(n902), .Z(n904) );
  NOR2_X1 U999 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(n983), .B(G286), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1002 ( .A(n984), .B(G171), .Z(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1005 ( .A(G2438), .B(G2435), .Z(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT116), .B(G2454), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1008 ( .A(G2427), .B(G2443), .Z(n913) );
  XNOR2_X1 U1009 ( .A(KEYINPUT115), .B(G2446), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT114), .B(G2451), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n920) );
  XOR2_X1 U1014 ( .A(G1341), .B(G1348), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G2430), .B(n918), .ZN(n919) );
  XOR2_X1 U1016 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1017 ( .A1(G14), .A2(n921), .ZN(n927) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n927), .ZN(G401) );
  XOR2_X1 U1027 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n931), .Z(n952) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n949) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT122), .B(n937), .ZN(n947) );
  INV_X1 U1037 ( .A(n938), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n943), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT123), .B(n950), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n953), .ZN(n954) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n976), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(G29), .ZN(n1034) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(G34), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT125), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G2084), .B(n957), .ZN(n974) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n972) );
  XNOR2_X1 U1054 ( .A(G1991), .B(G25), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G2067), .B(G26), .Z(n960) );
  NAND2_X1 U1058 ( .A1(n960), .A2(G28), .ZN(n964) );
  XOR2_X1 U1059 ( .A(G32), .B(n961), .Z(n962) );
  XNOR2_X1 U1060 ( .A(KEYINPUT124), .B(n962), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1063 ( .A(G27), .B(n967), .Z(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n970), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1069 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n979), .ZN(n1032) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT57), .ZN(n1003) );
  XNOR2_X1 U1076 ( .A(n983), .B(G1341), .ZN(n1001) );
  XNOR2_X1 U1077 ( .A(G301), .B(G1961), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n984), .B(G1348), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT126), .B(n987), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n990), .B(G1956), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(KEYINPUT127), .B(n999), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1030) );
  INV_X1 U1092 ( .A(G16), .ZN(n1028) );
  XNOR2_X1 U1093 ( .A(G20), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G6), .B(G1981), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1014), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1025) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

