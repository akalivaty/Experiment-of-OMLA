

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747;

  OR2_X1 U366 ( .A1(n511), .A2(n465), .ZN(n466) );
  XNOR2_X1 U367 ( .A(n575), .B(n574), .ZN(n584) );
  BUF_X1 U368 ( .A(n544), .Z(n346) );
  NOR2_X1 U369 ( .A1(n567), .A2(n494), .ZN(n430) );
  XNOR2_X1 U370 ( .A(n526), .B(KEYINPUT1), .ZN(n544) );
  AND2_X1 U371 ( .A1(n365), .A2(n364), .ZN(n363) );
  BUF_X1 U372 ( .A(G953), .Z(n345) );
  XNOR2_X1 U373 ( .A(n398), .B(n397), .ZN(n635) );
  XNOR2_X1 U374 ( .A(n456), .B(n396), .ZN(n397) );
  XNOR2_X1 U375 ( .A(n393), .B(n392), .ZN(n723) );
  XNOR2_X1 U376 ( .A(n348), .B(n386), .ZN(n407) );
  XNOR2_X1 U377 ( .A(n483), .B(n357), .ZN(n738) );
  XNOR2_X1 U378 ( .A(n448), .B(n391), .ZN(n483) );
  XNOR2_X1 U379 ( .A(n347), .B(G104), .ZN(n393) );
  XNOR2_X1 U380 ( .A(n400), .B(KEYINPUT15), .ZN(n605) );
  INV_X2 U381 ( .A(G107), .ZN(n347) );
  XNOR2_X1 U382 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n449) );
  NAND2_X2 U383 ( .A1(n379), .A2(n378), .ZN(n747) );
  NAND2_X1 U384 ( .A1(n493), .A2(n681), .ZN(n686) );
  XNOR2_X2 U385 ( .A(n424), .B(n423), .ZN(n493) );
  INV_X1 U386 ( .A(n453), .ZN(n451) );
  XNOR2_X1 U387 ( .A(n446), .B(n447), .ZN(n453) );
  INV_X1 U388 ( .A(G902), .ZN(n478) );
  XNOR2_X2 U389 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n444) );
  XNOR2_X2 U390 ( .A(n723), .B(n434), .ZN(n456) );
  XNOR2_X2 U391 ( .A(n522), .B(KEYINPUT19), .ZN(n555) );
  XNOR2_X1 U392 ( .A(n566), .B(KEYINPUT31), .ZN(n389) );
  NOR2_X1 U393 ( .A1(n565), .A2(n703), .ZN(n559) );
  XNOR2_X2 U394 ( .A(G146), .B(G125), .ZN(n406) );
  INV_X1 U395 ( .A(KEYINPUT75), .ZN(n351) );
  XNOR2_X2 U396 ( .A(G146), .B(G125), .ZN(n348) );
  AND2_X2 U397 ( .A1(n610), .A2(n676), .ZN(n639) );
  OR2_X1 U398 ( .A1(n565), .A2(n691), .ZN(n566) );
  NAND2_X1 U399 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U400 ( .A(n549), .B(n548), .ZN(n703) );
  XNOR2_X1 U401 ( .A(n563), .B(KEYINPUT109), .ZN(n546) );
  NAND2_X1 U402 ( .A1(n516), .A2(n695), .ZN(n506) );
  OR2_X1 U403 ( .A1(n616), .A2(G902), .ZN(n441) );
  XNOR2_X1 U404 ( .A(n449), .B(n358), .ZN(n357) );
  XNOR2_X1 U405 ( .A(G137), .B(G131), .ZN(n358) );
  XNOR2_X2 U406 ( .A(n595), .B(n594), .ZN(n625) );
  INV_X1 U407 ( .A(n398), .ZN(n349) );
  INV_X1 U408 ( .A(n362), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n738), .B(G146), .ZN(n431) );
  XNOR2_X1 U410 ( .A(n674), .B(n351), .ZN(n352) );
  OR2_X1 U411 ( .A1(n526), .A2(n686), .ZN(n567) );
  XOR2_X2 U412 ( .A(n417), .B(n416), .Z(n611) );
  INV_X1 U413 ( .A(KEYINPUT18), .ZN(n385) );
  AND2_X1 U414 ( .A1(G469), .A2(n478), .ZN(n361) );
  INV_X1 U415 ( .A(G237), .ZN(n442) );
  XNOR2_X1 U416 ( .A(G119), .B(G128), .ZN(n410) );
  INV_X1 U417 ( .A(G140), .ZN(n386) );
  INV_X1 U418 ( .A(KEYINPUT84), .ZN(n601) );
  XNOR2_X1 U419 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U420 ( .A(n372), .B(KEYINPUT76), .ZN(n471) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n372) );
  XNOR2_X1 U422 ( .A(n505), .B(n504), .ZN(n532) );
  INV_X1 U423 ( .A(KEYINPUT46), .ZN(n504) );
  NOR2_X1 U424 ( .A1(n747), .A2(n746), .ZN(n505) );
  XNOR2_X1 U425 ( .A(n420), .B(n419), .ZN(n422) );
  NAND2_X2 U426 ( .A1(n363), .A2(n360), .ZN(n526) );
  NAND2_X1 U427 ( .A1(n362), .A2(n361), .ZN(n360) );
  NAND2_X1 U428 ( .A1(G902), .A2(n399), .ZN(n364) );
  XNOR2_X1 U429 ( .A(G116), .B(G107), .ZN(n481) );
  INV_X1 U430 ( .A(KEYINPUT40), .ZN(n384) );
  NAND2_X1 U431 ( .A1(n661), .A2(n384), .ZN(n382) );
  XNOR2_X1 U432 ( .A(n443), .B(KEYINPUT30), .ZN(n377) );
  INV_X1 U433 ( .A(KEYINPUT0), .ZN(n556) );
  XNOR2_X1 U434 ( .A(n616), .B(KEYINPUT62), .ZN(n617) );
  INV_X2 U435 ( .A(G953), .ZN(n739) );
  NAND2_X1 U436 ( .A1(n356), .A2(n354), .ZN(n610) );
  XNOR2_X1 U437 ( .A(n628), .B(KEYINPUT59), .ZN(n629) );
  XNOR2_X1 U438 ( .A(n641), .B(n643), .ZN(n644) );
  NAND2_X1 U439 ( .A1(n380), .A2(n381), .ZN(n378) );
  AND2_X1 U440 ( .A1(n383), .A2(n382), .ZN(n379) );
  NOR2_X1 U441 ( .A1(n661), .A2(n384), .ZN(n381) );
  BUF_X1 U442 ( .A(n389), .Z(n355) );
  NOR2_X1 U443 ( .A1(n511), .A2(n377), .ZN(n353) );
  OR2_X1 U444 ( .A1(n605), .A2(n604), .ZN(n354) );
  NAND2_X1 U445 ( .A1(n603), .A2(n352), .ZN(n356) );
  XNOR2_X2 U446 ( .A(G143), .B(G128), .ZN(n448) );
  INV_X1 U447 ( .A(n635), .ZN(n362) );
  NAND2_X1 U448 ( .A1(n635), .A2(n399), .ZN(n365) );
  XNOR2_X1 U449 ( .A(n366), .B(KEYINPUT45), .ZN(n607) );
  NAND2_X1 U450 ( .A1(n368), .A2(n367), .ZN(n366) );
  XNOR2_X1 U451 ( .A(n369), .B(KEYINPUT87), .ZN(n367) );
  NAND2_X1 U452 ( .A1(n371), .A2(n370), .ZN(n368) );
  NAND2_X1 U453 ( .A1(n581), .A2(n582), .ZN(n369) );
  NAND2_X1 U454 ( .A1(n599), .A2(KEYINPUT44), .ZN(n370) );
  NAND2_X1 U455 ( .A1(n598), .A2(n597), .ZN(n371) );
  XNOR2_X1 U456 ( .A(n406), .B(n385), .ZN(n447) );
  XNOR2_X1 U457 ( .A(n349), .B(n373), .ZN(n616) );
  XNOR2_X1 U458 ( .A(n375), .B(n374), .ZN(n373) );
  XNOR2_X1 U459 ( .A(n432), .B(n433), .ZN(n374) );
  XNOR2_X1 U460 ( .A(n460), .B(n436), .ZN(n375) );
  NAND2_X1 U461 ( .A1(n376), .A2(n696), .ZN(n465) );
  INV_X1 U462 ( .A(n377), .ZN(n376) );
  INV_X1 U463 ( .A(n534), .ZN(n380) );
  XNOR2_X2 U464 ( .A(n466), .B(n467), .ZN(n534) );
  NAND2_X1 U465 ( .A1(n534), .A2(n384), .ZN(n383) );
  NAND2_X1 U466 ( .A1(n388), .A2(n387), .ZN(n570) );
  INV_X1 U467 ( .A(n650), .ZN(n387) );
  INV_X1 U468 ( .A(n389), .ZN(n388) );
  NAND2_X1 U469 ( .A1(n355), .A2(n666), .ZN(n667) );
  NAND2_X1 U470 ( .A1(n355), .A2(n668), .ZN(n669) );
  BUF_X1 U471 ( .A(n639), .Z(n718) );
  NOR2_X1 U472 ( .A1(n704), .A2(n703), .ZN(n390) );
  INV_X1 U473 ( .A(n627), .ZN(n596) );
  INV_X1 U474 ( .A(KEYINPUT68), .ZN(n529) );
  XNOR2_X1 U475 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U476 ( .A1(n555), .A2(n508), .ZN(n662) );
  INV_X1 U477 ( .A(KEYINPUT63), .ZN(n620) );
  INV_X1 U478 ( .A(KEYINPUT39), .ZN(n467) );
  INV_X1 U479 ( .A(G134), .ZN(n391) );
  INV_X1 U480 ( .A(n431), .ZN(n398) );
  XNOR2_X1 U481 ( .A(G110), .B(KEYINPUT91), .ZN(n392) );
  XNOR2_X1 U482 ( .A(KEYINPUT66), .B(G101), .ZN(n434) );
  XNOR2_X1 U483 ( .A(KEYINPUT95), .B(G140), .ZN(n395) );
  NAND2_X1 U484 ( .A1(n739), .A2(G227), .ZN(n394) );
  XNOR2_X1 U485 ( .A(n395), .B(n394), .ZN(n396) );
  INV_X1 U486 ( .A(G469), .ZN(n399) );
  XNOR2_X1 U487 ( .A(G902), .B(KEYINPUT90), .ZN(n400) );
  NAND2_X1 U488 ( .A1(n605), .A2(G234), .ZN(n401) );
  XNOR2_X1 U489 ( .A(n401), .B(KEYINPUT20), .ZN(n418) );
  AND2_X1 U490 ( .A1(n418), .A2(G221), .ZN(n403) );
  XNOR2_X1 U491 ( .A(KEYINPUT100), .B(KEYINPUT21), .ZN(n402) );
  XNOR2_X1 U492 ( .A(n403), .B(n402), .ZN(n681) );
  NAND2_X1 U493 ( .A1(n739), .A2(G234), .ZN(n405) );
  XNOR2_X1 U494 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n404) );
  XNOR2_X1 U495 ( .A(n405), .B(n404), .ZN(n485) );
  NAND2_X1 U496 ( .A1(n485), .A2(G221), .ZN(n409) );
  XOR2_X1 U497 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n408) );
  XNOR2_X2 U498 ( .A(n408), .B(n407), .ZN(n737) );
  XNOR2_X1 U499 ( .A(n409), .B(n737), .ZN(n417) );
  XOR2_X1 U500 ( .A(G110), .B(G137), .Z(n411) );
  XNOR2_X1 U501 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U502 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n413) );
  XNOR2_X1 U503 ( .A(KEYINPUT96), .B(KEYINPUT24), .ZN(n412) );
  XNOR2_X1 U504 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U505 ( .A(n415), .B(n414), .Z(n416) );
  NOR2_X1 U506 ( .A1(n611), .A2(G902), .ZN(n424) );
  NAND2_X1 U507 ( .A1(n418), .A2(G217), .ZN(n420) );
  XNOR2_X1 U508 ( .A(KEYINPUT98), .B(KEYINPUT25), .ZN(n419) );
  XOR2_X1 U509 ( .A(KEYINPUT99), .B(KEYINPUT78), .Z(n421) );
  XOR2_X1 U510 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n426) );
  NAND2_X1 U511 ( .A1(G237), .A2(G234), .ZN(n425) );
  XNOR2_X1 U512 ( .A(n426), .B(n425), .ZN(n427) );
  NAND2_X1 U513 ( .A1(G952), .A2(n427), .ZN(n708) );
  NOR2_X1 U514 ( .A1(n345), .A2(n708), .ZN(n552) );
  NAND2_X1 U515 ( .A1(G902), .A2(n427), .ZN(n550) );
  OR2_X1 U516 ( .A1(n739), .A2(n550), .ZN(n428) );
  NOR2_X1 U517 ( .A1(G900), .A2(n428), .ZN(n429) );
  NOR2_X1 U518 ( .A1(n552), .A2(n429), .ZN(n494) );
  XNOR2_X1 U519 ( .A(n430), .B(KEYINPUT77), .ZN(n511) );
  XOR2_X1 U520 ( .A(KEYINPUT5), .B(KEYINPUT101), .Z(n433) );
  NAND2_X1 U521 ( .A1(n471), .A2(G210), .ZN(n432) );
  XNOR2_X1 U522 ( .A(KEYINPUT74), .B(KEYINPUT102), .ZN(n435) );
  XNOR2_X1 U523 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U524 ( .A(G119), .B(G116), .ZN(n438) );
  XNOR2_X1 U525 ( .A(G113), .B(KEYINPUT69), .ZN(n437) );
  XNOR2_X1 U526 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U527 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n439) );
  XNOR2_X1 U528 ( .A(n440), .B(n439), .ZN(n460) );
  XNOR2_X2 U529 ( .A(n441), .B(G472), .ZN(n585) );
  NAND2_X1 U530 ( .A1(n478), .A2(n442), .ZN(n462) );
  NAND2_X1 U531 ( .A1(n462), .A2(G214), .ZN(n695) );
  NAND2_X1 U532 ( .A1(n585), .A2(n695), .ZN(n443) );
  NAND2_X1 U533 ( .A1(G224), .A2(n739), .ZN(n445) );
  XNOR2_X1 U534 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U535 ( .A(n449), .B(n448), .ZN(n452) );
  INV_X1 U536 ( .A(n452), .ZN(n450) );
  NAND2_X1 U537 ( .A1(n451), .A2(n450), .ZN(n455) );
  NAND2_X1 U538 ( .A1(n453), .A2(n452), .ZN(n454) );
  NAND2_X1 U539 ( .A1(n455), .A2(n454), .ZN(n457) );
  XNOR2_X1 U540 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U541 ( .A(KEYINPUT16), .B(G122), .ZN(n458) );
  XNOR2_X1 U542 ( .A(n458), .B(KEYINPUT72), .ZN(n459) );
  XNOR2_X1 U543 ( .A(n460), .B(n459), .ZN(n725) );
  XNOR2_X1 U544 ( .A(n461), .B(n725), .ZN(n640) );
  NAND2_X1 U545 ( .A1(n640), .A2(n605), .ZN(n464) );
  AND2_X1 U546 ( .A1(n462), .A2(G210), .ZN(n463) );
  XNOR2_X2 U547 ( .A(n464), .B(n463), .ZN(n516) );
  INV_X1 U548 ( .A(n516), .ZN(n540) );
  XNOR2_X1 U549 ( .A(n540), .B(KEYINPUT38), .ZN(n696) );
  XOR2_X1 U550 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n469) );
  XNOR2_X1 U551 ( .A(G122), .B(KEYINPUT103), .ZN(n468) );
  XNOR2_X1 U552 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U553 ( .A(n737), .B(n470), .Z(n477) );
  AND2_X1 U554 ( .A1(n471), .A2(G214), .ZN(n473) );
  XNOR2_X1 U555 ( .A(G143), .B(G131), .ZN(n472) );
  XNOR2_X1 U556 ( .A(n473), .B(n472), .ZN(n475) );
  XOR2_X1 U557 ( .A(G104), .B(G113), .Z(n474) );
  XNOR2_X1 U558 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U559 ( .A(n477), .B(n476), .ZN(n628) );
  NAND2_X1 U560 ( .A1(n628), .A2(n478), .ZN(n480) );
  XOR2_X1 U561 ( .A(KEYINPUT13), .B(G475), .Z(n479) );
  XNOR2_X1 U562 ( .A(n480), .B(n479), .ZN(n513) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(G122), .Z(n482) );
  XNOR2_X1 U564 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U565 ( .A(n484), .B(n483), .ZN(n491) );
  NAND2_X1 U566 ( .A1(G217), .A2(n485), .ZN(n489) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n487) );
  XNOR2_X1 U568 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n486) );
  XNOR2_X1 U569 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U570 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U571 ( .A(n491), .B(n490), .ZN(n719) );
  NOR2_X1 U572 ( .A1(G902), .A2(n719), .ZN(n492) );
  XNOR2_X1 U573 ( .A(G478), .B(n492), .ZN(n509) );
  AND2_X1 U574 ( .A1(n513), .A2(n509), .ZN(n666) );
  INV_X1 U575 ( .A(n666), .ZN(n661) );
  NOR2_X1 U576 ( .A1(n494), .A2(n493), .ZN(n495) );
  NAND2_X1 U577 ( .A1(n495), .A2(n681), .ZN(n519) );
  INV_X1 U578 ( .A(n519), .ZN(n496) );
  NAND2_X1 U579 ( .A1(n585), .A2(n496), .ZN(n498) );
  INV_X1 U580 ( .A(KEYINPUT28), .ZN(n497) );
  XNOR2_X1 U581 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U582 ( .A(n526), .B(KEYINPUT113), .ZN(n499) );
  NAND2_X1 U583 ( .A1(n500), .A2(n499), .ZN(n507) );
  INV_X1 U584 ( .A(n509), .ZN(n512) );
  OR2_X1 U585 ( .A1(n513), .A2(n512), .ZN(n698) );
  NAND2_X1 U586 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U587 ( .A1(n698), .A2(n699), .ZN(n502) );
  XNOR2_X1 U588 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n501) );
  XNOR2_X1 U589 ( .A(n502), .B(n501), .ZN(n710) );
  NOR2_X1 U590 ( .A1(n507), .A2(n710), .ZN(n503) );
  XNOR2_X1 U591 ( .A(n503), .B(KEYINPUT42), .ZN(n746) );
  XNOR2_X2 U592 ( .A(n506), .B(KEYINPUT88), .ZN(n522) );
  INV_X1 U593 ( .A(n507), .ZN(n508) );
  OR2_X1 U594 ( .A1(n513), .A2(n509), .ZN(n657) );
  INV_X1 U595 ( .A(n657), .ZN(n668) );
  XNOR2_X1 U596 ( .A(KEYINPUT107), .B(n668), .ZN(n535) );
  AND2_X1 U597 ( .A1(n535), .A2(n661), .ZN(n700) );
  NOR2_X1 U598 ( .A1(n662), .A2(n700), .ZN(n510) );
  XNOR2_X1 U599 ( .A(n510), .B(KEYINPUT47), .ZN(n518) );
  NAND2_X1 U600 ( .A1(n513), .A2(n512), .ZN(n515) );
  INV_X1 U601 ( .A(KEYINPUT110), .ZN(n514) );
  XNOR2_X1 U602 ( .A(n515), .B(n514), .ZN(n560) );
  AND2_X1 U603 ( .A1(n516), .A2(n560), .ZN(n517) );
  NAND2_X1 U604 ( .A1(n353), .A2(n517), .ZN(n660) );
  AND2_X1 U605 ( .A1(n518), .A2(n660), .ZN(n528) );
  XNOR2_X1 U606 ( .A(n585), .B(KEYINPUT6), .ZN(n589) );
  OR2_X1 U607 ( .A1(n589), .A2(n519), .ZN(n520) );
  XNOR2_X1 U608 ( .A(n520), .B(KEYINPUT111), .ZN(n521) );
  AND2_X1 U609 ( .A1(n521), .A2(n666), .ZN(n537) );
  INV_X1 U610 ( .A(n522), .ZN(n523) );
  NAND2_X1 U611 ( .A1(n537), .A2(n523), .ZN(n525) );
  INV_X1 U612 ( .A(KEYINPUT36), .ZN(n524) );
  XNOR2_X1 U613 ( .A(n525), .B(n524), .ZN(n527) );
  INV_X1 U614 ( .A(n346), .ZN(n590) );
  NAND2_X1 U615 ( .A1(n527), .A2(n590), .ZN(n670) );
  AND2_X1 U616 ( .A1(n528), .A2(n670), .ZN(n530) );
  NOR2_X2 U617 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U618 ( .A(n533), .B(KEYINPUT48), .ZN(n543) );
  NOR2_X1 U619 ( .A1(n535), .A2(n534), .ZN(n672) );
  AND2_X1 U620 ( .A1(n346), .A2(n695), .ZN(n536) );
  NAND2_X1 U621 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U622 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n538) );
  XNOR2_X1 U623 ( .A(n539), .B(n538), .ZN(n541) );
  AND2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n624) );
  NOR2_X1 U625 ( .A1(n672), .A2(n624), .ZN(n542) );
  AND2_X2 U626 ( .A1(n543), .A2(n542), .ZN(n674) );
  OR2_X2 U627 ( .A1(n544), .A2(n686), .ZN(n563) );
  INV_X1 U628 ( .A(n589), .ZN(n545) );
  NAND2_X1 U629 ( .A1(n546), .A2(n545), .ZN(n549) );
  INV_X1 U630 ( .A(KEYINPUT70), .ZN(n547) );
  XNOR2_X1 U631 ( .A(n547), .B(KEYINPUT33), .ZN(n548) );
  XNOR2_X1 U632 ( .A(G898), .B(KEYINPUT93), .ZN(n732) );
  NAND2_X1 U633 ( .A1(n345), .A2(n732), .ZN(n726) );
  NOR2_X1 U634 ( .A1(n550), .A2(n726), .ZN(n551) );
  OR2_X1 U635 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U636 ( .A(n553), .B(KEYINPUT94), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X2 U638 ( .A(n557), .B(n556), .ZN(n573) );
  INV_X1 U639 ( .A(n573), .ZN(n565) );
  XOR2_X1 U640 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n558) );
  XNOR2_X1 U641 ( .A(n559), .B(n558), .ZN(n561) );
  NAND2_X1 U642 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X2 U643 ( .A(n562), .B(KEYINPUT35), .ZN(n627) );
  NAND2_X1 U644 ( .A1(n627), .A2(KEYINPUT44), .ZN(n582) );
  INV_X1 U645 ( .A(n563), .ZN(n564) );
  NAND2_X1 U646 ( .A1(n564), .A2(n585), .ZN(n691) );
  NOR2_X1 U647 ( .A1(n567), .A2(n585), .ZN(n568) );
  AND2_X1 U648 ( .A1(n573), .A2(n568), .ZN(n650) );
  INV_X1 U649 ( .A(n700), .ZN(n569) );
  NAND2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n580) );
  INV_X1 U651 ( .A(n698), .ZN(n571) );
  AND2_X1 U652 ( .A1(n571), .A2(n681), .ZN(n572) );
  XNOR2_X1 U653 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n574) );
  BUF_X1 U654 ( .A(n584), .Z(n576) );
  INV_X1 U655 ( .A(n576), .ZN(n579) );
  AND2_X1 U656 ( .A1(n589), .A2(n493), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n577), .A2(n346), .ZN(n578) );
  OR2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n623) );
  AND2_X1 U659 ( .A1(n580), .A2(n623), .ZN(n581) );
  INV_X1 U660 ( .A(n493), .ZN(n583) );
  AND2_X2 U661 ( .A1(n584), .A2(n583), .ZN(n593) );
  INV_X1 U662 ( .A(n585), .ZN(n684) );
  AND2_X1 U663 ( .A1(n346), .A2(n684), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n593), .A2(n586), .ZN(n588) );
  INV_X1 U665 ( .A(KEYINPUT108), .ZN(n587) );
  XNOR2_X1 U666 ( .A(n588), .B(n587), .ZN(n626) );
  XNOR2_X1 U667 ( .A(n589), .B(KEYINPUT80), .ZN(n591) );
  AND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n595) );
  INV_X1 U670 ( .A(KEYINPUT32), .ZN(n594) );
  NOR2_X2 U671 ( .A1(n626), .A2(n625), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n599), .A2(n596), .ZN(n598) );
  INV_X1 U673 ( .A(KEYINPUT44), .ZN(n597) );
  INV_X1 U674 ( .A(n605), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n607), .A2(n600), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(n601), .ZN(n603) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n674), .A2(KEYINPUT2), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT85), .ZN(n609) );
  BUF_X1 U680 ( .A(n607), .Z(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n676) );
  NAND2_X1 U682 ( .A1(n639), .A2(G217), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U684 ( .A(G952), .ZN(n613) );
  AND2_X1 U685 ( .A1(n613), .A2(n345), .ZN(n722) );
  NOR2_X2 U686 ( .A1(n614), .A2(n722), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n615), .B(KEYINPUT126), .ZN(G66) );
  NAND2_X1 U688 ( .A1(n639), .A2(G472), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X2 U690 ( .A1(n619), .A2(n722), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G57) );
  XOR2_X1 U692 ( .A(G101), .B(KEYINPUT115), .Z(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(G3) );
  XOR2_X1 U694 ( .A(G140), .B(n624), .Z(G42) );
  XOR2_X1 U695 ( .A(n625), .B(G119), .Z(G21) );
  XOR2_X1 U696 ( .A(G110), .B(n626), .Z(G12) );
  XOR2_X1 U697 ( .A(n627), .B(G122), .Z(G24) );
  NAND2_X1 U698 ( .A1(n639), .A2(G475), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U700 ( .A1(n631), .A2(n722), .ZN(n633) );
  XOR2_X1 U701 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n632) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(G60) );
  NAND2_X1 U703 ( .A1(n718), .A2(G469), .ZN(n637) );
  XOR2_X1 U704 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n634) );
  XNOR2_X1 U705 ( .A(n350), .B(n634), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U707 ( .A1(n638), .A2(n722), .ZN(G54) );
  NAND2_X1 U708 ( .A1(n639), .A2(G210), .ZN(n645) );
  BUF_X1 U709 ( .A(n640), .Z(n641) );
  XNOR2_X1 U710 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n642) );
  XOR2_X1 U711 ( .A(n642), .B(KEYINPUT55), .Z(n643) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X2 U713 ( .A1(n646), .A2(n722), .ZN(n648) );
  XNOR2_X1 U714 ( .A(KEYINPUT86), .B(KEYINPUT56), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(G51) );
  NAND2_X1 U716 ( .A1(n650), .A2(n666), .ZN(n649) );
  XNOR2_X1 U717 ( .A(n649), .B(G104), .ZN(G6) );
  NAND2_X1 U718 ( .A1(n650), .A2(n668), .ZN(n656) );
  XOR2_X1 U719 ( .A(KEYINPUT118), .B(KEYINPUT27), .Z(n652) );
  XNOR2_X1 U720 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n654) );
  XOR2_X1 U722 ( .A(G107), .B(KEYINPUT26), .Z(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(G9) );
  NOR2_X1 U725 ( .A1(n662), .A2(n657), .ZN(n659) );
  XNOR2_X1 U726 ( .A(G128), .B(KEYINPUT29), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(G30) );
  XNOR2_X1 U728 ( .A(G143), .B(n660), .ZN(G45) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n664) );
  XNOR2_X1 U730 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U732 ( .A(G146), .B(n665), .ZN(G48) );
  XNOR2_X1 U733 ( .A(n667), .B(G113), .ZN(G15) );
  XNOR2_X1 U734 ( .A(n669), .B(G116), .ZN(G18) );
  XOR2_X1 U735 ( .A(G125), .B(n670), .Z(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U737 ( .A(G134), .B(n672), .Z(G36) );
  NOR2_X1 U738 ( .A1(n608), .A2(KEYINPUT2), .ZN(n673) );
  XOR2_X1 U739 ( .A(KEYINPUT82), .B(n673), .Z(n680) );
  NOR2_X1 U740 ( .A1(n674), .A2(KEYINPUT2), .ZN(n675) );
  XOR2_X1 U741 ( .A(KEYINPUT83), .B(n675), .Z(n678) );
  INV_X1 U742 ( .A(n676), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n715) );
  NOR2_X1 U745 ( .A1(n681), .A2(n493), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT121), .B(n682), .Z(n683) );
  XNOR2_X1 U747 ( .A(KEYINPUT49), .B(n683), .ZN(n685) );
  AND2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n690) );
  XOR2_X1 U749 ( .A(KEYINPUT50), .B(KEYINPUT122), .Z(n688) );
  NAND2_X1 U750 ( .A1(n346), .A2(n686), .ZN(n687) );
  XOR2_X1 U751 ( .A(n688), .B(n687), .Z(n689) );
  NAND2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n693), .ZN(n694) );
  NOR2_X1 U755 ( .A1(n710), .A2(n694), .ZN(n705) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n705), .A2(n390), .ZN(n706) );
  XNOR2_X1 U761 ( .A(n706), .B(KEYINPUT52), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT123), .ZN(n712) );
  OR2_X1 U764 ( .A1(n710), .A2(n703), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U766 ( .A(KEYINPUT124), .B(n713), .Z(n714) );
  NAND2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n716), .A2(n345), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n717), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U770 ( .A1(n718), .A2(G478), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n722), .A2(n721), .ZN(G63) );
  XNOR2_X1 U773 ( .A(n723), .B(G101), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(n726), .ZN(n736) );
  INV_X1 U776 ( .A(n608), .ZN(n728) );
  NOR2_X1 U777 ( .A1(n728), .A2(n345), .ZN(n734) );
  NAND2_X1 U778 ( .A1(G224), .A2(n345), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n729), .B(KEYINPUT61), .ZN(n730) );
  XNOR2_X1 U780 ( .A(n730), .B(KEYINPUT127), .ZN(n731) );
  NOR2_X1 U781 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n738), .B(n737), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n674), .B(n741), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n745) );
  XOR2_X1 U787 ( .A(G227), .B(n741), .Z(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(n345), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n745), .A2(n744), .ZN(G72) );
  XOR2_X1 U791 ( .A(G137), .B(n746), .Z(G39) );
  XOR2_X1 U792 ( .A(n747), .B(G131), .Z(G33) );
endmodule

