

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766;

  NAND2_X1 U367 ( .A1(n554), .A2(n700), .ZN(n583) );
  OR2_X1 U368 ( .A1(n661), .A2(G902), .ZN(n426) );
  XNOR2_X1 U369 ( .A(n504), .B(KEYINPUT4), .ZN(n470) );
  INV_X2 U370 ( .A(G953), .ZN(n757) );
  XNOR2_X1 U371 ( .A(n538), .B(KEYINPUT1), .ZN(n569) );
  NOR2_X1 U372 ( .A1(n540), .A2(n539), .ZN(n736) );
  XNOR2_X2 U373 ( .A(n639), .B(n638), .ZN(n745) );
  AND2_X1 U374 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U375 ( .A(n566), .B(n565), .ZN(n407) );
  XNOR2_X1 U376 ( .A(n604), .B(n382), .ZN(n739) );
  NOR2_X1 U377 ( .A1(n630), .A2(n396), .ZN(n625) );
  XNOR2_X1 U378 ( .A(n520), .B(n519), .ZN(n717) );
  XNOR2_X1 U379 ( .A(n432), .B(n431), .ZN(n582) );
  XNOR2_X1 U380 ( .A(n426), .B(n349), .ZN(n521) );
  XNOR2_X1 U381 ( .A(n444), .B(n443), .ZN(n538) );
  BUF_X1 U382 ( .A(n582), .Z(n601) );
  INV_X1 U383 ( .A(KEYINPUT103), .ZN(n618) );
  XNOR2_X1 U384 ( .A(n412), .B(G110), .ZN(n464) );
  INV_X1 U385 ( .A(G119), .ZN(n412) );
  NAND2_X1 U386 ( .A1(n663), .A2(n355), .ZN(n393) );
  NAND2_X1 U387 ( .A1(n739), .A2(n348), .ZN(n380) );
  NAND2_X1 U388 ( .A1(n376), .A2(n375), .ZN(n374) );
  NOR2_X1 U389 ( .A1(n739), .A2(n606), .ZN(n375) );
  NOR2_X1 U390 ( .A1(n407), .A2(KEYINPUT79), .ZN(n406) );
  NAND2_X1 U391 ( .A1(n404), .A2(n400), .ZN(n399) );
  AND2_X1 U392 ( .A1(n401), .A2(n651), .ZN(n400) );
  NAND2_X1 U393 ( .A1(n407), .A2(n405), .ZN(n404) );
  NAND2_X1 U394 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U395 ( .A(n362), .B(n361), .ZN(n621) );
  XNOR2_X1 U396 ( .A(n470), .B(n434), .ZN(n756) );
  XNOR2_X1 U397 ( .A(G134), .B(G131), .ZN(n433) );
  OR2_X1 U398 ( .A1(n672), .A2(G902), .ZN(n444) );
  OR2_X2 U399 ( .A1(n399), .A2(n406), .ZN(n579) );
  XOR2_X1 U400 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n472) );
  XNOR2_X1 U401 ( .A(n568), .B(KEYINPUT111), .ZN(n369) );
  INV_X1 U402 ( .A(n569), .ZN(n613) );
  XNOR2_X1 U403 ( .A(n467), .B(n466), .ZN(n360) );
  AND2_X1 U404 ( .A1(n393), .A2(n346), .ZN(n384) );
  AND2_X1 U405 ( .A1(n381), .A2(n378), .ZN(n377) );
  AND2_X1 U406 ( .A1(n380), .A2(n379), .ZN(n378) );
  NAND2_X1 U407 ( .A1(n705), .A2(KEYINPUT101), .ZN(n379) );
  INV_X1 U408 ( .A(n743), .ZN(n403) );
  INV_X1 U409 ( .A(KEYINPUT79), .ZN(n402) );
  AND2_X1 U410 ( .A1(n743), .A2(KEYINPUT79), .ZN(n405) );
  INV_X1 U411 ( .A(KEYINPUT83), .ZN(n361) );
  XNOR2_X1 U412 ( .A(G116), .B(G119), .ZN(n446) );
  XNOR2_X1 U413 ( .A(G131), .B(G143), .ZN(n492) );
  XNOR2_X1 U414 ( .A(n394), .B(KEYINPUT33), .ZN(n708) );
  NAND2_X1 U415 ( .A1(n395), .A2(n601), .ZN(n394) );
  AND2_X1 U416 ( .A1(n396), .A2(n569), .ZN(n395) );
  XNOR2_X1 U417 ( .A(KEYINPUT16), .B(KEYINPUT70), .ZN(n461) );
  XNOR2_X1 U418 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n413) );
  XNOR2_X1 U419 ( .A(G128), .B(KEYINPUT91), .ZN(n415) );
  XNOR2_X1 U420 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n414) );
  NOR2_X1 U421 ( .A1(n392), .A2(n682), .ZN(n391) );
  NOR2_X1 U422 ( .A1(n410), .A2(G475), .ZN(n392) );
  XNOR2_X1 U423 ( .A(n756), .B(G146), .ZN(n450) );
  XNOR2_X1 U424 ( .A(G140), .B(G137), .ZN(n436) );
  XNOR2_X1 U425 ( .A(G110), .B(G104), .ZN(n439) );
  NAND2_X1 U426 ( .A1(n372), .A2(n745), .ZN(n363) );
  INV_X1 U427 ( .A(n579), .ZN(n372) );
  INV_X1 U428 ( .A(n759), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n477), .B(n360), .ZN(n680) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n365) );
  INV_X1 U431 ( .A(KEYINPUT36), .ZN(n366) );
  NAND2_X1 U432 ( .A1(n369), .A2(n368), .ZN(n367) );
  INV_X1 U433 ( .A(KEYINPUT31), .ZN(n382) );
  XNOR2_X1 U434 ( .A(n614), .B(KEYINPUT81), .ZN(n616) );
  NAND2_X1 U435 ( .A1(n384), .A2(n383), .ZN(n385) );
  AND2_X2 U436 ( .A1(n645), .A2(n644), .ZN(n663) );
  AND2_X1 U437 ( .A1(n645), .A2(n359), .ZN(n345) );
  AND2_X1 U438 ( .A1(n391), .A2(KEYINPUT60), .ZN(n346) );
  AND2_X1 U439 ( .A1(n644), .A2(G210), .ZN(n347) );
  NOR2_X1 U440 ( .A1(n705), .A2(KEYINPUT101), .ZN(n348) );
  XOR2_X1 U441 ( .A(n425), .B(KEYINPUT25), .Z(n349) );
  NOR2_X1 U442 ( .A1(n557), .A2(n556), .ZN(n350) );
  AND2_X1 U443 ( .A1(n645), .A2(n347), .ZN(n351) );
  XOR2_X1 U444 ( .A(KEYINPUT5), .B(G137), .Z(n352) );
  XNOR2_X1 U445 ( .A(n534), .B(n533), .ZN(n612) );
  INV_X1 U446 ( .A(n612), .ZN(n396) );
  OR2_X1 U447 ( .A1(n636), .A2(n635), .ZN(n353) );
  XNOR2_X1 U448 ( .A(KEYINPUT62), .B(n647), .ZN(n354) );
  INV_X1 U449 ( .A(KEYINPUT101), .ZN(n606) );
  AND2_X1 U450 ( .A1(n410), .A2(G475), .ZN(n355) );
  NOR2_X1 U451 ( .A1(n360), .A2(n744), .ZN(n356) );
  NAND2_X1 U452 ( .A1(n685), .A2(KEYINPUT72), .ZN(n357) );
  AND2_X1 U453 ( .A1(n659), .A2(n408), .ZN(n358) );
  NOR2_X1 U454 ( .A1(n757), .A2(G952), .ZN(n682) );
  INV_X1 U455 ( .A(n682), .ZN(n409) );
  AND2_X1 U456 ( .A1(n644), .A2(G472), .ZN(n359) );
  INV_X1 U457 ( .A(KEYINPUT60), .ZN(n408) );
  NAND2_X1 U458 ( .A1(n631), .A2(KEYINPUT44), .ZN(n362) );
  XNOR2_X2 U459 ( .A(n594), .B(KEYINPUT35), .ZN(n631) );
  NAND2_X1 U460 ( .A1(n363), .A2(KEYINPUT2), .ZN(n641) );
  XNOR2_X1 U461 ( .A(n363), .B(n685), .ZN(n721) );
  XNOR2_X2 U462 ( .A(G143), .B(G128), .ZN(n504) );
  NOR2_X1 U463 ( .A1(n535), .A2(n612), .ZN(n536) );
  XNOR2_X2 U464 ( .A(n364), .B(n646), .ZN(n534) );
  OR2_X2 U465 ( .A1(n647), .A2(G902), .ZN(n364) );
  NAND2_X1 U466 ( .A1(n365), .A2(n569), .ZN(n653) );
  INV_X1 U467 ( .A(n583), .ZN(n368) );
  INV_X1 U468 ( .A(n399), .ZN(n370) );
  NAND2_X1 U469 ( .A1(n371), .A2(n370), .ZN(n580) );
  NOR2_X1 U470 ( .A1(n406), .A2(n357), .ZN(n371) );
  XNOR2_X1 U471 ( .A(n579), .B(n373), .ZN(n758) );
  NOR2_X2 U472 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U473 ( .A1(n377), .A2(n374), .ZN(n617) );
  INV_X1 U474 ( .A(n725), .ZN(n376) );
  NAND2_X1 U475 ( .A1(n725), .A2(n348), .ZN(n381) );
  XNOR2_X1 U476 ( .A(n599), .B(n600), .ZN(n725) );
  NAND2_X1 U477 ( .A1(n393), .A2(n391), .ZN(n390) );
  NAND2_X1 U478 ( .A1(n389), .A2(n659), .ZN(n383) );
  NAND2_X1 U479 ( .A1(n386), .A2(n385), .ZN(G60) );
  NAND2_X1 U480 ( .A1(n389), .A2(n358), .ZN(n387) );
  NAND2_X1 U481 ( .A1(n390), .A2(n408), .ZN(n388) );
  INV_X1 U482 ( .A(n663), .ZN(n389) );
  XNOR2_X1 U483 ( .A(n397), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U484 ( .A1(n398), .A2(n409), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n345), .B(n354), .ZN(n398) );
  INV_X1 U486 ( .A(n659), .ZN(n410) );
  XNOR2_X1 U487 ( .A(n595), .B(KEYINPUT105), .ZN(n459) );
  INV_X1 U488 ( .A(n503), .ZN(n462) );
  XNOR2_X1 U489 ( .A(n517), .B(n516), .ZN(n654) );
  XOR2_X1 U490 ( .A(n465), .B(n447), .Z(n411) );
  INV_X1 U491 ( .A(KEYINPUT72), .ZN(n578) );
  XNOR2_X1 U492 ( .A(n531), .B(KEYINPUT46), .ZN(n563) );
  INV_X1 U493 ( .A(KEYINPUT30), .ZN(n451) );
  INV_X1 U494 ( .A(KEYINPUT82), .ZN(n622) );
  INV_X1 U495 ( .A(KEYINPUT34), .ZN(n591) );
  BUF_X1 U496 ( .A(n654), .Z(n655) );
  AND2_X2 U497 ( .A1(n616), .A2(n522), .ZN(n660) );
  XNOR2_X1 U498 ( .A(n464), .B(n413), .ZN(n417) );
  XNOR2_X1 U499 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U500 ( .A(n417), .B(n416), .ZN(n421) );
  XNOR2_X1 U501 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n419) );
  NAND2_X1 U502 ( .A1(n757), .A2(G234), .ZN(n418) );
  XNOR2_X1 U503 ( .A(n419), .B(n418), .ZN(n502) );
  NAND2_X1 U504 ( .A1(n502), .A2(G221), .ZN(n420) );
  XNOR2_X1 U505 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X1 U506 ( .A(G146), .B(G125), .ZN(n468) );
  XNOR2_X1 U507 ( .A(n468), .B(KEYINPUT10), .ZN(n488) );
  INV_X1 U508 ( .A(n436), .ZN(n422) );
  XNOR2_X1 U509 ( .A(n488), .B(n422), .ZN(n755) );
  XNOR2_X1 U510 ( .A(n423), .B(n755), .ZN(n661) );
  XNOR2_X1 U511 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  NAND2_X1 U512 ( .A1(G234), .A2(n643), .ZN(n424) );
  XNOR2_X1 U513 ( .A(KEYINPUT20), .B(n424), .ZN(n427) );
  NAND2_X1 U514 ( .A1(n427), .A2(G217), .ZN(n425) );
  NAND2_X1 U515 ( .A1(n427), .A2(G221), .ZN(n430) );
  INV_X1 U516 ( .A(KEYINPUT92), .ZN(n428) );
  XNOR2_X1 U517 ( .A(n428), .B(KEYINPUT21), .ZN(n429) );
  XNOR2_X1 U518 ( .A(n430), .B(n429), .ZN(n686) );
  NAND2_X1 U519 ( .A1(n521), .A2(n686), .ZN(n432) );
  INV_X1 U520 ( .A(KEYINPUT64), .ZN(n431) );
  XNOR2_X1 U521 ( .A(n433), .B(KEYINPUT66), .ZN(n434) );
  NAND2_X1 U522 ( .A1(n757), .A2(G227), .ZN(n435) );
  XNOR2_X1 U523 ( .A(n435), .B(KEYINPUT69), .ZN(n437) );
  XNOR2_X1 U524 ( .A(n437), .B(n436), .ZN(n441) );
  XNOR2_X1 U525 ( .A(G101), .B(G107), .ZN(n438) );
  XNOR2_X1 U526 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U527 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U528 ( .A(n450), .B(n442), .ZN(n672) );
  XNOR2_X1 U529 ( .A(KEYINPUT68), .B(G469), .ZN(n443) );
  NAND2_X1 U530 ( .A1(n582), .A2(n538), .ZN(n595) );
  XNOR2_X1 U531 ( .A(G113), .B(G101), .ZN(n445) );
  XNOR2_X1 U532 ( .A(n445), .B(KEYINPUT3), .ZN(n465) );
  XNOR2_X1 U533 ( .A(n352), .B(n446), .ZN(n447) );
  NOR2_X1 U534 ( .A1(G953), .A2(G237), .ZN(n485) );
  NAND2_X1 U535 ( .A1(n485), .A2(G210), .ZN(n448) );
  XNOR2_X1 U536 ( .A(n411), .B(n448), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n450), .B(n449), .ZN(n647) );
  INV_X1 U538 ( .A(G472), .ZN(n646) );
  OR2_X1 U539 ( .A1(G237), .A2(G902), .ZN(n478) );
  NAND2_X1 U540 ( .A1(G214), .A2(n478), .ZN(n700) );
  INV_X1 U541 ( .A(n700), .ZN(n567) );
  NOR2_X1 U542 ( .A1(n534), .A2(n567), .ZN(n452) );
  XNOR2_X1 U543 ( .A(n452), .B(n451), .ZN(n457) );
  NAND2_X1 U544 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U545 ( .A(n453), .B(KEYINPUT14), .ZN(n713) );
  NOR2_X1 U546 ( .A1(G900), .A2(n757), .ZN(n454) );
  NAND2_X1 U547 ( .A1(n454), .A2(G902), .ZN(n455) );
  NAND2_X1 U548 ( .A1(G952), .A2(n757), .ZN(n584) );
  NAND2_X1 U549 ( .A1(n455), .A2(n584), .ZN(n456) );
  NAND2_X1 U550 ( .A1(n713), .A2(n456), .ZN(n523) );
  NOR2_X1 U551 ( .A1(n457), .A2(n523), .ZN(n458) );
  NAND2_X1 U552 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X2 U553 ( .A(n460), .B(KEYINPUT73), .ZN(n552) );
  XOR2_X2 U554 ( .A(G122), .B(G104), .Z(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(n461), .ZN(n463) );
  XOR2_X1 U556 ( .A(G116), .B(G107), .Z(n503) );
  XNOR2_X1 U557 ( .A(n463), .B(n462), .ZN(n467) );
  XNOR2_X1 U558 ( .A(n464), .B(n465), .ZN(n466) );
  XNOR2_X1 U559 ( .A(n468), .B(KEYINPUT74), .ZN(n469) );
  XNOR2_X1 U560 ( .A(n470), .B(n469), .ZN(n476) );
  NAND2_X1 U561 ( .A1(G224), .A2(n757), .ZN(n471) );
  XNOR2_X1 U562 ( .A(n472), .B(n471), .ZN(n474) );
  XOR2_X1 U563 ( .A(KEYINPUT69), .B(KEYINPUT17), .Z(n473) );
  XNOR2_X1 U564 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U565 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U566 ( .A1(n680), .A2(n643), .ZN(n481) );
  INV_X1 U567 ( .A(n478), .ZN(n479) );
  INV_X1 U568 ( .A(G210), .ZN(n676) );
  NOR2_X1 U569 ( .A1(n479), .A2(n676), .ZN(n480) );
  XNOR2_X2 U570 ( .A(n481), .B(n480), .ZN(n554) );
  XNOR2_X1 U571 ( .A(KEYINPUT71), .B(KEYINPUT38), .ZN(n482) );
  XNOR2_X1 U572 ( .A(n554), .B(n482), .ZN(n701) );
  NAND2_X1 U573 ( .A1(n552), .A2(n701), .ZN(n484) );
  INV_X1 U574 ( .A(KEYINPUT39), .ZN(n483) );
  XNOR2_X1 U575 ( .A(n484), .B(n483), .ZN(n574) );
  INV_X1 U576 ( .A(n574), .ZN(n515) );
  XOR2_X1 U577 ( .A(G140), .B(G113), .Z(n487) );
  NAND2_X1 U578 ( .A1(G214), .A2(n485), .ZN(n486) );
  XNOR2_X1 U579 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U580 ( .A(n489), .B(n488), .ZN(n497) );
  XOR2_X1 U581 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n491) );
  XNOR2_X1 U582 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n490) );
  XNOR2_X1 U583 ( .A(n491), .B(n490), .ZN(n495) );
  XNOR2_X1 U584 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U585 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U586 ( .A(n497), .B(n496), .ZN(n658) );
  INV_X1 U587 ( .A(G902), .ZN(n498) );
  NAND2_X1 U588 ( .A1(n658), .A2(n498), .ZN(n500) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(G475), .ZN(n499) );
  XNOR2_X1 U590 ( .A(n500), .B(n499), .ZN(n556) );
  INV_X1 U591 ( .A(KEYINPUT96), .ZN(n501) );
  XNOR2_X1 U592 ( .A(n556), .B(n501), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n502), .A2(G217), .ZN(n506) );
  XNOR2_X1 U594 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U595 ( .A(n506), .B(n505), .ZN(n512) );
  XOR2_X1 U596 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n508) );
  XNOR2_X1 U597 ( .A(G134), .B(G122), .ZN(n507) );
  XNOR2_X1 U598 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U599 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n509) );
  XNOR2_X1 U600 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U601 ( .A(n512), .B(n511), .ZN(n666) );
  OR2_X1 U602 ( .A1(n666), .A2(G902), .ZN(n514) );
  XNOR2_X1 U603 ( .A(KEYINPUT99), .B(G478), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n514), .B(n513), .ZN(n557) );
  AND2_X1 U605 ( .A1(n541), .A2(n557), .ZN(n738) );
  NAND2_X1 U606 ( .A1(n515), .A2(n738), .ZN(n517) );
  XNOR2_X1 U607 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n516) );
  NAND2_X1 U608 ( .A1(n701), .A2(n700), .ZN(n518) );
  XNOR2_X1 U609 ( .A(KEYINPUT108), .B(n518), .ZN(n704) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n703) );
  OR2_X1 U611 ( .A1(n704), .A2(n703), .ZN(n520) );
  XNOR2_X1 U612 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n519) );
  BUF_X1 U613 ( .A(n521), .Z(n522) );
  INV_X1 U614 ( .A(n522), .ZN(n615) );
  INV_X1 U615 ( .A(n686), .ZN(n524) );
  NOR2_X1 U616 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U617 ( .A1(n615), .A2(n525), .ZN(n535) );
  NOR2_X1 U618 ( .A1(n534), .A2(n535), .ZN(n527) );
  XNOR2_X1 U619 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U621 ( .A1(n528), .A2(n538), .ZN(n540) );
  NOR2_X1 U622 ( .A1(n717), .A2(n540), .ZN(n530) );
  XNOR2_X1 U623 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n529) );
  XNOR2_X1 U624 ( .A(n530), .B(n529), .ZN(n764) );
  NOR2_X2 U625 ( .A1(n654), .A2(n764), .ZN(n531) );
  INV_X1 U626 ( .A(KEYINPUT102), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT6), .ZN(n533) );
  XNOR2_X1 U628 ( .A(KEYINPUT104), .B(n536), .ZN(n537) );
  NAND2_X1 U629 ( .A1(n537), .A2(n738), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT19), .B(n583), .Z(n539) );
  INV_X1 U631 ( .A(KEYINPUT76), .ZN(n543) );
  NAND2_X1 U632 ( .A1(n736), .A2(n543), .ZN(n546) );
  OR2_X1 U633 ( .A1(n541), .A2(n557), .ZN(n649) );
  INV_X1 U634 ( .A(KEYINPUT100), .ZN(n542) );
  XNOR2_X1 U635 ( .A(n649), .B(n542), .ZN(n576) );
  OR2_X1 U636 ( .A1(n576), .A2(n738), .ZN(n605) );
  NAND2_X1 U637 ( .A1(n605), .A2(KEYINPUT47), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U640 ( .A1(n605), .A2(n736), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n547), .B(KEYINPUT47), .ZN(n548) );
  NAND2_X1 U642 ( .A1(n548), .A2(KEYINPUT76), .ZN(n549) );
  AND2_X1 U643 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U644 ( .A1(n653), .A2(n551), .ZN(n561) );
  BUF_X1 U645 ( .A(n552), .Z(n553) );
  INV_X1 U646 ( .A(n553), .ZN(n559) );
  BUF_X1 U647 ( .A(n554), .Z(n555) );
  INV_X1 U648 ( .A(n555), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n555), .A2(n350), .ZN(n558) );
  OR2_X1 U650 ( .A1(n559), .A2(n558), .ZN(n648) );
  XNOR2_X1 U651 ( .A(n648), .B(KEYINPUT77), .ZN(n560) );
  NOR2_X1 U652 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U653 ( .A1(n563), .A2(n562), .ZN(n566) );
  XNOR2_X1 U654 ( .A(KEYINPUT80), .B(KEYINPUT48), .ZN(n564) );
  XNOR2_X1 U655 ( .A(n564), .B(KEYINPUT67), .ZN(n565) );
  NOR2_X1 U656 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n570), .A2(n613), .ZN(n571) );
  XNOR2_X1 U658 ( .A(n571), .B(KEYINPUT43), .ZN(n573) );
  NAND2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n743) );
  BUF_X1 U660 ( .A(n574), .Z(n575) );
  INV_X1 U661 ( .A(n575), .ZN(n577) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n651) );
  NAND2_X1 U663 ( .A1(n579), .A2(n578), .ZN(n581) );
  INV_X1 U664 ( .A(KEYINPUT2), .ZN(n685) );
  NAND2_X1 U665 ( .A1(n581), .A2(n580), .ZN(n640) );
  XNOR2_X1 U666 ( .A(n583), .B(KEYINPUT19), .ZN(n588) );
  XOR2_X1 U667 ( .A(G898), .B(KEYINPUT87), .Z(n749) );
  NOR2_X1 U668 ( .A1(n749), .A2(n757), .ZN(n744) );
  NAND2_X1 U669 ( .A1(n744), .A2(G902), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n585), .A2(n584), .ZN(n586) );
  AND2_X1 U671 ( .A1(n586), .A2(n713), .ZN(n587) );
  NAND2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X2 U673 ( .A(n589), .B(KEYINPUT0), .ZN(n609) );
  XNOR2_X1 U674 ( .A(n609), .B(KEYINPUT88), .ZN(n598) );
  INV_X1 U675 ( .A(n598), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n708), .A2(n590), .ZN(n592) );
  XNOR2_X1 U677 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n593), .A2(n350), .ZN(n594) );
  INV_X1 U679 ( .A(KEYINPUT93), .ZN(n600) );
  INV_X1 U680 ( .A(n595), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n596), .A2(n534), .ZN(n597) );
  NOR2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U683 ( .A(n534), .ZN(n602) );
  AND2_X1 U684 ( .A1(n601), .A2(n602), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n569), .A2(n603), .ZN(n694) );
  NOR2_X1 U686 ( .A1(n609), .A2(n694), .ZN(n604) );
  INV_X1 U687 ( .A(n605), .ZN(n705) );
  INV_X1 U688 ( .A(n703), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n686), .A2(n607), .ZN(n608) );
  NOR2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n611) );
  INV_X1 U691 ( .A(KEYINPUT22), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n611), .B(n610), .ZN(n630) );
  NAND2_X1 U693 ( .A1(n625), .A2(n613), .ZN(n614) );
  NOR2_X1 U694 ( .A1(n617), .A2(n660), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(n637) );
  AND2_X1 U698 ( .A1(n615), .A2(n569), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U700 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n765) );
  NAND2_X1 U702 ( .A1(n534), .A2(n615), .ZN(n628) );
  OR2_X1 U703 ( .A1(n569), .A2(n628), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n732) );
  OR2_X1 U705 ( .A1(n765), .A2(n732), .ZN(n634) );
  NOR2_X1 U706 ( .A1(n634), .A2(n631), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n632), .A2(KEYINPUT44), .ZN(n636) );
  INV_X1 U708 ( .A(KEYINPUT44), .ZN(n633) );
  NOR2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n637), .A2(n353), .ZN(n639) );
  XNOR2_X1 U711 ( .A(KEYINPUT78), .B(KEYINPUT45), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n640), .A2(n745), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n645) );
  INV_X1 U714 ( .A(n643), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n648), .B(G143), .ZN(G45) );
  INV_X1 U716 ( .A(n649), .ZN(n733) );
  NAND2_X1 U717 ( .A1(n739), .A2(n733), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(G116), .ZN(G18) );
  XNOR2_X1 U719 ( .A(n651), .B(G134), .ZN(G36) );
  XOR2_X1 U720 ( .A(G125), .B(KEYINPUT37), .Z(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(G27) );
  XOR2_X1 U722 ( .A(n655), .B(G131), .Z(G33) );
  XOR2_X1 U723 ( .A(G122), .B(KEYINPUT126), .Z(n656) );
  XNOR2_X1 U724 ( .A(n631), .B(n656), .ZN(G24) );
  XOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n657) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(n660), .B(G101), .Z(G3) );
  BUF_X1 U728 ( .A(n661), .Z(n662) );
  NAND2_X1 U729 ( .A1(n663), .A2(G217), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n662), .B(n664), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n665), .A2(n682), .ZN(G66) );
  NAND2_X1 U732 ( .A1(n663), .A2(G478), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n666), .B(KEYINPUT122), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n669), .A2(n682), .ZN(G63) );
  NAND2_X1 U736 ( .A1(n663), .A2(G469), .ZN(n674) );
  XOR2_X1 U737 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT58), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n675), .A2(n682), .ZN(G54) );
  XNOR2_X1 U742 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n678) );
  XNOR2_X1 U743 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n351), .B(n681), .ZN(n683) );
  XNOR2_X1 U747 ( .A(n684), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U748 ( .A1(n522), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n688), .B(n687), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n689), .A2(n534), .ZN(n692) );
  NOR2_X1 U752 ( .A1(n569), .A2(n601), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n690), .B(KEYINPUT50), .ZN(n691) );
  NOR2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U755 ( .A(KEYINPUT117), .B(n693), .Z(n696) );
  INV_X1 U756 ( .A(n694), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U758 ( .A(n697), .B(KEYINPUT51), .Z(n698) );
  NOR2_X1 U759 ( .A1(n717), .A2(n698), .ZN(n699) );
  XNOR2_X1 U760 ( .A(n699), .B(KEYINPUT118), .ZN(n711) );
  NOR2_X1 U761 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U765 ( .A(n708), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n709), .A2(n716), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n712), .B(KEYINPUT52), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n713), .A2(G952), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n722), .B(KEYINPUT119), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n723), .A2(n757), .ZN(n724) );
  XOR2_X1 U776 ( .A(KEYINPUT53), .B(n724), .Z(G75) );
  NAND2_X1 U777 ( .A1(n725), .A2(n738), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n726), .B(G104), .ZN(G6) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n728) );
  NAND2_X1 U780 ( .A1(n725), .A2(n733), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n728), .B(n727), .ZN(n729) );
  XOR2_X1 U782 ( .A(n729), .B(KEYINPUT26), .Z(n731) );
  XNOR2_X1 U783 ( .A(G107), .B(KEYINPUT112), .ZN(n730) );
  XNOR2_X1 U784 ( .A(n731), .B(n730), .ZN(G9) );
  XOR2_X1 U785 ( .A(G110), .B(n732), .Z(G12) );
  XOR2_X1 U786 ( .A(G128), .B(KEYINPUT29), .Z(n735) );
  NAND2_X1 U787 ( .A1(n736), .A2(n733), .ZN(n734) );
  XNOR2_X1 U788 ( .A(n735), .B(n734), .ZN(G30) );
  NAND2_X1 U789 ( .A1(n736), .A2(n738), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n737), .B(G146), .ZN(G48) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT114), .ZN(n741) );
  XNOR2_X1 U793 ( .A(G113), .B(n741), .ZN(G15) );
  XOR2_X1 U794 ( .A(G140), .B(KEYINPUT115), .Z(n742) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(G42) );
  NAND2_X1 U796 ( .A1(n745), .A2(n757), .ZN(n752) );
  XOR2_X1 U797 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n747) );
  NAND2_X1 U798 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U800 ( .A(KEYINPUT123), .B(n748), .ZN(n750) );
  NAND2_X1 U801 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U803 ( .A(n753), .B(KEYINPUT125), .Z(n754) );
  XNOR2_X1 U804 ( .A(n356), .B(n754), .ZN(G69) );
  XOR2_X1 U805 ( .A(n756), .B(n755), .Z(n759) );
  NAND2_X1 U806 ( .A1(n758), .A2(n757), .ZN(n763) );
  XOR2_X1 U807 ( .A(G227), .B(n759), .Z(n760) );
  NAND2_X1 U808 ( .A1(n760), .A2(G900), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(G953), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n763), .A2(n762), .ZN(G72) );
  XOR2_X1 U811 ( .A(n764), .B(G137), .Z(G39) );
  XNOR2_X1 U812 ( .A(G119), .B(KEYINPUT127), .ZN(n766) );
  XNOR2_X1 U813 ( .A(n766), .B(n765), .ZN(G21) );
endmodule

