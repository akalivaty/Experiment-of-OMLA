//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT1), .B2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT73), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT74), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n208), .B(new_n210), .C1(G113gat), .C2(new_n209), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n205), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217));
  XNOR2_X1  g016(.A(G141gat), .B(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(G155gat), .B2(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G155gat), .B(G162gat), .ZN(new_n222));
  XOR2_X1   g021(.A(new_n221), .B(new_n222), .Z(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT4), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT81), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n205), .A2(new_n215), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n226), .B2(new_n223), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n229), .B(new_n223), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT5), .B1(new_n234), .B2(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n225), .A2(new_n231), .A3(KEYINPUT5), .A4(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT0), .ZN(new_n240));
  XNOR2_X1  g039(.A(G57gat), .B(G85gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n240), .B(new_n241), .Z(new_n242));
  AOI21_X1  g041(.A(KEYINPUT6), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n242), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n244), .A3(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n236), .A2(KEYINPUT6), .A3(new_n244), .A4(new_n237), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G169gat), .ZN(new_n253));
  INV_X1    g052(.A(G176gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT23), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G169gat), .B2(G176gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT67), .Z(new_n261));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT24), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n263), .B2(new_n262), .ZN(new_n265));
  INV_X1    g064(.A(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT71), .B1(new_n266), .B2(new_n267), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n261), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n249), .B1(new_n258), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n272), .A2(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT24), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n277), .A2(new_n268), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n252), .A2(new_n249), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n260), .B(KEYINPUT67), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT66), .B(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(KEYINPUT23), .A3(new_n253), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n266), .B2(KEYINPUT27), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n267), .B(new_n288), .C1(new_n289), .C2(new_n287), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G190gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n290), .A2(new_n291), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n252), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n262), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n276), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n276), .A2(new_n298), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT29), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n303), .B2(new_n300), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT78), .B(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n308), .B2(KEYINPUT22), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n311), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n301), .B(new_n316), .C1(new_n303), .C2(new_n300), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(KEYINPUT79), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n315), .B1(new_n312), .B2(new_n317), .ZN(new_n325));
  INV_X1    g124(.A(new_n318), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(KEYINPUT30), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n248), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G22gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n311), .B1(new_n228), .B2(KEYINPUT29), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT81), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n227), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n316), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT84), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n226), .B1(new_n311), .B2(KEYINPUT29), .ZN(new_n341));
  INV_X1    g140(.A(new_n223), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n343), .A2(KEYINPUT83), .ZN(new_n344));
  INV_X1    g143(.A(G228gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  AOI211_X1 g145(.A(new_n345), .B(new_n346), .C1(new_n343), .C2(KEYINPUT83), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n335), .A2(new_n340), .A3(new_n344), .A4(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT31), .B(G50gat), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n311), .A2(KEYINPUT82), .ZN(new_n351));
  INV_X1    g150(.A(new_n310), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n309), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n351), .B(new_n338), .C1(KEYINPUT82), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n223), .B1(new_n354), .B2(new_n226), .ZN(new_n355));
  OAI22_X1  g154(.A1(new_n339), .A2(new_n355), .B1(new_n345), .B2(new_n346), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n348), .A2(new_n350), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n350), .B1(new_n348), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n332), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n349), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n348), .A2(new_n350), .A3(new_n356), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n331), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n299), .A2(new_n216), .ZN(new_n364));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT64), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n302), .A2(new_n229), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT32), .ZN(new_n369));
  XNOR2_X1  g168(.A(G15gat), .B(G43gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT77), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n368), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n368), .B2(new_n375), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n369), .B(new_n373), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(KEYINPUT33), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n367), .ZN(new_n382));
  INV_X1    g181(.A(new_n366), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT34), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n384), .B(KEYINPUT34), .Z(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n380), .A3(new_n378), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n359), .A2(new_n363), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT35), .B1(new_n329), .B2(new_n389), .ZN(new_n390));
  AND4_X1   g189(.A1(new_n386), .A2(new_n359), .A3(new_n363), .A4(new_n388), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT35), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n248), .A4(new_n328), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT85), .B(KEYINPUT40), .Z(new_n395));
  INV_X1    g194(.A(KEYINPUT39), .ZN(new_n396));
  INV_X1    g195(.A(new_n232), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n224), .B(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n228), .A2(new_n230), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n396), .B(new_n397), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n242), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n234), .A2(new_n232), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT39), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n225), .A2(new_n231), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(new_n397), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n395), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT86), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(new_n395), .C1(new_n402), .C2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n324), .A2(new_n327), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n402), .A2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT40), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n245), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n359), .A2(new_n363), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n312), .A2(new_n317), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT37), .ZN(new_n419));
  INV_X1    g218(.A(new_n315), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n312), .A2(new_n421), .A3(new_n317), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n326), .B1(new_n423), .B2(KEYINPUT38), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT38), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n419), .A2(new_n425), .A3(new_n420), .A4(new_n422), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n246), .A2(new_n424), .A3(new_n247), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n329), .A2(new_n416), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT36), .ZN(new_n430));
  INV_X1    g229(.A(new_n388), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n387), .B1(new_n378), .B2(new_n380), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n386), .A2(KEYINPUT36), .A3(new_n388), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n394), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G197gat), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT11), .B(G169gat), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT12), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G22gat), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(G1gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G8gat), .ZN(new_n448));
  INV_X1    g247(.A(G1gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT16), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  OAI21_X1  g252(.A(G8gat), .B1(new_n453), .B2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n452), .B2(new_n454), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G50gat), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n459), .A2(G43gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(G43gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT15), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(G29gat), .A2(G36gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT14), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(KEYINPUT15), .A3(new_n461), .ZN(new_n468));
  NAND2_X1  g267(.A1(G29gat), .A2(G36gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n468), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n465), .B(KEYINPUT14), .ZN(new_n473));
  INV_X1    g272(.A(new_n469), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n471), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n471), .B2(new_n475), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n443), .B1(new_n458), .B2(new_n479), .ZN(new_n480));
  OAI221_X1 g279(.A(KEYINPUT90), .B1(new_n477), .B2(new_n478), .C1(new_n456), .C2(new_n457), .ZN(new_n481));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n452), .A2(new_n454), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n471), .A2(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT18), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n442), .B1(new_n488), .B2(KEYINPUT91), .ZN(new_n489));
  INV_X1    g288(.A(new_n457), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n484), .A2(KEYINPUT17), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n475), .A3(new_n476), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n494), .A2(KEYINPUT90), .B1(new_n484), .B2(new_n483), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(KEYINPUT18), .A3(new_n482), .A4(new_n480), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n483), .B(new_n484), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT13), .Z(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n488), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n486), .A2(new_n487), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n486), .B2(new_n487), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n502), .B(new_n496), .C1(new_n504), .C2(new_n442), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT7), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(G85gat), .A3(G92gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513));
  INV_X1    g312(.A(G85gat), .ZN(new_n514));
  INV_X1    g313(.A(G92gat), .ZN(new_n515));
  AOI22_X1  g314(.A1(KEYINPUT8), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G99gat), .B(G106gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n512), .B2(new_n516), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n484), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT41), .ZN(new_n523));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT96), .ZN(new_n525));
  OAI221_X1 g324(.A(new_n522), .B1(new_n523), .B2(new_n525), .C1(new_n479), .C2(new_n521), .ZN(new_n526));
  XOR2_X1   g325(.A(G190gat), .B(G218gat), .Z(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n523), .ZN(new_n529));
  XOR2_X1   g328(.A(G134gat), .B(G162gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(new_n531), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  XNOR2_X1  g337(.A(G71gat), .B(G78gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n541));
  INV_X1    g340(.A(G57gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G57gat), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(KEYINPUT93), .B(new_n540), .C1(new_n546), .C2(KEYINPUT92), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548));
  NAND2_X1  g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n544), .A2(G57gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n542), .A2(G64gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n539), .B1(new_n546), .B2(KEYINPUT93), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n547), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n521), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n512), .A2(new_n516), .ZN(new_n560));
  INV_X1    g359(.A(new_n517), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n518), .ZN(new_n563));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n548), .B1(new_n564), .B2(new_n541), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n545), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT92), .B1(new_n566), .B2(new_n551), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n539), .B(new_n565), .C1(new_n567), .C2(new_n548), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n568), .A3(new_n547), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n559), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT98), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n576), .A3(new_n569), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n521), .A3(KEYINPUT10), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n571), .B(KEYINPUT99), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI211_X1 g381(.A(KEYINPUT100), .B(new_n580), .C1(new_n577), .C2(new_n578), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n538), .B1(new_n574), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n577), .A2(KEYINPUT97), .A3(new_n578), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT97), .B1(new_n577), .B2(new_n578), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n586), .A2(new_n587), .A3(new_n571), .ZN(new_n588));
  INV_X1    g387(.A(new_n538), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n588), .A2(new_n573), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n558), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(G231gat), .B(G233gat), .C1(new_n558), .C2(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n597), .A2(new_n599), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G183gat), .B(G211gat), .Z(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n454), .B(new_n452), .C1(new_n592), .C2(new_n593), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n608), .B2(new_n612), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n535), .B(new_n591), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n437), .A2(new_n507), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(new_n248), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(new_n449), .ZN(G1324gat));
  XNOR2_X1  g419(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n621));
  INV_X1    g420(.A(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n412), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT16), .B(G8gat), .Z(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT102), .Z(new_n625));
  OAI21_X1  g424(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(G8gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(KEYINPUT42), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n626), .B(new_n627), .C1(new_n623), .C2(new_n628), .ZN(G1325gat));
  NOR2_X1   g428(.A1(new_n431), .A2(new_n432), .ZN(new_n630));
  AOI21_X1  g429(.A(G15gat), .B1(new_n622), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n435), .A2(KEYINPUT103), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n433), .A2(new_n434), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G15gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT104), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n631), .B1(new_n622), .B2(new_n637), .ZN(G1326gat));
  OR3_X1    g437(.A1(new_n618), .A2(KEYINPUT105), .A3(new_n417), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT105), .B1(new_n618), .B2(new_n417), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT43), .B(G22gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  NOR2_X1   g442(.A1(new_n614), .A2(new_n615), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n591), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g446(.A1(new_n437), .A2(new_n507), .A3(new_n534), .A4(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G29gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n248), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT45), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n534), .A2(KEYINPUT44), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n437), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n647), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n506), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n632), .A2(new_n428), .A3(new_n429), .A4(new_n634), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n535), .B1(new_n657), .B2(new_n394), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n654), .B(new_n656), .C1(new_n658), .C2(KEYINPUT44), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n659), .A2(new_n660), .A3(new_n248), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n659), .B2(new_n248), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G29gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n652), .B1(new_n661), .B2(new_n663), .ZN(G1328gat));
  AOI21_X1  g463(.A(G36gat), .B1(KEYINPUT107), .B2(KEYINPUT46), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n412), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G36gat), .B1(new_n659), .B2(new_n328), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1329gat));
  INV_X1    g469(.A(new_n634), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n633), .B1(new_n433), .B2(new_n434), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G43gat), .B1(new_n659), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G43gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n648), .A2(new_n677), .A3(new_n630), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n674), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(G1330gat));
  OAI21_X1  g480(.A(G50gat), .B1(new_n659), .B2(new_n417), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT48), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n648), .A2(new_n459), .A3(new_n416), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(G1331gat));
  NAND2_X1  g486(.A1(new_n657), .A2(new_n394), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n608), .A2(new_n612), .ZN(new_n689));
  INV_X1    g488(.A(new_n611), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n534), .B1(new_n691), .B2(new_n613), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n692), .A2(new_n506), .A3(new_n646), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n248), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n542), .ZN(G1332gat));
  AND2_X1   g495(.A1(new_n688), .A2(new_n693), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n698));
  AND2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n697), .B(new_n412), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n694), .A2(new_n328), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n698), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n702), .A2(new_n698), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n705), .B2(new_n700), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(G1333gat));
  NAND3_X1  g506(.A1(new_n697), .A2(G71gat), .A3(new_n635), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n630), .B(KEYINPUT110), .Z(new_n709));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(G71gat), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n416), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g513(.A1(new_n650), .A2(new_n514), .A3(new_n646), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT112), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n645), .A2(new_n507), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n658), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n658), .A2(KEYINPUT51), .A3(new_n717), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n720), .A2(KEYINPUT111), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT111), .B1(new_n720), .B2(new_n721), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n645), .A2(new_n507), .A3(new_n591), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n654), .B(new_n725), .C1(new_n658), .C2(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n248), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(G1336gat));
  OAI21_X1  g527(.A(G92gat), .B1(new_n726), .B2(new_n328), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n328), .A2(G92gat), .A3(new_n591), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n658), .A2(KEYINPUT51), .A3(new_n717), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT51), .B1(new_n658), .B2(new_n717), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT52), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(G1337gat));
  NOR4_X1   g537(.A1(new_n431), .A2(new_n432), .A3(G99gat), .A4(new_n591), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n722), .B2(new_n723), .ZN(new_n740));
  OAI21_X1  g539(.A(G99gat), .B1(new_n726), .B2(new_n673), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1338gat));
  OAI21_X1  g541(.A(G106gat), .B1(new_n726), .B2(new_n417), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n417), .A2(G106gat), .A3(new_n591), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n731), .B2(new_n732), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT53), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n743), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1339gat));
  NAND3_X1  g549(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT54), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT114), .B1(new_n588), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT97), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n571), .B1(new_n579), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n577), .A2(KEYINPUT97), .A3(new_n578), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  INV_X1    g557(.A(new_n752), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n582), .B2(new_n583), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n589), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n763), .A2(KEYINPUT55), .A3(new_n589), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n590), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n507), .B(new_n768), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n482), .B1(new_n495), .B2(new_n480), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n497), .A2(new_n498), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n441), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n442), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n500), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n591), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n534), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n768), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n761), .A2(new_n769), .ZN(new_n783));
  INV_X1    g582(.A(new_n590), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n535), .A2(new_n778), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n644), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n616), .B2(new_n507), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n692), .A2(KEYINPUT113), .A3(new_n506), .A4(new_n591), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n389), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n248), .A2(new_n412), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n507), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT116), .B(G113gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1340gat));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n646), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n645), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g605(.A(new_n535), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n808), .B(new_n809), .Z(G1343gat));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n632), .A2(new_n634), .A3(new_n798), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n792), .A2(new_n796), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n506), .A2(G141gat), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n416), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n815), .B2(KEYINPUT119), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(KEYINPUT119), .B2(new_n815), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT57), .B1(new_n813), .B2(new_n416), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n416), .A2(KEYINPUT57), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n764), .B1(new_n753), .B2(new_n760), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n783), .B(new_n784), .C1(new_n820), .C2(KEYINPUT55), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n768), .A2(KEYINPUT117), .A3(new_n770), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n507), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n534), .B1(new_n825), .B2(new_n780), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n644), .B1(new_n826), .B2(new_n791), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n819), .B1(new_n827), .B2(new_n796), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n507), .B(new_n812), .C1(new_n818), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G141gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n817), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n815), .B(KEYINPUT118), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(G141gat), .B2(new_n829), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n833), .B2(new_n811), .ZN(G1344gat));
  INV_X1    g633(.A(G148gat), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(KEYINPUT59), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n812), .B1(new_n818), .B2(new_n828), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n591), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT121), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n836), .C1(new_n837), .C2(new_n591), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n616), .A2(new_n507), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n417), .B1(new_n827), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n789), .A2(new_n790), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n779), .B1(new_n789), .B2(new_n507), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n534), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(new_n644), .B1(new_n794), .B2(new_n795), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n844), .A2(KEYINPUT57), .B1(new_n848), .B2(new_n819), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n812), .A2(new_n646), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT59), .B1(new_n851), .B2(new_n835), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n839), .A2(new_n841), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n848), .A2(new_n417), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n854), .A3(new_n835), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT120), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(G1345gat));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n812), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n644), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(G155gat), .ZN(new_n860));
  INV_X1    g659(.A(new_n837), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n645), .A2(G155gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(G1346gat));
  OR3_X1    g662(.A1(new_n858), .A2(G162gat), .A3(new_n535), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT122), .B1(new_n837), .B2(new_n535), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G162gat), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n837), .A2(KEYINPUT122), .A3(new_n535), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n650), .A2(new_n328), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n709), .A2(new_n416), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n813), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n253), .A3(new_n506), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n797), .A2(KEYINPUT123), .A3(new_n869), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT123), .B1(new_n797), .B2(new_n869), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n507), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n873), .B1(new_n878), .B2(new_n253), .ZN(G1348gat));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880));
  AOI21_X1  g679(.A(G176gat), .B1(new_n877), .B2(new_n646), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n872), .A2(new_n284), .A3(new_n591), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n876), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n874), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n254), .B1(new_n885), .B2(new_n591), .ZN(new_n886));
  INV_X1    g685(.A(new_n882), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(KEYINPUT124), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n883), .A2(new_n888), .ZN(G1349gat));
  NOR2_X1   g688(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n890));
  OAI21_X1  g689(.A(G183gat), .B1(new_n872), .B2(new_n644), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n797), .A2(new_n289), .A3(new_n645), .A4(new_n869), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n872), .B2(new_n535), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n267), .A3(new_n534), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1351gat));
  NOR4_X1   g698(.A1(new_n848), .A2(new_n417), .A3(new_n635), .A4(new_n870), .ZN(new_n900));
  INV_X1    g699(.A(G197gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n507), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n673), .A2(new_n507), .A3(new_n869), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n506), .B1(new_n821), .B2(new_n822), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n779), .B1(new_n905), .B2(new_n824), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n845), .B1(new_n906), .B2(new_n534), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n842), .B1(new_n907), .B2(new_n644), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(new_n417), .ZN(new_n909));
  INV_X1    g708(.A(new_n819), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n813), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n903), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913));
  OAI21_X1  g712(.A(G197gat), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT126), .B(new_n903), .C1(new_n909), .C2(new_n911), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT127), .B(new_n902), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1352gat));
  INV_X1    g719(.A(G204gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n900), .A2(new_n921), .A3(new_n646), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n635), .A2(new_n870), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n849), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(new_n646), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n923), .B(new_n924), .C1(new_n927), .C2(new_n921), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n900), .A2(new_n307), .A3(new_n645), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n849), .A2(new_n645), .A3(new_n925), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n900), .B2(new_n534), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n535), .A2(new_n306), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n926), .B2(new_n935), .ZN(G1355gat));
endmodule


