//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT96), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(new_n211), .B2(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n215), .A2(KEYINPUT94), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n214), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT94), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n212), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT95), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT17), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT17), .B1(new_n226), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n209), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n207), .B(G8gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n226), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n222), .A2(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n223), .B2(new_n222), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n239), .A2(new_n212), .B1(new_n213), .B2(new_n216), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n241), .A3(KEYINPUT98), .ZN(new_n242));
  OR3_X1    g041(.A1(new_n209), .A2(KEYINPUT98), .A3(new_n240), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT97), .B(KEYINPUT13), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(new_n232), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n234), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n237), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G169gat), .B(G197gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT93), .ZN(new_n250));
  XOR2_X1   g049(.A(G113gat), .B(G141gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT12), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT99), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n237), .A2(new_n246), .A3(new_n255), .A4(new_n247), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n248), .A2(KEYINPUT99), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G78gat), .B(G106gat), .Z(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT31), .B(G50gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  INV_X1    g066(.A(G148gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(G141gat), .ZN(new_n269));
  INV_X1    g068(.A(G141gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(G141gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT77), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n269), .A2(new_n271), .A3(new_n275), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285));
  INV_X1    g084(.A(new_n281), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n278), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n270), .A2(G148gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n272), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT78), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n291), .B1(new_n277), .B2(new_n283), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT78), .A3(new_n285), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G211gat), .B(G218gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(G211gat), .ZN(new_n302));
  INV_X1    g101(.A(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT73), .B(new_n300), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G211gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n303), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n311), .B2(KEYINPUT22), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n299), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n266), .B1(new_n298), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT78), .B1(new_n296), .B2(new_n285), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n282), .B1(new_n274), .B2(new_n276), .ZN(new_n319));
  NOR4_X1   g118(.A1(new_n319), .A2(new_n294), .A3(KEYINPUT3), .A4(new_n291), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n306), .A2(new_n314), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT84), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n285), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n284), .A2(new_n292), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n316), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G22gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n324), .B(KEYINPUT82), .Z(new_n330));
  NAND2_X1  g129(.A1(new_n295), .A2(new_n297), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n315), .B1(new_n331), .B2(new_n317), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n312), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n304), .A2(KEYINPUT83), .A3(new_n305), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n300), .A3(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(new_n317), .C1(new_n300), .C2(new_n334), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n296), .B1(new_n337), .B2(new_n285), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n330), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n328), .A2(new_n329), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n329), .B1(new_n328), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n265), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT85), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344));
  INV_X1    g143(.A(new_n324), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT3), .B1(new_n315), .B2(new_n317), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n296), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n322), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n266), .ZN(new_n349));
  INV_X1    g148(.A(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n348), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n349), .A2(new_n323), .B1(new_n351), .B2(new_n330), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n344), .B1(new_n352), .B2(new_n329), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n265), .B1(new_n352), .B2(new_n329), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n341), .A2(KEYINPUT86), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(new_n265), .C1(new_n340), .C2(new_n341), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(G169gat), .ZN(new_n364));
  INV_X1    g163(.A(G176gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT23), .ZN(new_n366));
  AND3_X1   g165(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT65), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT24), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(G183gat), .A3(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n372), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n366), .B(KEYINPUT65), .C1(new_n367), .C2(new_n368), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT23), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n371), .A2(new_n381), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n374), .A2(new_n376), .B1(new_n372), .B2(new_n373), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n366), .B(new_n384), .C1(new_n367), .C2(new_n368), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n378), .A2(new_n379), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT27), .B(G183gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n372), .A2(KEYINPUT27), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G183gat), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n396), .A3(new_n398), .A4(new_n379), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n393), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n372), .A2(new_n373), .ZN(new_n402));
  NOR2_X1   g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT26), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n367), .A2(new_n368), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n386), .A2(new_n390), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n363), .B1(new_n407), .B2(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n390), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n401), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n363), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n408), .A2(new_n413), .A3(new_n322), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n322), .B1(new_n408), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n362), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT74), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT74), .B(new_n362), .C1(new_n414), .C2(new_n415), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n414), .A2(new_n415), .A3(new_n362), .ZN(new_n422));
  INV_X1    g221(.A(new_n362), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n315), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n413), .A3(new_n322), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n422), .B1(KEYINPUT30), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT0), .ZN(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  XOR2_X1   g232(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n434));
  INV_X1    g233(.A(G120gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G113gat), .ZN(new_n436));
  INV_X1    g235(.A(G113gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G120gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440));
  INV_X1    g239(.A(G134gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G127gat), .ZN(new_n442));
  INV_X1    g241(.A(G127gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G134gat), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n439), .A2(new_n440), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n444), .ZN(new_n446));
  XNOR2_X1  g245(.A(G113gat), .B(G120gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n318), .B2(new_n320), .ZN(new_n452));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n284), .A2(new_n292), .A3(new_n450), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n296), .A2(KEYINPUT4), .A3(new_n450), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT4), .B1(new_n296), .B2(new_n450), .ZN(new_n462));
  NOR4_X1   g261(.A1(new_n319), .A2(new_n449), .A3(new_n458), .A4(new_n291), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT79), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n452), .B(new_n455), .C1(new_n461), .C2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n449), .B1(new_n319), .B2(new_n291), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n449), .B1(new_n296), .B2(new_n285), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n295), .B2(new_n297), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(new_n460), .A3(new_n453), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT5), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n433), .B(new_n434), .C1(new_n465), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n465), .A2(new_n472), .ZN(new_n474));
  INV_X1    g273(.A(new_n433), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n472), .A3(new_n433), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n434), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n477), .A2(new_n434), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT81), .A3(new_n476), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n429), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n409), .A2(new_n450), .A3(new_n410), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n450), .B1(new_n409), .B2(new_n410), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G43gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n488), .B(KEYINPUT32), .C1(new_n489), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n488), .B2(KEYINPUT32), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n411), .A2(new_n449), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n407), .A2(new_n450), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n484), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT33), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT68), .B1(new_n488), .B2(new_n489), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n494), .B(new_n495), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n499), .B1(new_n498), .B2(KEYINPUT33), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n488), .A2(KEYINPUT68), .A3(new_n489), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n494), .B1(new_n506), .B2(new_n495), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n493), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n486), .A2(new_n487), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n484), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n484), .B2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n515), .A3(new_n484), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n511), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n511), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n508), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n519), .B(new_n493), .C1(new_n507), .C2(new_n503), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n359), .A2(new_n483), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n421), .A2(new_n527), .A3(new_n428), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n421), .B2(new_n428), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT90), .B1(new_n474), .B2(new_n475), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532));
  AOI211_X1 g331(.A(new_n532), .B(new_n433), .C1(new_n465), .C2(new_n472), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n473), .B1(new_n534), .B2(new_n481), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n526), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n429), .A2(KEYINPUT87), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n421), .A2(new_n527), .A3(new_n428), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n531), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n474), .A2(KEYINPUT90), .A3(new_n475), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n481), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n473), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n545), .A3(KEYINPUT91), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n537), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n359), .A2(new_n523), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n525), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT37), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n425), .B2(new_n426), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n423), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT38), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n535), .A2(new_n418), .A3(new_n420), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT39), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n452), .B1(new_n461), .B2(new_n464), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n454), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n559), .B1(new_n558), .B2(new_n454), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n467), .A2(KEYINPUT89), .A3(new_n454), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n557), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT89), .B1(new_n467), .B2(new_n454), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n568), .A3(new_n560), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n569), .A3(new_n433), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n563), .A2(new_n569), .A3(KEYINPUT40), .A4(new_n433), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n538), .A2(new_n534), .A3(new_n539), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n556), .B(new_n359), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n521), .A2(KEYINPUT36), .A3(new_n522), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT36), .B1(new_n521), .B2(new_n522), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n359), .A2(new_n483), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n262), .B1(new_n549), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  OAI211_X1 g385(.A(KEYINPUT106), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G99gat), .ZN(new_n588));
  INV_X1    g387(.A(G106gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT8), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n586), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n584), .A2(KEYINPUT106), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n584), .A2(KEYINPUT106), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n593), .A2(G85gat), .A3(G92gat), .A4(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT107), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n592), .B(new_n595), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n596), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n598), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G71gat), .ZN(new_n602));
  INV_X1    g401(.A(G78gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(KEYINPUT100), .ZN(new_n607));
  INV_X1    g406(.A(G57gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G64gat), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G57gat), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n606), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n607), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n601), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n614), .B(KEYINPUT108), .C1(new_n601), .C2(new_n616), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n616), .A2(new_n601), .A3(KEYINPUT108), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT10), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n601), .A3(KEYINPUT10), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n583), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n617), .A2(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(new_n583), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n622), .A2(new_n625), .A3(new_n629), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT109), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT109), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n626), .A2(new_n634), .A3(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n613), .B(KEYINPUT101), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n233), .B1(KEYINPUT21), .B2(new_n616), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n645), .A2(new_n653), .A3(new_n648), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n655), .B2(new_n658), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n638), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n656), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n637), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(G134gat), .B(G162gat), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n240), .B2(KEYINPUT95), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n601), .B1(new_n671), .B2(new_n228), .ZN(new_n672));
  AND2_X1   g471(.A1(G232gat), .A2(G233gat), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n601), .A2(new_n226), .B1(KEYINPUT41), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G190gat), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n601), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n229), .B2(new_n230), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n373), .A3(new_n674), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n669), .B1(new_n680), .B2(new_n303), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n673), .A2(KEYINPUT41), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n676), .A2(new_n679), .A3(G218gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n681), .B2(new_n684), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n668), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n684), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n682), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n667), .A3(new_n685), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n582), .A2(new_n636), .A3(new_n666), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n480), .A2(new_n482), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n204), .ZN(G1324gat));
  XOR2_X1   g495(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n697));
  NOR2_X1   g496(.A1(new_n693), .A2(new_n540), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT111), .Z(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n702), .B(new_n703), .C1(new_n208), .C2(new_n698), .ZN(G1325gat));
  OAI21_X1  g503(.A(G15gat), .B1(new_n693), .B2(new_n579), .ZN(new_n705));
  INV_X1    g504(.A(new_n523), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n693), .B2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n359), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n549), .A2(new_n712), .A3(new_n581), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n549), .B2(new_n581), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n688), .A2(new_n691), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n713), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n692), .B1(new_n549), .B2(new_n581), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n716), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n661), .A2(new_n665), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n636), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n262), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n694), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n719), .A2(new_n724), .ZN(new_n727));
  INV_X1    g526(.A(new_n694), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n218), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1328gat));
  OAI21_X1  g530(.A(G36gat), .B1(new_n725), .B2(new_n540), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n219), .A3(new_n530), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT46), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1329gat));
  INV_X1    g534(.A(new_n579), .ZN(new_n736));
  AND4_X1   g535(.A1(G43gat), .A2(new_n721), .A3(new_n736), .A4(new_n724), .ZN(new_n737));
  AOI21_X1  g536(.A(G43gat), .B1(new_n727), .B2(new_n523), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1330gat));
  NOR3_X1   g540(.A1(new_n723), .A2(G50gat), .A3(new_n692), .ZN(new_n742));
  INV_X1    g541(.A(new_n359), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n582), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n725), .A2(new_n359), .ZN(new_n745));
  INV_X1    g544(.A(G50gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(KEYINPUT48), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1331gat));
  NAND3_X1  g550(.A1(new_n692), .A2(new_n262), .A3(new_n666), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n713), .A2(new_n714), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n636), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n694), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n608), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n540), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n755), .B2(new_n579), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n706), .A2(new_n636), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n753), .A2(new_n602), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g566(.A1(new_n755), .A2(new_n359), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n603), .ZN(G1335gat));
  NAND2_X1  g568(.A1(new_n722), .A2(new_n262), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n549), .A2(new_n581), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT113), .B1(new_n774), .B2(new_n715), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776));
  AOI211_X1 g575(.A(new_n776), .B(new_n692), .C1(new_n549), .C2(new_n581), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n771), .A2(new_n772), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n779), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(new_n773), .C1(new_n775), .C2(new_n777), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(new_n585), .A3(new_n728), .A4(new_n754), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n770), .A2(new_n636), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n721), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n694), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1336gat));
  OAI21_X1  g587(.A(G92gat), .B1(new_n786), .B2(new_n540), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n636), .A2(G92gat), .A3(new_n540), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT115), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g593(.A1(new_n783), .A2(new_n588), .A3(new_n764), .ZN(new_n795));
  OAI21_X1  g594(.A(G99gat), .B1(new_n786), .B2(new_n579), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1338gat));
  OAI211_X1 g596(.A(new_n743), .B(new_n785), .C1(new_n718), .C2(new_n720), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n798), .B2(G106gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n636), .A2(new_n359), .A3(G106gat), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n780), .A2(KEYINPUT117), .A3(new_n782), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n782), .A3(new_n800), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT118), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  AND4_X1   g605(.A1(KEYINPUT118), .A2(new_n805), .A3(new_n801), .A4(new_n799), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n798), .A2(G106gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(KEYINPUT53), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n810), .A2(new_n808), .A3(KEYINPUT53), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n806), .A2(new_n807), .B1(new_n811), .B2(new_n812), .ZN(G1339gat));
  AOI21_X1  g612(.A(new_n245), .B1(new_n242), .B2(new_n243), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n232), .B1(new_n231), .B2(new_n234), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n254), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n259), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n633), .A2(new_n635), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n624), .B(new_n620), .C1(new_n623), .C2(KEYINPUT10), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n622), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n822), .B(new_n583), .C1(new_n619), .C2(new_n621), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n630), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n824), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n622), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n632), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n818), .B1(new_n829), .B2(new_n262), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n692), .ZN(new_n831));
  INV_X1    g630(.A(new_n829), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n715), .A2(new_n832), .A3(new_n817), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n666), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n692), .A2(new_n666), .A3(new_n262), .A4(new_n636), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n694), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n548), .A2(new_n530), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n262), .ZN(new_n842));
  AOI21_X1  g641(.A(G113gat), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n837), .A2(new_n743), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n694), .A2(new_n530), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n706), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n262), .A2(new_n437), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  AOI21_X1  g648(.A(G120gat), .B1(new_n841), .B2(new_n754), .ZN(new_n850));
  INV_X1    g649(.A(new_n846), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n706), .A2(new_n636), .A3(new_n435), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(G1341gat));
  NAND3_X1  g652(.A1(new_n841), .A2(new_n443), .A3(new_n666), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n846), .A2(new_n706), .A3(new_n722), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n443), .ZN(G1342gat));
  NOR3_X1   g655(.A1(new_n840), .A2(G134gat), .A3(new_n692), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT56), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n846), .A2(new_n706), .A3(new_n692), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n441), .B2(new_n859), .ZN(G1343gat));
  NOR3_X1   g659(.A1(new_n736), .A2(new_n359), .A3(new_n530), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n838), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n270), .B1(new_n862), .B2(new_n262), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n579), .A2(new_n845), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n837), .A2(new_n359), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n828), .A2(new_n632), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT55), .B1(new_n826), .B2(new_n827), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n825), .A2(KEYINPUT119), .A3(new_n828), .A4(new_n632), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n842), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n715), .B1(new_n873), .B2(new_n818), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n825), .A2(new_n632), .A3(new_n828), .A4(new_n817), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n688), .B2(new_n691), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n722), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n836), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n359), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n867), .B1(new_n881), .B2(new_n866), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n842), .A2(G141gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n863), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n884), .B(new_n885), .ZN(G1344gat));
  OAI211_X1 g685(.A(KEYINPUT57), .B(new_n743), .C1(new_n834), .C2(new_n836), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n876), .B1(new_n692), .B2(new_n830), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n835), .B1(new_n889), .B2(new_n666), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT57), .A4(new_n743), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n359), .B1(new_n877), .B2(new_n835), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n888), .B(new_n892), .C1(new_n893), .C2(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n864), .A2(new_n636), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(KEYINPUT122), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G148gat), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT122), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n268), .A2(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n882), .B2(new_n636), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n862), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n268), .A3(new_n754), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1345gat));
  AOI21_X1  g704(.A(G155gat), .B1(new_n903), .B2(new_n666), .ZN(new_n906));
  INV_X1    g705(.A(new_n882), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n666), .A2(G155gat), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT123), .Z(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n907), .B2(new_n909), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n903), .B2(new_n715), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n715), .A2(G162gat), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n907), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n837), .A2(new_n728), .ZN(new_n914));
  INV_X1    g713(.A(new_n548), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(new_n530), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n364), .A3(new_n842), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n694), .A2(new_n530), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n706), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n844), .A2(new_n842), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n922), .B2(G169gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n917), .A2(new_n919), .A3(new_n364), .A4(new_n842), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1348gat));
  NAND2_X1  g725(.A1(new_n844), .A2(new_n921), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n365), .A3(new_n636), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n917), .A2(new_n754), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n365), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n927), .B2(new_n722), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n666), .A2(new_n392), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n916), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n391), .A3(new_n715), .ZN(new_n935));
  OAI21_X1  g734(.A(G190gat), .B1(new_n927), .B2(new_n692), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1351gat));
  NAND3_X1  g737(.A1(new_n579), .A2(new_n743), .A3(new_n530), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT126), .Z(new_n940));
  NAND2_X1  g739(.A1(new_n914), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n842), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n736), .A2(new_n920), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n894), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n842), .A2(G197gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n636), .A2(G204gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n942), .B2(new_n950), .ZN(new_n951));
  NOR4_X1   g750(.A1(new_n941), .A2(KEYINPUT62), .A3(G204gat), .A4(new_n636), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n945), .B2(new_n636), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n302), .A3(new_n666), .ZN(new_n960));
  OAI21_X1  g759(.A(G211gat), .B1(new_n945), .B2(new_n722), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n945), .B2(new_n692), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n942), .A2(new_n303), .A3(new_n715), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


