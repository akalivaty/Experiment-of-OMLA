//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  INV_X1    g032(.A(new_n451), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(G2106), .B2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(new_n460), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n467), .B1(new_n464), .B2(new_n465), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G124), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AOI21_X1  g060(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(G138), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n467), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n487), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT68), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n494), .A2(new_n501), .A3(new_n505), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(new_n516), .A3(G62), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n520), .A2(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n518), .A2(new_n528), .ZN(G166));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n525), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n510), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n531), .A2(G51), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(new_n513), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n511), .B2(new_n512), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT72), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n523), .A2(new_n522), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n547), .B(new_n544), .C1(new_n548), .C2(new_n542), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n546), .A2(new_n549), .A3(new_n552), .A4(G651), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n520), .A2(new_n554), .B1(new_n526), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  XNOR2_X1  g135(.A(KEYINPUT75), .B(G81), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n520), .A2(new_n560), .B1(new_n526), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n548), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n508), .B1(new_n565), .B2(new_n566), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  AOI22_X1  g149(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n508), .B1(new_n576), .B2(new_n526), .ZN(new_n577));
  OAI211_X1 g152(.A(G53), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n526), .B2(new_n585), .C1(new_n586), .C2(new_n520), .ZN(G288));
  AOI22_X1  g162(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n508), .ZN(new_n589));
  INV_X1    g164(.A(G48), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n520), .A2(new_n590), .B1(new_n526), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n508), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n520), .A2(new_n597), .B1(new_n526), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n548), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n531), .B2(G54), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n526), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n513), .A2(new_n519), .A3(KEYINPUT10), .A4(G92), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G321));
  XOR2_X1   g189(.A(G321), .B(KEYINPUT76), .Z(G284));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n581), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NOR2_X1   g196(.A1(new_n569), .A2(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(G111), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G2105), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n477), .A2(G135), .ZN(new_n630));
  AOI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G123), .C2(new_n482), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT78), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n466), .A2(new_n461), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT79), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT80), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(new_n659), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT81), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n660), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n659), .A2(new_n662), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n658), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  AND2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT83), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n676), .A2(new_n683), .A3(new_n679), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT84), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  NAND2_X1  g269(.A1(new_n593), .A2(G16), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n696));
  OR2_X1    g271(.A1(G6), .A2(G16), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n700));
  OAI21_X1  g275(.A(G1981), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n703), .A3(new_n698), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(G16), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G1971), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n708), .A2(G1971), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n709), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n706), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n719), .A2(new_n720), .A3(new_n705), .A4(new_n709), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(KEYINPUT34), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n718), .A2(KEYINPUT86), .A3(KEYINPUT34), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(KEYINPUT34), .B1(new_n718), .B2(new_n721), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n477), .A2(G131), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(G107), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G119), .B2(new_n482), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G25), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n710), .A2(G24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n600), .B2(new_n710), .ZN(new_n741));
  INV_X1    g316(.A(G1986), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n727), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n726), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n726), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G26), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT87), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n477), .A2(G140), .ZN(new_n756));
  OAI21_X1  g331(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n757));
  INV_X1    g332(.A(G116), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G2105), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G128), .B2(new_n482), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n755), .B1(new_n762), .B2(new_n751), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT88), .B(G2067), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n710), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n581), .B2(new_n710), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n763), .A2(new_n765), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n710), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n619), .B2(new_n710), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n751), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n751), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT29), .B(G2090), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n763), .A2(new_n765), .B1(new_n766), .B2(new_n770), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT24), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G160), .B2(new_n751), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G19), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n569), .B2(G16), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(G1348), .B2(new_n773), .C1(new_n789), .C2(G1341), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n775), .A2(new_n779), .A3(new_n780), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n751), .A2(G27), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n751), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(G2078), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n477), .A2(G139), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT90), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n466), .A2(G127), .ZN(new_n800));
  AND2_X1   g375(.A1(G115), .A2(G2104), .ZN(new_n801));
  OAI21_X1  g376(.A(G2105), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n795), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G33), .B(new_n803), .S(G29), .Z(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G2072), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n804), .A2(G2072), .B1(G1341), .B2(new_n789), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n751), .A2(G32), .ZN(new_n807));
  NAND3_X1  g382(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT26), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n482), .A2(G129), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n461), .A2(G105), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n477), .B2(G141), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n751), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT27), .B(G1996), .Z(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  AND4_X1   g391(.A1(new_n794), .A2(new_n805), .A3(new_n806), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G171), .A2(new_n710), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G5), .B2(new_n710), .ZN(new_n819));
  INV_X1    g394(.A(G1961), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(G2078), .B2(new_n793), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n791), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n710), .A2(G21), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G168), .B2(new_n710), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(G1966), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n631), .A2(G29), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(G1966), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT30), .B(G28), .ZN(new_n830));
  OR2_X1    g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  NAND2_X1  g406(.A1(KEYINPUT31), .A2(G11), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n830), .A2(new_n751), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND4_X1   g408(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n824), .A2(KEYINPUT92), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT92), .B1(new_n824), .B2(new_n834), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n822), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(KEYINPUT93), .B1(new_n750), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n726), .A2(new_n745), .A3(new_n748), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n748), .B1(new_n726), .B2(new_n745), .ZN(new_n840));
  OAI211_X1 g415(.A(KEYINPUT93), .B(new_n837), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n838), .A2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n750), .A2(new_n837), .ZN(G150));
  NAND2_X1  g419(.A1(new_n619), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n508), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  INV_X1    g424(.A(G93), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n520), .A2(new_n849), .B1(new_n526), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n569), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n569), .B(new_n848), .C1(new_n853), .C2(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n846), .B(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n862), .A2(new_n863), .A3(G860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n855), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(G160), .B(KEYINPUT95), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n484), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n631), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n482), .A2(G130), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT97), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(G118), .B2(new_n467), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(KEYINPUT97), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n477), .B2(G142), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(new_n635), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n733), .ZN(new_n880));
  INV_X1    g455(.A(new_n813), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n803), .A2(KEYINPUT96), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n499), .B1(new_n493), .B2(new_n488), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n499), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n494), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n803), .A2(KEYINPUT96), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n761), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n761), .B1(new_n884), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n881), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n888), .A3(new_n813), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n880), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n893), .A3(new_n880), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n897), .B2(KEYINPUT98), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n871), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n897), .A2(new_n894), .A3(new_n870), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(G37), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT40), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G395));
  NAND2_X1  g482(.A1(new_n855), .A2(new_n612), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(new_n593), .ZN(new_n909));
  NAND2_X1  g484(.A1(G290), .A2(G288), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n712), .A2(new_n600), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT101), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n915), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n915), .B2(new_n917), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n919), .B1(new_n924), .B2(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n859), .B(new_n623), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT99), .B1(new_n581), .B2(new_n611), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n610), .B(new_n605), .C1(new_n577), .C2(new_n580), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n581), .A2(KEYINPUT99), .A3(new_n611), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT41), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n928), .A2(new_n935), .A3(new_n929), .A4(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n932), .B(KEYINPUT100), .C1(new_n926), .C2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(KEYINPUT100), .B2(new_n932), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n925), .B(new_n939), .Z(new_n940));
  OAI21_X1  g515(.A(new_n908), .B1(new_n940), .B2(new_n612), .ZN(G295));
  OAI21_X1  g516(.A(new_n908), .B1(new_n940), .B2(new_n612), .ZN(G331));
  NAND2_X1  g517(.A1(G301), .A2(G168), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT103), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n945));
  NAND3_X1  g520(.A1(G301), .A2(new_n945), .A3(G168), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n551), .A2(G286), .A3(new_n553), .A4(new_n557), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT104), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n556), .B1(new_n550), .B2(KEYINPUT73), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(G286), .A4(new_n553), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n859), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n945), .B1(G301), .B2(G168), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT103), .B(G286), .C1(new_n950), .C2(new_n553), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n953), .B(new_n859), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n959), .A2(new_n931), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n944), .A2(new_n946), .B1(new_n949), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT106), .B1(new_n961), .B2(new_n859), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n958), .A2(new_n957), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n949), .A2(new_n952), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n860), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n959), .ZN(new_n968));
  INV_X1    g543(.A(new_n937), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI211_X1 g545(.A(KEYINPUT105), .B(new_n937), .C1(new_n967), .C2(new_n959), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n923), .B(new_n963), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n974), .B2(new_n924), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n959), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n969), .B1(new_n978), .B2(new_n954), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n968), .A2(new_n964), .A3(new_n969), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n923), .B1(new_n982), .B2(new_n963), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT107), .B1(new_n983), .B2(G37), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n956), .A2(new_n962), .A3(new_n959), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n969), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n960), .A2(new_n967), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT108), .A3(new_n924), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n986), .A2(new_n969), .B1(new_n967), .B2(new_n960), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(new_n923), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G37), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n972), .A2(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n994), .A2(KEYINPUT43), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT44), .B1(new_n985), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n977), .B2(new_n984), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n994), .A2(new_n1000), .A3(new_n996), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(G397));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n883), .B2(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G160), .A2(G40), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n761), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n881), .A2(G1996), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1008), .A2(G1996), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT110), .Z(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1014), .B2(new_n813), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1008), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n734), .A2(new_n737), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n734), .A2(new_n737), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1008), .A2(new_n742), .A3(new_n600), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1008), .A2(G1986), .A3(G290), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT109), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n504), .A2(new_n1028), .A3(new_n506), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1005), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n883), .A2(G1384), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1007), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1027), .B1(new_n1033), .B2(G2078), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT123), .B(new_n1027), .C1(new_n1033), .C2(G2078), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT122), .B(G1961), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n886), .A2(new_n1040), .A3(new_n1028), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT111), .B1(new_n883), .B2(G1384), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n471), .A2(new_n472), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G2105), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n486), .A2(G137), .B1(G101), .B2(new_n461), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1046), .A2(G40), .A3(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1039), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1027), .B(G2078), .C1(new_n1031), .C2(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(KEYINPUT124), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n1046), .A3(G40), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1047), .A2(KEYINPUT124), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(KEYINPUT125), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(KEYINPUT125), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(new_n1006), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1051), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1038), .A2(new_n1060), .A3(G301), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1005), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1028), .A4(new_n506), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1048), .A3(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1066), .A2(new_n1027), .A3(G2078), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(new_n1051), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1038), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1026), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1038), .A2(new_n1068), .A3(G301), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1038), .A2(new_n1060), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1071), .B(KEYINPUT54), .C1(new_n1072), .C2(G301), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1041), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1075), .B(new_n1077), .C1(new_n1076), .C2(G288), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1074), .B(G8), .C1(new_n1076), .C2(G288), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT52), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n593), .A2(new_n703), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n589), .A2(new_n592), .A3(G1981), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT112), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT112), .B(new_n1085), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1075), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1078), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G166), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT55), .ZN(new_n1091));
  INV_X1    g666(.A(G1971), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1033), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G2090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1049), .A2(new_n1094), .A3(new_n1050), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1089), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1088), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1007), .B1(new_n1063), .B2(KEYINPUT50), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n504), .A2(new_n1043), .A3(new_n1028), .A4(new_n506), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1098), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1971), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1101));
  OAI21_X1  g676(.A(G8), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1091), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1066), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1050), .A2(new_n786), .A3(new_n1048), .A4(new_n1044), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1089), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G168), .A2(new_n1089), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT120), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(KEYINPUT51), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1109), .B2(KEYINPUT121), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1115), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1110), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1070), .A2(new_n1073), .A3(new_n1105), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1122));
  INV_X1    g697(.A(G1996), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1030), .A2(new_n1123), .A3(new_n1032), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1074), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n569), .B(new_n1122), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n581), .B(KEYINPUT57), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1030), .A2(new_n1032), .A3(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1132), .B(new_n1134), .C1(new_n1135), .C2(G1956), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1134), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1956), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(KEYINPUT61), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1130), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1124), .A2(new_n1125), .B1(new_n1074), .B2(new_n1127), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n856), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1145));
  OAI211_X1 g720(.A(new_n1131), .B(new_n1141), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT117), .B(KEYINPUT61), .Z(new_n1147));
  INV_X1    g722(.A(new_n1136), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1140), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(KEYINPUT118), .B(new_n1147), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1146), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1348), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1074), .A2(G2067), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT114), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1348), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT114), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1157), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1155), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(KEYINPUT119), .A3(new_n611), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n619), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1154), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1169), .A2(new_n1148), .A3(new_n611), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(new_n1149), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1120), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1117), .A2(new_n1180), .A3(new_n1118), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1069), .A2(new_n1104), .A3(new_n1097), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT113), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1089), .B(G286), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1186), .A2(G8), .A3(new_n1091), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1078), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1104), .A2(new_n1185), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1109), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1096), .A2(new_n1091), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1097), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(G288), .A2(G1976), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1087), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1082), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1075), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(new_n1187), .B2(new_n1088), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1184), .B1(new_n1195), .B2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g778(.A(KEYINPUT113), .B(new_n1201), .C1(new_n1191), .C2(new_n1194), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1183), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1025), .B1(new_n1178), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1015), .A2(new_n1017), .B1(new_n1009), .B2(new_n762), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1207), .A2(new_n1008), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT126), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1022), .B(KEYINPUT48), .Z(new_n1210));
  NAND2_X1  g785(.A1(new_n1020), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1010), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1016), .B1(new_n1212), .B2(new_n881), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1014), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1209), .A2(new_n1211), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1206), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g796(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1223));
  NAND3_X1  g797(.A1(new_n673), .A2(G319), .A3(new_n654), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1224), .A2(G229), .ZN(new_n1225));
  INV_X1    g799(.A(new_n904), .ZN(new_n1226));
  OAI21_X1  g800(.A(new_n1225), .B1(new_n1226), .B2(new_n901), .ZN(new_n1227));
  NOR2_X1   g801(.A1(new_n1223), .A2(new_n1227), .ZN(G308));
  OAI221_X1 g802(.A(new_n1225), .B1(new_n1226), .B2(new_n901), .C1(new_n1001), .C2(new_n1002), .ZN(G225));
endmodule


