// Benchmark "locked_c3540" written by ABC on Sat Dec 16 11:14:50 2023

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41,
    G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132,
    G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226,
    G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311,
    G317, G322, G326, G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13,
    G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124,
    G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213,
    G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283,
    G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137, new_n138, new_n139, new_n140, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n174, new_n175,
    new_n176, new_n177, new_n178, new_n179, new_n180, new_n181, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n192, new_n193, new_n194, new_n195, new_n196, new_n197,
    new_n198, new_n199, new_n200, new_n201, new_n202, new_n203, new_n204,
    new_n205, new_n206, new_n207, new_n208, new_n209, new_n210, new_n211,
    new_n212, new_n213, new_n214, new_n215, new_n216, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223, new_n224, new_n225,
    new_n226, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023;
  INV_X1    g000(.A(G50), .ZN(new_n137));
  INV_X1    g001(.A(G58), .ZN(new_n138));
  INV_X1    g002(.A(G68), .ZN(new_n139));
  NAND3_X1  g003(.A1(new_n137), .A2(new_n138), .A3(new_n139), .ZN(new_n140));
  NOR2_X1   g004(.A1(new_n140), .A2(G77), .ZN(G353));
  OAI21_X1  g005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n143));
  INV_X1    g007(.A(G20), .ZN(new_n144));
  NAND2_X1  g008(.A1(G1), .A2(G13), .ZN(new_n145));
  NOR3_X1   g009(.A1(new_n143), .A2(new_n144), .A3(new_n145), .ZN(new_n146));
  INV_X1    g010(.A(G1), .ZN(new_n147));
  NOR3_X1   g011(.A1(new_n147), .A2(new_n144), .A3(G13), .ZN(new_n148));
  OAI211_X1 g012(.A(new_n148), .B(G250), .C1(G257), .C2(G264), .ZN(new_n149));
  XNOR2_X1  g013(.A(new_n149), .B(KEYINPUT0), .ZN(new_n150));
  AOI22_X1  g014(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n151));
  NAND2_X1  g015(.A1(G87), .A2(G250), .ZN(new_n152));
  NAND2_X1  g016(.A1(G116), .A2(G270), .ZN(new_n153));
  NAND3_X1  g017(.A1(new_n151), .A2(new_n152), .A3(new_n153), .ZN(new_n154));
  AOI21_X1  g018(.A(new_n154), .B1(G50), .B2(G226), .ZN(new_n155));
  INV_X1    g019(.A(G232), .ZN(new_n156));
  INV_X1    g020(.A(G107), .ZN(new_n157));
  INV_X1    g021(.A(G264), .ZN(new_n158));
  OAI221_X1 g022(.A(new_n155), .B1(new_n138), .B2(new_n156), .C1(new_n157), .C2(new_n158), .ZN(new_n159));
  AND2_X1   g023(.A1(G77), .A2(G244), .ZN(new_n160));
  OAI22_X1  g024(.A1(new_n159), .A2(new_n160), .B1(new_n147), .B2(new_n144), .ZN(new_n161));
  OAI21_X1  g025(.A(new_n150), .B1(new_n161), .B2(KEYINPUT1), .ZN(new_n162));
  AOI211_X1 g026(.A(new_n146), .B(new_n162), .C1(KEYINPUT1), .C2(new_n161), .ZN(G361));
  XNOR2_X1  g027(.A(G238), .B(G244), .ZN(new_n164));
  XNOR2_X1  g028(.A(new_n164), .B(KEYINPUT2), .ZN(new_n165));
  INV_X1    g029(.A(G226), .ZN(new_n166));
  XNOR2_X1  g030(.A(new_n165), .B(new_n166), .ZN(new_n167));
  XNOR2_X1  g031(.A(new_n167), .B(new_n156), .ZN(new_n168));
  XNOR2_X1  g032(.A(G264), .B(G270), .ZN(new_n169));
  XNOR2_X1  g033(.A(new_n169), .B(G250), .ZN(new_n170));
  INV_X1    g034(.A(G257), .ZN(new_n171));
  XNOR2_X1  g035(.A(new_n170), .B(new_n171), .ZN(new_n172));
  XNOR2_X1  g036(.A(new_n168), .B(new_n172), .ZN(G358));
  XNOR2_X1  g037(.A(G87), .B(G97), .ZN(new_n174));
  XNOR2_X1  g038(.A(new_n174), .B(new_n157), .ZN(new_n175));
  INV_X1    g039(.A(G116), .ZN(new_n176));
  XNOR2_X1  g040(.A(new_n175), .B(new_n176), .ZN(new_n177));
  XNOR2_X1  g041(.A(G58), .B(G68), .ZN(new_n178));
  XNOR2_X1  g042(.A(new_n178), .B(G50), .ZN(new_n179));
  INV_X1    g043(.A(G77), .ZN(new_n180));
  XNOR2_X1  g044(.A(new_n179), .B(new_n180), .ZN(new_n181));
  XOR2_X1   g045(.A(new_n177), .B(new_n181), .Z(G351));
  INV_X1    g046(.A(G33), .ZN(new_n183));
  NAND2_X1  g047(.A1(new_n183), .A2(KEYINPUT3), .ZN(new_n184));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n185));
  NAND2_X1  g049(.A1(new_n185), .A2(G33), .ZN(new_n186));
  NAND2_X1  g050(.A1(new_n184), .A2(new_n186), .ZN(new_n187));
  AOI21_X1  g051(.A(KEYINPUT7), .B1(new_n187), .B2(new_n144), .ZN(new_n188));
  INV_X1    g052(.A(KEYINPUT7), .ZN(new_n189));
  AOI211_X1 g053(.A(new_n189), .B(G20), .C1(new_n184), .C2(new_n186), .ZN(new_n190));
  OAI21_X1  g054(.A(G68), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  NOR2_X1   g055(.A1(G20), .A2(G33), .ZN(new_n192));
  NAND2_X1  g056(.A1(new_n192), .A2(G159), .ZN(new_n193));
  NAND2_X1  g057(.A1(new_n178), .A2(G20), .ZN(new_n194));
  NAND3_X1  g058(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g059(.A(KEYINPUT16), .ZN(new_n196));
  NAND2_X1  g060(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n198));
  NAND2_X1  g062(.A1(new_n198), .A2(new_n145), .ZN(new_n199));
  NAND4_X1  g063(.A1(new_n191), .A2(KEYINPUT16), .A3(new_n193), .A4(new_n194), .ZN(new_n200));
  NAND3_X1  g064(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g065(.A(KEYINPUT8), .B(G58), .ZN(new_n202));
  NAND3_X1  g066(.A1(new_n147), .A2(G13), .A3(G20), .ZN(new_n203));
  INV_X1    g067(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g068(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g069(.A(new_n199), .B1(new_n147), .B2(G20), .ZN(new_n206));
  INV_X1    g070(.A(new_n202), .ZN(new_n207));
  NAND2_X1  g071(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g072(.A1(new_n201), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g073(.A(new_n145), .ZN(new_n210));
  NAND2_X1  g074(.A1(G33), .A2(G41), .ZN(new_n211));
  NAND2_X1  g075(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g076(.A(new_n147), .B1(G41), .B2(G45), .ZN(new_n213));
  NAND2_X1  g077(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g078(.A(G274), .ZN(new_n215));
  OAI22_X1  g079(.A1(new_n214), .A2(new_n156), .B1(new_n215), .B2(new_n213), .ZN(new_n216));
  XNOR2_X1  g080(.A(KEYINPUT3), .B(G33), .ZN(new_n217));
  INV_X1    g081(.A(G1698), .ZN(new_n218));
  NAND3_X1  g082(.A1(new_n217), .A2(G223), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g083(.A1(G33), .A2(G87), .ZN(new_n220));
  NAND2_X1  g084(.A1(new_n217), .A2(G1698), .ZN(new_n221));
  OAI211_X1 g085(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n166), .ZN(new_n222));
  INV_X1    g086(.A(new_n212), .ZN(new_n223));
  AOI21_X1  g087(.A(new_n216), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g088(.A1(new_n224), .A2(G179), .ZN(new_n225));
  INV_X1    g089(.A(G169), .ZN(new_n226));
  OAI21_X1  g090(.A(new_n225), .B1(new_n226), .B2(new_n224), .ZN(new_n227));
  NAND2_X1  g091(.A1(new_n209), .A2(new_n227), .ZN(new_n228));
  INV_X1    g092(.A(KEYINPUT18), .ZN(new_n229));
  NAND2_X1  g093(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g094(.A1(new_n209), .A2(KEYINPUT18), .A3(new_n227), .ZN(new_n231));
  NAND2_X1  g095(.A1(new_n222), .A2(new_n223), .ZN(new_n232));
  INV_X1    g096(.A(G190), .ZN(new_n233));
  INV_X1    g097(.A(new_n216), .ZN(new_n234));
  NAND3_X1  g098(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g099(.A(new_n235), .B1(G200), .B2(new_n224), .ZN(new_n236));
  NAND4_X1  g100(.A1(new_n201), .A2(new_n236), .A3(new_n205), .A4(new_n208), .ZN(new_n237));
  OR2_X1    g101(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g102(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n239));
  AOI22_X1  g103(.A1(new_n230), .A2(new_n231), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI22_X1  g104(.A1(new_n140), .A2(G20), .B1(G150), .B2(new_n192), .ZN(new_n241));
  NAND2_X1  g105(.A1(new_n144), .A2(G33), .ZN(new_n242));
  OAI21_X1  g106(.A(new_n241), .B1(new_n242), .B2(new_n202), .ZN(new_n243));
  NAND2_X1  g107(.A1(new_n243), .A2(new_n199), .ZN(new_n244));
  NAND2_X1  g108(.A1(new_n204), .A2(new_n137), .ZN(new_n245));
  NAND2_X1  g109(.A1(new_n206), .A2(G50), .ZN(new_n246));
  NAND3_X1  g110(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g111(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g112(.A1(new_n213), .A2(new_n215), .ZN(new_n249));
  NAND3_X1  g113(.A1(new_n217), .A2(G222), .A3(new_n218), .ZN(new_n250));
  INV_X1    g114(.A(G223), .ZN(new_n251));
  OAI221_X1 g115(.A(new_n250), .B1(new_n180), .B2(new_n217), .C1(new_n221), .C2(new_n251), .ZN(new_n252));
  AOI21_X1  g116(.A(new_n249), .B1(new_n252), .B2(new_n223), .ZN(new_n253));
  OAI21_X1  g117(.A(new_n253), .B1(new_n166), .B2(new_n214), .ZN(new_n254));
  INV_X1    g118(.A(G179), .ZN(new_n255));
  OR2_X1    g119(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g120(.A1(new_n254), .A2(G169), .ZN(new_n257));
  AOI21_X1  g121(.A(new_n248), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g122(.A1(new_n254), .A2(new_n233), .ZN(new_n259));
  XNOR2_X1  g123(.A(new_n247), .B(KEYINPUT9), .ZN(new_n260));
  NAND2_X1  g124(.A1(new_n254), .A2(G200), .ZN(new_n261));
  NAND3_X1  g125(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g126(.A1(new_n262), .A2(KEYINPUT10), .ZN(new_n263));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n264));
  NAND4_X1  g128(.A1(new_n259), .A2(new_n264), .A3(new_n260), .A4(new_n261), .ZN(new_n265));
  AOI21_X1  g129(.A(new_n258), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g130(.A1(new_n240), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g131(.A1(new_n192), .A2(G50), .B1(G20), .B2(new_n139), .ZN(new_n268));
  OAI21_X1  g132(.A(new_n268), .B1(new_n180), .B2(new_n242), .ZN(new_n269));
  NAND2_X1  g133(.A1(new_n269), .A2(new_n199), .ZN(new_n270));
  XNOR2_X1  g134(.A(new_n270), .B(KEYINPUT11), .ZN(new_n271));
  NAND2_X1  g135(.A1(new_n204), .A2(new_n139), .ZN(new_n272));
  XNOR2_X1  g136(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  INV_X1    g137(.A(new_n206), .ZN(new_n274));
  OAI211_X1 g138(.A(new_n271), .B(new_n273), .C1(new_n139), .C2(new_n274), .ZN(new_n275));
  INV_X1    g139(.A(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g140(.A1(new_n217), .A2(G226), .A3(new_n218), .ZN(new_n277));
  NAND2_X1  g141(.A1(G33), .A2(G97), .ZN(new_n278));
  OAI211_X1 g142(.A(new_n277), .B(new_n278), .C1(new_n221), .C2(new_n156), .ZN(new_n279));
  AOI21_X1  g143(.A(new_n249), .B1(new_n279), .B2(new_n223), .ZN(new_n280));
  INV_X1    g144(.A(new_n214), .ZN(new_n281));
  NAND2_X1  g145(.A1(new_n281), .A2(G238), .ZN(new_n282));
  AOI21_X1  g146(.A(new_n276), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g147(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g148(.A1(new_n280), .A2(new_n276), .A3(new_n282), .ZN(new_n285));
  NAND2_X1  g149(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g150(.A(G200), .ZN(new_n287));
  NAND2_X1  g151(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g152(.A1(new_n284), .A2(new_n233), .A3(new_n285), .ZN(new_n289));
  AOI21_X1  g153(.A(new_n275), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g154(.A(new_n285), .ZN(new_n291));
  OAI21_X1  g155(.A(G169), .B1(new_n291), .B2(new_n283), .ZN(new_n292));
  NAND2_X1  g156(.A1(new_n292), .A2(KEYINPUT14), .ZN(new_n293));
  INV_X1    g157(.A(KEYINPUT14), .ZN(new_n294));
  NAND3_X1  g158(.A1(new_n286), .A2(new_n294), .A3(G169), .ZN(new_n295));
  NAND3_X1  g159(.A1(new_n284), .A2(G179), .A3(new_n285), .ZN(new_n296));
  NAND3_X1  g160(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g161(.A(new_n290), .B1(new_n297), .B2(new_n275), .ZN(new_n298));
  AOI22_X1  g162(.A1(new_n207), .A2(new_n192), .B1(G20), .B2(G77), .ZN(new_n299));
  XNOR2_X1  g163(.A(KEYINPUT15), .B(G87), .ZN(new_n300));
  OAI21_X1  g164(.A(new_n299), .B1(new_n242), .B2(new_n300), .ZN(new_n301));
  AOI22_X1  g165(.A1(new_n301), .A2(new_n199), .B1(G77), .B2(new_n206), .ZN(new_n302));
  NAND2_X1  g166(.A1(new_n204), .A2(new_n180), .ZN(new_n303));
  NAND2_X1  g167(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g168(.A1(new_n217), .A2(G232), .A3(new_n218), .ZN(new_n305));
  INV_X1    g169(.A(G238), .ZN(new_n306));
  OAI221_X1 g170(.A(new_n305), .B1(new_n157), .B2(new_n217), .C1(new_n221), .C2(new_n306), .ZN(new_n307));
  AOI21_X1  g171(.A(new_n249), .B1(new_n307), .B2(new_n223), .ZN(new_n308));
  NAND2_X1  g172(.A1(new_n281), .A2(G244), .ZN(new_n309));
  NAND2_X1  g173(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g174(.A1(new_n310), .A2(new_n255), .ZN(new_n311));
  AOI21_X1  g175(.A(new_n226), .B1(new_n308), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g176(.A(new_n304), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g177(.A(new_n304), .ZN(new_n314));
  NOR2_X1   g178(.A1(new_n310), .A2(G190), .ZN(new_n315));
  AOI21_X1  g179(.A(G200), .B1(new_n308), .B2(new_n309), .ZN(new_n316));
  OAI21_X1  g180(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g181(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g182(.A1(new_n267), .A2(new_n298), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g183(.A(KEYINPUT5), .B(G41), .ZN(new_n320));
  NAND3_X1  g184(.A1(new_n147), .A2(G45), .A3(G274), .ZN(new_n321));
  INV_X1    g185(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g186(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g187(.A(G41), .ZN(new_n324));
  NAND2_X1  g188(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n325));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n326));
  NAND2_X1  g190(.A1(new_n326), .A2(G41), .ZN(new_n327));
  NAND2_X1  g191(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g192(.A1(new_n147), .A2(G45), .ZN(new_n329));
  OAI21_X1  g193(.A(new_n212), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g194(.A(new_n323), .B1(new_n330), .B2(new_n158), .ZN(new_n331));
  NAND3_X1  g195(.A1(new_n217), .A2(G250), .A3(new_n218), .ZN(new_n332));
  NAND2_X1  g196(.A1(G33), .A2(G294), .ZN(new_n333));
  OAI211_X1 g197(.A(new_n332), .B(new_n333), .C1(new_n221), .C2(new_n171), .ZN(new_n334));
  AOI21_X1  g198(.A(new_n331), .B1(new_n223), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g199(.A1(new_n335), .A2(G179), .ZN(new_n336));
  OAI21_X1  g200(.A(new_n336), .B1(new_n226), .B2(new_n335), .ZN(new_n337));
  NAND4_X1  g201(.A1(new_n184), .A2(new_n186), .A3(new_n144), .A4(G87), .ZN(new_n338));
  NAND2_X1  g202(.A1(new_n338), .A2(KEYINPUT22), .ZN(new_n339));
  INV_X1    g203(.A(KEYINPUT22), .ZN(new_n340));
  NAND4_X1  g204(.A1(new_n217), .A2(new_n340), .A3(new_n144), .A4(G87), .ZN(new_n341));
  NAND2_X1  g205(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g206(.A1(G33), .A2(G116), .ZN(new_n343));
  NOR2_X1   g207(.A1(new_n343), .A2(G20), .ZN(new_n344));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n345));
  OAI21_X1  g209(.A(new_n345), .B1(new_n144), .B2(G107), .ZN(new_n346));
  NAND3_X1  g210(.A1(new_n157), .A2(KEYINPUT23), .A3(G20), .ZN(new_n347));
  AOI21_X1  g211(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g212(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g213(.A(KEYINPUT24), .ZN(new_n350));
  NAND2_X1  g214(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g215(.A1(new_n342), .A2(KEYINPUT24), .A3(new_n348), .ZN(new_n352));
  NAND3_X1  g216(.A1(new_n351), .A2(new_n199), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g217(.A1(new_n203), .A2(G107), .ZN(new_n354));
  XNOR2_X1  g218(.A(new_n354), .B(KEYINPUT25), .ZN(new_n355));
  NAND2_X1  g219(.A1(new_n147), .A2(G33), .ZN(new_n356));
  NAND3_X1  g220(.A1(new_n356), .A2(new_n145), .A3(new_n198), .ZN(new_n357));
  NOR2_X1   g221(.A1(new_n357), .A2(new_n204), .ZN(new_n358));
  NAND2_X1  g222(.A1(new_n358), .A2(G107), .ZN(new_n359));
  NAND3_X1  g223(.A1(new_n353), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g224(.A1(new_n337), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g225(.A1(new_n334), .A2(new_n223), .ZN(new_n362));
  NOR2_X1   g226(.A1(new_n328), .A2(new_n321), .ZN(new_n363));
  INV_X1    g227(.A(new_n329), .ZN(new_n364));
  AOI22_X1  g228(.A1(new_n320), .A2(new_n364), .B1(new_n210), .B2(new_n211), .ZN(new_n365));
  AOI21_X1  g229(.A(new_n363), .B1(new_n365), .B2(G264), .ZN(new_n366));
  NAND3_X1  g230(.A1(new_n362), .A2(new_n233), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g231(.A(new_n367), .B1(new_n335), .B2(G200), .ZN(new_n368));
  NAND4_X1  g232(.A1(new_n368), .A2(new_n355), .A3(new_n359), .A4(new_n353), .ZN(new_n369));
  NAND2_X1  g233(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g234(.A1(new_n330), .A2(new_n171), .ZN(new_n371));
  NAND4_X1  g235(.A1(new_n184), .A2(new_n186), .A3(G244), .A4(new_n218), .ZN(new_n372));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g237(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g238(.A1(new_n217), .A2(KEYINPUT4), .A3(G244), .A4(new_n218), .ZN(new_n375));
  NAND2_X1  g239(.A1(G33), .A2(G283), .ZN(new_n376));
  NAND3_X1  g240(.A1(new_n217), .A2(G250), .A3(G1698), .ZN(new_n377));
  NAND4_X1  g241(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g242(.A(new_n371), .B1(new_n378), .B2(new_n223), .ZN(new_n379));
  NAND3_X1  g243(.A1(new_n379), .A2(new_n233), .A3(new_n323), .ZN(new_n380));
  AOI211_X1 g244(.A(new_n363), .B(new_n371), .C1(new_n223), .C2(new_n378), .ZN(new_n381));
  OAI21_X1  g245(.A(new_n380), .B1(new_n381), .B2(G200), .ZN(new_n382));
  NOR2_X1   g246(.A1(new_n203), .A2(G97), .ZN(new_n383));
  INV_X1    g247(.A(new_n383), .ZN(new_n384));
  INV_X1    g248(.A(new_n358), .ZN(new_n385));
  INV_X1    g249(.A(G97), .ZN(new_n386));
  NOR2_X1   g250(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g251(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g252(.A(new_n189), .B1(new_n217), .B2(G20), .ZN(new_n389));
  NAND3_X1  g253(.A1(new_n187), .A2(KEYINPUT7), .A3(new_n144), .ZN(new_n390));
  AOI21_X1  g254(.A(new_n157), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n392));
  OAI21_X1  g256(.A(new_n392), .B1(new_n386), .B2(G107), .ZN(new_n393));
  NAND3_X1  g257(.A1(new_n157), .A2(KEYINPUT6), .A3(G97), .ZN(new_n394));
  NAND2_X1  g258(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g259(.A1(new_n386), .A2(G107), .ZN(new_n396));
  AND3_X1   g260(.A1(new_n395), .A2(G20), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g261(.A1(new_n192), .A2(G77), .ZN(new_n398));
  INV_X1    g262(.A(new_n398), .ZN(new_n399));
  NOR3_X1   g263(.A1(new_n391), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g264(.A(new_n199), .ZN(new_n401));
  OAI211_X1 g265(.A(new_n384), .B(new_n388), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g266(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g267(.A1(new_n382), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g268(.A1(new_n184), .A2(new_n186), .A3(G238), .A4(new_n218), .ZN(new_n405));
  NAND4_X1  g269(.A1(new_n184), .A2(new_n186), .A3(G244), .A4(G1698), .ZN(new_n406));
  NAND3_X1  g270(.A1(new_n405), .A2(new_n406), .A3(new_n343), .ZN(new_n407));
  NAND2_X1  g271(.A1(new_n407), .A2(new_n223), .ZN(new_n408));
  AND2_X1   g272(.A1(G33), .A2(G41), .ZN(new_n409));
  OAI211_X1 g273(.A(new_n329), .B(G250), .C1(new_n409), .C2(new_n145), .ZN(new_n410));
  NAND3_X1  g274(.A1(new_n408), .A2(new_n321), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g275(.A1(new_n411), .A2(new_n226), .ZN(new_n412));
  INV_X1    g276(.A(new_n410), .ZN(new_n413));
  AOI211_X1 g277(.A(new_n322), .B(new_n413), .C1(new_n407), .C2(new_n223), .ZN(new_n414));
  NAND4_X1  g278(.A1(new_n184), .A2(new_n186), .A3(new_n144), .A4(G68), .ZN(new_n415));
  INV_X1    g279(.A(KEYINPUT19), .ZN(new_n416));
  OAI21_X1  g280(.A(new_n416), .B1(new_n242), .B2(new_n386), .ZN(new_n417));
  INV_X1    g281(.A(G87), .ZN(new_n418));
  NAND3_X1  g282(.A1(new_n418), .A2(new_n386), .A3(new_n157), .ZN(new_n419));
  NAND2_X1  g283(.A1(new_n419), .A2(G20), .ZN(new_n420));
  NAND4_X1  g284(.A1(new_n144), .A2(KEYINPUT19), .A3(G33), .A4(G97), .ZN(new_n421));
  NAND4_X1  g285(.A1(new_n415), .A2(new_n417), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  AOI22_X1  g286(.A1(new_n422), .A2(new_n199), .B1(new_n204), .B2(new_n300), .ZN(new_n423));
  INV_X1    g287(.A(new_n300), .ZN(new_n424));
  NAND2_X1  g288(.A1(new_n358), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g289(.A1(new_n414), .A2(new_n255), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g290(.A1(new_n408), .A2(new_n233), .A3(new_n321), .A4(new_n410), .ZN(new_n427));
  OAI21_X1  g291(.A(new_n427), .B1(new_n414), .B2(G200), .ZN(new_n428));
  NAND2_X1  g292(.A1(new_n358), .A2(G87), .ZN(new_n429));
  AND2_X1   g293(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g294(.A1(new_n412), .A2(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g295(.A1(new_n378), .A2(new_n223), .ZN(new_n432));
  INV_X1    g296(.A(new_n371), .ZN(new_n433));
  NAND3_X1  g297(.A1(new_n432), .A2(new_n323), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g298(.A1(new_n434), .A2(new_n226), .ZN(new_n435));
  NAND3_X1  g299(.A1(new_n379), .A2(new_n255), .A3(new_n323), .ZN(new_n436));
  NAND3_X1  g300(.A1(new_n402), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g301(.A1(new_n404), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g302(.A1(new_n203), .A2(G116), .ZN(new_n439));
  NOR3_X1   g303(.A1(new_n357), .A2(new_n204), .A3(new_n176), .ZN(new_n440));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n441));
  NOR2_X1   g305(.A1(new_n144), .A2(new_n176), .ZN(new_n442));
  OAI21_X1  g306(.A(new_n376), .B1(new_n386), .B2(G33), .ZN(new_n443));
  AOI21_X1  g307(.A(new_n442), .B1(new_n443), .B2(new_n144), .ZN(new_n444));
  OAI21_X1  g308(.A(new_n441), .B1(new_n444), .B2(new_n401), .ZN(new_n445));
  NAND2_X1  g309(.A1(new_n183), .A2(G97), .ZN(new_n446));
  AOI21_X1  g310(.A(G20), .B1(new_n446), .B2(new_n376), .ZN(new_n447));
  OAI211_X1 g311(.A(KEYINPUT20), .B(new_n199), .C1(new_n447), .C2(new_n442), .ZN(new_n448));
  AOI211_X1 g312(.A(new_n439), .B(new_n440), .C1(new_n445), .C2(new_n448), .ZN(new_n449));
  NAND4_X1  g313(.A1(new_n184), .A2(new_n186), .A3(G264), .A4(G1698), .ZN(new_n450));
  NAND4_X1  g314(.A1(new_n184), .A2(new_n186), .A3(G257), .A4(new_n218), .ZN(new_n451));
  INV_X1    g315(.A(G303), .ZN(new_n452));
  OAI211_X1 g316(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n217), .ZN(new_n453));
  NAND2_X1  g317(.A1(new_n453), .A2(new_n223), .ZN(new_n454));
  AOI21_X1  g318(.A(new_n363), .B1(new_n365), .B2(G270), .ZN(new_n455));
  NAND2_X1  g319(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g320(.A1(new_n456), .A2(G190), .ZN(new_n457));
  AOI21_X1  g321(.A(G200), .B1(new_n454), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g322(.A(new_n449), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g323(.A(KEYINPUT21), .ZN(new_n460));
  NAND2_X1  g324(.A1(new_n456), .A2(G169), .ZN(new_n461));
  OAI21_X1  g325(.A(new_n460), .B1(new_n461), .B2(new_n449), .ZN(new_n462));
  AOI21_X1  g326(.A(new_n439), .B1(new_n445), .B2(new_n448), .ZN(new_n463));
  OAI21_X1  g327(.A(new_n463), .B1(new_n176), .B2(new_n385), .ZN(new_n464));
  AOI21_X1  g328(.A(new_n226), .B1(new_n454), .B2(new_n455), .ZN(new_n465));
  NAND3_X1  g329(.A1(new_n464), .A2(KEYINPUT21), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g330(.A1(new_n456), .A2(new_n255), .ZN(new_n467));
  NAND2_X1  g331(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  NAND4_X1  g332(.A1(new_n459), .A2(new_n462), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NOR4_X1   g333(.A1(new_n319), .A2(new_n370), .A3(new_n438), .A4(new_n469), .ZN(G372));
  INV_X1    g334(.A(new_n258), .ZN(new_n471));
  INV_X1    g335(.A(new_n313), .ZN(new_n472));
  NAND4_X1  g336(.A1(new_n240), .A2(new_n298), .A3(new_n266), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g337(.A1(new_n297), .A2(new_n275), .ZN(new_n474));
  INV_X1    g338(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g339(.A1(new_n475), .A2(new_n240), .A3(new_n266), .ZN(new_n476));
  NAND2_X1  g340(.A1(new_n263), .A2(new_n265), .ZN(new_n477));
  AND3_X1   g341(.A1(new_n209), .A2(KEYINPUT18), .A3(new_n227), .ZN(new_n478));
  AOI21_X1  g342(.A(KEYINPUT18), .B1(new_n209), .B2(new_n227), .ZN(new_n479));
  NOR2_X1   g343(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g344(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AND4_X1   g345(.A1(new_n471), .A2(new_n473), .A3(new_n476), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g346(.A1(new_n423), .A2(new_n425), .ZN(new_n483));
  AOI21_X1  g347(.A(new_n322), .B1(new_n407), .B2(new_n223), .ZN(new_n484));
  NAND3_X1  g348(.A1(new_n484), .A2(new_n255), .A3(new_n410), .ZN(new_n485));
  NAND3_X1  g349(.A1(new_n412), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g350(.A1(new_n462), .A2(new_n466), .A3(new_n468), .ZN(new_n487));
  AOI22_X1  g351(.A1(new_n487), .A2(new_n369), .B1(new_n360), .B2(new_n337), .ZN(new_n488));
  OAI21_X1  g352(.A(new_n486), .B1(new_n488), .B2(new_n438), .ZN(new_n489));
  INV_X1    g353(.A(KEYINPUT26), .ZN(new_n490));
  AND4_X1   g354(.A1(new_n233), .A2(new_n408), .A3(new_n321), .A4(new_n410), .ZN(new_n491));
  AOI21_X1  g355(.A(G200), .B1(new_n484), .B2(new_n410), .ZN(new_n492));
  OAI21_X1  g356(.A(new_n430), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g357(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  OAI21_X1  g358(.A(new_n490), .B1(new_n437), .B2(new_n494), .ZN(new_n495));
  AND4_X1   g359(.A1(new_n255), .A2(new_n432), .A3(new_n323), .A4(new_n433), .ZN(new_n496));
  AOI21_X1  g360(.A(G169), .B1(new_n379), .B2(new_n323), .ZN(new_n497));
  NOR2_X1   g361(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g362(.A1(new_n431), .A2(KEYINPUT26), .A3(new_n498), .A4(new_n402), .ZN(new_n499));
  AND2_X1   g363(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g364(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g365(.A(new_n482), .B1(new_n319), .B2(new_n501), .ZN(G369));
  NAND3_X1  g366(.A1(new_n147), .A2(new_n144), .A3(G13), .ZN(new_n503));
  OR2_X1    g367(.A1(new_n503), .A2(KEYINPUT27), .ZN(new_n504));
  NAND2_X1  g368(.A1(new_n503), .A2(KEYINPUT27), .ZN(new_n505));
  NAND3_X1  g369(.A1(new_n504), .A2(G213), .A3(new_n505), .ZN(new_n506));
  INV_X1    g370(.A(G343), .ZN(new_n507));
  NOR2_X1   g371(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g372(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g373(.A1(new_n487), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g374(.A1(new_n360), .A2(new_n508), .ZN(new_n511));
  OR2_X1    g375(.A1(new_n370), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g376(.A1(new_n511), .A2(new_n337), .ZN(new_n513));
  AOI21_X1  g377(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g378(.A1(new_n449), .A2(new_n509), .ZN(new_n515));
  OR2_X1    g379(.A1(new_n469), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g380(.A1(new_n487), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g381(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g382(.A1(new_n518), .A2(G330), .ZN(new_n519));
  NAND2_X1  g383(.A1(new_n512), .A2(new_n513), .ZN(new_n520));
  AOI21_X1  g384(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g385(.A(new_n521), .B1(new_n361), .B2(new_n508), .ZN(G399));
  INV_X1    g386(.A(new_n148), .ZN(new_n523));
  NOR2_X1   g387(.A1(new_n523), .A2(G41), .ZN(new_n524));
  OR2_X1    g388(.A1(new_n419), .A2(G116), .ZN(new_n525));
  NOR3_X1   g389(.A1(new_n524), .A2(new_n147), .A3(new_n525), .ZN(new_n526));
  INV_X1    g390(.A(new_n143), .ZN(new_n527));
  AOI21_X1  g391(.A(new_n526), .B1(new_n527), .B2(new_n524), .ZN(new_n528));
  XOR2_X1   g392(.A(new_n528), .B(KEYINPUT28), .Z(new_n529));
  OAI21_X1  g393(.A(new_n509), .B1(new_n489), .B2(new_n500), .ZN(new_n530));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n531));
  NAND2_X1  g395(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g396(.A(KEYINPUT29), .B(new_n509), .C1(new_n489), .C2(new_n500), .ZN(new_n533));
  AND3_X1   g397(.A1(new_n404), .A2(new_n431), .A3(new_n437), .ZN(new_n534));
  INV_X1    g398(.A(new_n370), .ZN(new_n535));
  INV_X1    g399(.A(new_n469), .ZN(new_n536));
  NAND4_X1  g400(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n509), .ZN(new_n537));
  NAND4_X1  g401(.A1(new_n381), .A2(new_n467), .A3(new_n335), .A4(new_n414), .ZN(new_n538));
  INV_X1    g402(.A(KEYINPUT30), .ZN(new_n539));
  NAND2_X1  g403(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g404(.A1(new_n456), .A2(new_n411), .A3(new_n255), .ZN(new_n541));
  NAND4_X1  g405(.A1(new_n541), .A2(KEYINPUT30), .A3(new_n335), .A4(new_n381), .ZN(new_n542));
  NOR2_X1   g406(.A1(new_n335), .A2(G179), .ZN(new_n543));
  NAND4_X1  g407(.A1(new_n543), .A2(new_n411), .A3(new_n434), .A4(new_n456), .ZN(new_n544));
  NAND3_X1  g408(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g409(.A1(new_n545), .A2(new_n508), .ZN(new_n546));
  INV_X1    g410(.A(KEYINPUT31), .ZN(new_n547));
  NAND2_X1  g411(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g412(.A1(new_n545), .A2(KEYINPUT31), .A3(new_n508), .ZN(new_n549));
  NAND3_X1  g413(.A1(new_n537), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g414(.A1(new_n532), .A2(new_n533), .B1(G330), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g415(.A(new_n529), .B1(new_n551), .B2(G1), .ZN(G364));
  INV_X1    g416(.A(G13), .ZN(new_n553));
  NOR2_X1   g417(.A1(new_n553), .A2(G20), .ZN(new_n554));
  AOI21_X1  g418(.A(new_n147), .B1(new_n554), .B2(G45), .ZN(new_n555));
  INV_X1    g419(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g420(.A1(new_n524), .A2(new_n556), .ZN(new_n557));
  INV_X1    g421(.A(new_n557), .ZN(new_n558));
  INV_X1    g422(.A(new_n518), .ZN(new_n559));
  NOR2_X1   g423(.A1(G13), .A2(G33), .ZN(new_n560));
  INV_X1    g424(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g425(.A1(new_n561), .A2(G20), .ZN(new_n562));
  AOI21_X1  g426(.A(new_n558), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g427(.A(new_n145), .B1(G20), .B2(new_n226), .ZN(new_n564));
  NOR2_X1   g428(.A1(new_n144), .A2(new_n255), .ZN(new_n565));
  NAND2_X1  g429(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NOR2_X1   g430(.A1(new_n566), .A2(G190), .ZN(new_n567));
  XNOR2_X1  g431(.A(KEYINPUT33), .B(G317), .ZN(new_n568));
  NOR2_X1   g432(.A1(new_n144), .A2(new_n287), .ZN(new_n569));
  NAND3_X1  g433(.A1(new_n569), .A2(new_n255), .A3(G190), .ZN(new_n570));
  INV_X1    g434(.A(new_n570), .ZN(new_n571));
  AOI22_X1  g435(.A1(new_n567), .A2(new_n568), .B1(new_n571), .B2(G303), .ZN(new_n572));
  INV_X1    g436(.A(G311), .ZN(new_n573));
  NAND3_X1  g437(.A1(new_n565), .A2(new_n233), .A3(new_n287), .ZN(new_n574));
  OAI211_X1 g438(.A(new_n572), .B(new_n187), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g439(.A1(new_n566), .A2(new_n233), .ZN(new_n576));
  NAND3_X1  g440(.A1(new_n569), .A2(new_n255), .A3(new_n233), .ZN(new_n577));
  INV_X1    g441(.A(new_n577), .ZN(new_n578));
  AOI22_X1  g442(.A1(G326), .A2(new_n576), .B1(new_n578), .B2(G283), .ZN(new_n579));
  NOR2_X1   g443(.A1(G179), .A2(G200), .ZN(new_n580));
  NAND3_X1  g444(.A1(new_n580), .A2(G20), .A3(new_n233), .ZN(new_n581));
  INV_X1    g445(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g446(.A1(new_n582), .A2(G329), .ZN(new_n583));
  INV_X1    g447(.A(G294), .ZN(new_n584));
  AOI21_X1  g448(.A(new_n144), .B1(new_n580), .B2(G190), .ZN(new_n585));
  OAI211_X1 g449(.A(new_n579), .B(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g450(.A1(new_n565), .A2(G190), .A3(new_n287), .ZN(new_n587));
  INV_X1    g451(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g452(.A(new_n575), .B(new_n586), .C1(G322), .C2(new_n588), .ZN(new_n589));
  AOI22_X1  g453(.A1(G50), .A2(new_n576), .B1(new_n567), .B2(G68), .ZN(new_n590));
  INV_X1    g454(.A(new_n574), .ZN(new_n591));
  NAND2_X1  g455(.A1(new_n591), .A2(G77), .ZN(new_n592));
  NAND2_X1  g456(.A1(new_n571), .A2(G87), .ZN(new_n593));
  INV_X1    g457(.A(G159), .ZN(new_n594));
  OAI21_X1  g458(.A(KEYINPUT32), .B1(new_n581), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g459(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g460(.A1(new_n585), .A2(new_n386), .ZN(new_n597));
  AOI21_X1  g461(.A(new_n597), .B1(G58), .B2(new_n588), .ZN(new_n598));
  NAND2_X1  g462(.A1(new_n578), .A2(G107), .ZN(new_n599));
  OR3_X1    g463(.A1(new_n581), .A2(KEYINPUT32), .A3(new_n594), .ZN(new_n600));
  NAND4_X1  g464(.A1(new_n598), .A2(new_n217), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g465(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g466(.A(new_n564), .B1(new_n589), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g467(.A1(new_n562), .A2(new_n564), .ZN(new_n604));
  INV_X1    g468(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g469(.A1(new_n217), .A2(new_n148), .A3(G355), .ZN(new_n606));
  NOR2_X1   g470(.A1(new_n527), .A2(G45), .ZN(new_n607));
  AOI21_X1  g471(.A(new_n607), .B1(new_n181), .B2(G45), .ZN(new_n608));
  NOR2_X1   g472(.A1(new_n523), .A2(new_n217), .ZN(new_n609));
  INV_X1    g473(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g474(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g475(.A(new_n611), .B1(new_n176), .B2(new_n523), .ZN(new_n612));
  OAI211_X1 g476(.A(new_n563), .B(new_n603), .C1(new_n605), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g477(.A1(new_n518), .A2(G330), .ZN(new_n614));
  OR3_X1    g478(.A1(new_n519), .A2(new_n614), .A3(new_n557), .ZN(new_n615));
  NAND2_X1  g479(.A1(new_n613), .A2(new_n615), .ZN(G396));
  AOI22_X1  g480(.A1(new_n588), .A2(G143), .B1(new_n591), .B2(G159), .ZN(new_n617));
  INV_X1    g481(.A(G137), .ZN(new_n618));
  INV_X1    g482(.A(new_n576), .ZN(new_n619));
  INV_X1    g483(.A(G150), .ZN(new_n620));
  INV_X1    g484(.A(new_n567), .ZN(new_n621));
  OAI221_X1 g485(.A(new_n617), .B1(new_n618), .B2(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g486(.A(KEYINPUT34), .ZN(new_n623));
  AOI22_X1  g487(.A1(new_n622), .A2(new_n623), .B1(G50), .B2(new_n571), .ZN(new_n624));
  INV_X1    g488(.A(G132), .ZN(new_n625));
  OAI221_X1 g489(.A(new_n217), .B1(new_n581), .B2(new_n625), .C1(new_n138), .C2(new_n585), .ZN(new_n626));
  AOI21_X1  g490(.A(new_n626), .B1(G68), .B2(new_n578), .ZN(new_n627));
  OAI211_X1 g491(.A(new_n624), .B(new_n627), .C1(new_n623), .C2(new_n622), .ZN(new_n628));
  OAI22_X1  g492(.A1(new_n619), .A2(new_n452), .B1(new_n157), .B2(new_n570), .ZN(new_n629));
  AOI211_X1 g493(.A(new_n597), .B(new_n629), .C1(G294), .C2(new_n588), .ZN(new_n630));
  NOR2_X1   g494(.A1(new_n577), .A2(new_n418), .ZN(new_n631));
  INV_X1    g495(.A(G283), .ZN(new_n632));
  OAI21_X1  g496(.A(new_n187), .B1(new_n621), .B2(new_n632), .ZN(new_n633));
  AOI211_X1 g497(.A(new_n631), .B(new_n633), .C1(G116), .C2(new_n591), .ZN(new_n634));
  OAI211_X1 g498(.A(new_n630), .B(new_n634), .C1(new_n573), .C2(new_n581), .ZN(new_n635));
  NAND2_X1  g499(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g500(.A1(new_n636), .A2(new_n564), .ZN(new_n637));
  NOR2_X1   g501(.A1(new_n564), .A2(new_n560), .ZN(new_n638));
  AOI21_X1  g502(.A(new_n558), .B1(new_n180), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g503(.A1(new_n304), .A2(new_n508), .ZN(new_n640));
  NAND3_X1  g504(.A1(new_n313), .A2(new_n317), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g505(.A(new_n304), .B(new_n508), .C1(new_n311), .C2(new_n312), .ZN(new_n642));
  NAND2_X1  g506(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g507(.A(new_n637), .B(new_n639), .C1(new_n643), .C2(new_n561), .ZN(new_n644));
  NAND3_X1  g508(.A1(new_n530), .A2(new_n641), .A3(new_n642), .ZN(new_n645));
  OAI211_X1 g509(.A(new_n509), .B(new_n643), .C1(new_n489), .C2(new_n500), .ZN(new_n646));
  NAND2_X1  g510(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g511(.A1(new_n550), .A2(G330), .ZN(new_n648));
  XNOR2_X1  g512(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OAI21_X1  g513(.A(new_n644), .B1(new_n649), .B2(new_n557), .ZN(G384));
  AND2_X1   g514(.A1(new_n550), .A2(new_n643), .ZN(new_n651));
  NAND2_X1  g515(.A1(new_n275), .A2(new_n508), .ZN(new_n652));
  NAND2_X1  g516(.A1(new_n298), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g517(.A1(new_n297), .A2(new_n275), .A3(new_n508), .ZN(new_n654));
  NAND2_X1  g518(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g519(.A(new_n506), .ZN(new_n656));
  NAND2_X1  g520(.A1(new_n209), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g521(.A1(new_n230), .A2(new_n231), .ZN(new_n658));
  NAND2_X1  g522(.A1(new_n238), .A2(new_n239), .ZN(new_n659));
  AOI21_X1  g523(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g524(.A(new_n209), .B1(new_n227), .B2(new_n656), .ZN(new_n661));
  INV_X1    g525(.A(KEYINPUT37), .ZN(new_n662));
  AND3_X1   g526(.A1(new_n661), .A2(new_n662), .A3(new_n237), .ZN(new_n663));
  AOI21_X1  g527(.A(new_n662), .B1(new_n661), .B2(new_n237), .ZN(new_n664));
  NOR2_X1   g528(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g529(.A(KEYINPUT38), .ZN(new_n666));
  NOR3_X1   g530(.A1(new_n660), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g531(.A(new_n657), .ZN(new_n668));
  INV_X1    g532(.A(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g533(.A(new_n237), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g534(.A(new_n668), .B1(new_n480), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g535(.A1(new_n661), .A2(new_n237), .ZN(new_n672));
  NAND2_X1  g536(.A1(new_n672), .A2(KEYINPUT37), .ZN(new_n673));
  NAND3_X1  g537(.A1(new_n661), .A2(new_n662), .A3(new_n237), .ZN(new_n674));
  NAND2_X1  g538(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g539(.A(KEYINPUT38), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g540(.A(new_n651), .B(new_n655), .C1(new_n667), .C2(new_n676), .ZN(new_n677));
  INV_X1    g541(.A(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g542(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g543(.A(new_n666), .B1(new_n660), .B2(new_n665), .ZN(new_n680));
  NAND3_X1  g544(.A1(new_n671), .A2(new_n675), .A3(KEYINPUT38), .ZN(new_n681));
  NAND2_X1  g545(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g546(.A1(new_n682), .A2(KEYINPUT40), .A3(new_n655), .A4(new_n651), .ZN(new_n683));
  NAND2_X1  g547(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g548(.A(new_n319), .ZN(new_n685));
  NAND2_X1  g549(.A1(new_n685), .A2(new_n550), .ZN(new_n686));
  XOR2_X1   g550(.A(new_n684), .B(new_n686), .Z(new_n687));
  NAND2_X1  g551(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NOR2_X1   g552(.A1(new_n474), .A2(new_n508), .ZN(new_n689));
  INV_X1    g553(.A(new_n689), .ZN(new_n690));
  INV_X1    g554(.A(KEYINPUT39), .ZN(new_n691));
  AOI21_X1  g555(.A(new_n691), .B1(new_n680), .B2(new_n681), .ZN(new_n692));
  INV_X1    g556(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g557(.A1(new_n680), .A2(new_n691), .A3(new_n681), .ZN(new_n694));
  AOI21_X1  g558(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g559(.A(new_n682), .ZN(new_n696));
  NAND2_X1  g560(.A1(new_n472), .A2(new_n509), .ZN(new_n697));
  NAND2_X1  g561(.A1(new_n646), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g562(.A1(new_n698), .A2(new_n655), .ZN(new_n699));
  OAI22_X1  g563(.A1(new_n696), .A2(new_n699), .B1(new_n658), .B2(new_n656), .ZN(new_n700));
  NOR2_X1   g564(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g565(.A1(new_n532), .A2(new_n533), .ZN(new_n702));
  OAI21_X1  g566(.A(new_n482), .B1(new_n319), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g567(.A(new_n701), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g568(.A(new_n688), .B(new_n704), .ZN(new_n705));
  OAI21_X1  g569(.A(new_n705), .B1(new_n147), .B2(new_n554), .ZN(new_n706));
  AND2_X1   g570(.A1(new_n395), .A2(new_n396), .ZN(new_n707));
  AOI21_X1  g571(.A(new_n176), .B1(new_n707), .B2(KEYINPUT35), .ZN(new_n708));
  NOR2_X1   g572(.A1(new_n145), .A2(new_n144), .ZN(new_n709));
  OAI211_X1 g573(.A(new_n708), .B(new_n709), .C1(KEYINPUT35), .C2(new_n707), .ZN(new_n710));
  XNOR2_X1  g574(.A(new_n710), .B(KEYINPUT36), .ZN(new_n711));
  OR2_X1    g575(.A1(new_n178), .A2(new_n137), .ZN(new_n712));
  OAI22_X1  g576(.A1(new_n712), .A2(new_n180), .B1(G50), .B2(new_n139), .ZN(new_n713));
  NAND3_X1  g577(.A1(new_n713), .A2(G1), .A3(new_n553), .ZN(new_n714));
  NAND3_X1  g578(.A1(new_n706), .A2(new_n711), .A3(new_n714), .ZN(G367));
  OAI211_X1 g579(.A(new_n404), .B(new_n437), .C1(new_n403), .C2(new_n509), .ZN(new_n716));
  NAND3_X1  g580(.A1(new_n498), .A2(new_n402), .A3(new_n508), .ZN(new_n717));
  NAND2_X1  g581(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g582(.A1(new_n514), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g583(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  INV_X1    g584(.A(new_n718), .ZN(new_n721));
  OAI21_X1  g585(.A(new_n437), .B1(new_n721), .B2(new_n361), .ZN(new_n722));
  NAND2_X1  g586(.A1(new_n722), .A2(new_n509), .ZN(new_n723));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n724));
  NAND3_X1  g588(.A1(new_n514), .A2(new_n724), .A3(new_n718), .ZN(new_n725));
  NAND3_X1  g589(.A1(new_n720), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n727));
  NAND2_X1  g591(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g592(.A1(new_n430), .A2(new_n509), .ZN(new_n729));
  NAND2_X1  g593(.A1(new_n431), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g594(.A(new_n730), .B1(new_n486), .B2(new_n729), .ZN(new_n731));
  INV_X1    g595(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g596(.A1(new_n720), .A2(new_n723), .A3(KEYINPUT43), .A4(new_n725), .ZN(new_n733));
  NAND3_X1  g597(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g598(.A1(new_n726), .A2(new_n727), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g599(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g600(.A1(new_n519), .A2(new_n520), .ZN(new_n737));
  NOR2_X1   g601(.A1(new_n737), .A2(new_n721), .ZN(new_n738));
  XNOR2_X1  g602(.A(new_n736), .B(new_n738), .ZN(new_n739));
  XOR2_X1   g603(.A(new_n524), .B(KEYINPUT41), .Z(new_n740));
  NOR2_X1   g604(.A1(new_n361), .A2(new_n508), .ZN(new_n741));
  NOR3_X1   g605(.A1(new_n514), .A2(new_n741), .A3(new_n721), .ZN(new_n742));
  XNOR2_X1  g606(.A(new_n742), .B(KEYINPUT45), .ZN(new_n743));
  OAI21_X1  g607(.A(new_n721), .B1(new_n514), .B2(new_n741), .ZN(new_n744));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n745));
  XNOR2_X1  g609(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g610(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g611(.A(new_n737), .ZN(new_n748));
  NAND2_X1  g612(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g613(.A(new_n510), .ZN(new_n750));
  NOR3_X1   g614(.A1(new_n519), .A2(new_n520), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g615(.A1(new_n748), .A2(new_n751), .A3(new_n514), .ZN(new_n752));
  NAND2_X1  g616(.A1(new_n752), .A2(new_n551), .ZN(new_n753));
  INV_X1    g617(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g618(.A1(new_n743), .A2(new_n746), .A3(new_n737), .ZN(new_n755));
  NAND3_X1  g619(.A1(new_n749), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g620(.A(new_n740), .B1(new_n756), .B2(new_n551), .ZN(new_n757));
  OAI21_X1  g621(.A(new_n739), .B1(new_n757), .B2(new_n556), .ZN(new_n758));
  OR3_X1    g622(.A1(new_n570), .A2(KEYINPUT46), .A3(new_n176), .ZN(new_n759));
  OAI21_X1  g623(.A(KEYINPUT46), .B1(new_n570), .B2(new_n176), .ZN(new_n760));
  NAND2_X1  g624(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g625(.A(new_n761), .B1(new_n584), .B2(new_n621), .ZN(new_n762));
  AOI211_X1 g626(.A(new_n217), .B(new_n762), .C1(G317), .C2(new_n582), .ZN(new_n763));
  OAI221_X1 g627(.A(new_n763), .B1(new_n386), .B2(new_n577), .C1(new_n632), .C2(new_n574), .ZN(new_n764));
  INV_X1    g628(.A(new_n585), .ZN(new_n765));
  AOI22_X1  g629(.A1(new_n588), .A2(G303), .B1(new_n765), .B2(G107), .ZN(new_n766));
  OAI21_X1  g630(.A(new_n766), .B1(new_n573), .B2(new_n619), .ZN(new_n767));
  AOI22_X1  g631(.A1(new_n571), .A2(G58), .B1(new_n591), .B2(G50), .ZN(new_n768));
  NAND2_X1  g632(.A1(new_n576), .A2(G143), .ZN(new_n769));
  OAI211_X1 g633(.A(new_n768), .B(new_n769), .C1(new_n620), .C2(new_n587), .ZN(new_n770));
  AOI21_X1  g634(.A(new_n770), .B1(G159), .B2(new_n567), .ZN(new_n771));
  NAND2_X1  g635(.A1(new_n765), .A2(G68), .ZN(new_n772));
  NAND3_X1  g636(.A1(new_n771), .A2(new_n217), .A3(new_n772), .ZN(new_n773));
  OAI22_X1  g637(.A1(new_n577), .A2(new_n180), .B1(new_n618), .B2(new_n581), .ZN(new_n774));
  OAI22_X1  g638(.A1(new_n764), .A2(new_n767), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g639(.A(new_n775), .B(KEYINPUT47), .ZN(new_n776));
  NAND2_X1  g640(.A1(new_n776), .A2(new_n564), .ZN(new_n777));
  NAND2_X1  g641(.A1(new_n732), .A2(new_n562), .ZN(new_n778));
  OAI221_X1 g642(.A(new_n604), .B1(new_n148), .B2(new_n300), .C1(new_n172), .C2(new_n610), .ZN(new_n779));
  NAND4_X1  g643(.A1(new_n777), .A2(new_n557), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g644(.A1(new_n758), .A2(new_n780), .ZN(G387));
  NAND2_X1  g645(.A1(new_n752), .A2(new_n556), .ZN(new_n782));
  OAI21_X1  g646(.A(new_n187), .B1(new_n577), .B2(new_n176), .ZN(new_n783));
  AOI22_X1  g647(.A1(G311), .A2(new_n567), .B1(new_n588), .B2(G317), .ZN(new_n784));
  AOI22_X1  g648(.A1(G322), .A2(new_n576), .B1(new_n591), .B2(G303), .ZN(new_n785));
  NAND2_X1  g649(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g650(.A(KEYINPUT48), .ZN(new_n787));
  AOI22_X1  g651(.A1(new_n786), .A2(new_n787), .B1(G294), .B2(new_n571), .ZN(new_n788));
  OAI221_X1 g652(.A(new_n788), .B1(new_n787), .B2(new_n786), .C1(new_n632), .C2(new_n585), .ZN(new_n789));
  XOR2_X1   g653(.A(new_n789), .B(KEYINPUT49), .Z(new_n790));
  AOI211_X1 g654(.A(new_n783), .B(new_n790), .C1(G326), .C2(new_n582), .ZN(new_n791));
  NAND2_X1  g655(.A1(new_n765), .A2(new_n424), .ZN(new_n792));
  NAND2_X1  g656(.A1(new_n792), .A2(new_n217), .ZN(new_n793));
  NOR2_X1   g657(.A1(new_n570), .A2(new_n180), .ZN(new_n794));
  OAI22_X1  g658(.A1(new_n577), .A2(new_n386), .B1(new_n587), .B2(new_n137), .ZN(new_n795));
  AOI211_X1 g659(.A(new_n794), .B(new_n795), .C1(G159), .C2(new_n576), .ZN(new_n796));
  OAI221_X1 g660(.A(new_n796), .B1(new_n620), .B2(new_n581), .C1(new_n202), .C2(new_n621), .ZN(new_n797));
  AOI211_X1 g661(.A(new_n793), .B(new_n797), .C1(G68), .C2(new_n591), .ZN(new_n798));
  OAI21_X1  g662(.A(new_n564), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g663(.A1(new_n525), .A2(new_n148), .A3(new_n217), .ZN(new_n800));
  INV_X1    g664(.A(G45), .ZN(new_n801));
  NOR2_X1   g665(.A1(new_n168), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g666(.A(new_n525), .B1(G68), .B2(G77), .ZN(new_n803));
  AOI21_X1  g667(.A(KEYINPUT50), .B1(new_n207), .B2(new_n137), .ZN(new_n804));
  AND3_X1   g668(.A1(new_n207), .A2(KEYINPUT50), .A3(new_n137), .ZN(new_n805));
  OAI211_X1 g669(.A(new_n803), .B(new_n801), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g670(.A1(new_n806), .A2(new_n609), .ZN(new_n807));
  OAI221_X1 g671(.A(new_n800), .B1(G107), .B2(new_n148), .C1(new_n802), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g672(.A1(new_n808), .A2(new_n604), .ZN(new_n809));
  NAND3_X1  g673(.A1(new_n512), .A2(new_n513), .A3(new_n562), .ZN(new_n810));
  NAND4_X1  g674(.A1(new_n799), .A2(new_n557), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g675(.A(new_n524), .B1(new_n752), .B2(new_n551), .ZN(new_n812));
  OAI211_X1 g676(.A(new_n782), .B(new_n811), .C1(new_n754), .C2(new_n812), .ZN(G393));
  AND3_X1   g677(.A1(new_n743), .A2(new_n737), .A3(new_n746), .ZN(new_n814));
  AOI21_X1  g678(.A(new_n737), .B1(new_n743), .B2(new_n746), .ZN(new_n815));
  OAI21_X1  g679(.A(new_n753), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g680(.A1(new_n816), .A2(new_n756), .A3(new_n524), .ZN(new_n817));
  AND2_X1   g681(.A1(new_n177), .A2(new_n609), .ZN(new_n818));
  OAI21_X1  g682(.A(new_n604), .B1(new_n386), .B2(new_n148), .ZN(new_n819));
  INV_X1    g683(.A(new_n562), .ZN(new_n820));
  OAI221_X1 g684(.A(new_n557), .B1(new_n818), .B2(new_n819), .C1(new_n718), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g685(.A1(G317), .A2(new_n576), .B1(new_n588), .B2(G311), .ZN(new_n822));
  XNOR2_X1  g686(.A(new_n822), .B(KEYINPUT52), .ZN(new_n823));
  AOI21_X1  g687(.A(new_n823), .B1(G116), .B2(new_n765), .ZN(new_n824));
  NAND2_X1  g688(.A1(new_n571), .A2(G283), .ZN(new_n825));
  OAI221_X1 g689(.A(new_n187), .B1(new_n584), .B2(new_n574), .C1(new_n621), .C2(new_n452), .ZN(new_n826));
  AOI21_X1  g690(.A(new_n826), .B1(G322), .B2(new_n582), .ZN(new_n827));
  NAND4_X1  g691(.A1(new_n824), .A2(new_n599), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  AOI22_X1  g692(.A1(G150), .A2(new_n576), .B1(new_n588), .B2(G159), .ZN(new_n829));
  XNOR2_X1  g693(.A(new_n829), .B(KEYINPUT51), .ZN(new_n830));
  AOI21_X1  g694(.A(new_n830), .B1(G68), .B2(new_n571), .ZN(new_n831));
  NAND2_X1  g695(.A1(new_n765), .A2(G77), .ZN(new_n832));
  NAND2_X1  g696(.A1(new_n591), .A2(new_n207), .ZN(new_n833));
  OAI221_X1 g697(.A(new_n217), .B1(new_n418), .B2(new_n577), .C1(new_n621), .C2(new_n137), .ZN(new_n834));
  AOI21_X1  g698(.A(new_n834), .B1(G143), .B2(new_n582), .ZN(new_n835));
  NAND4_X1  g699(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g700(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g701(.A(new_n821), .B1(new_n564), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g702(.A1(new_n814), .A2(new_n815), .ZN(new_n839));
  AOI21_X1  g703(.A(new_n838), .B1(new_n839), .B2(new_n556), .ZN(new_n840));
  AND2_X1   g704(.A1(new_n817), .A2(new_n840), .ZN(new_n841));
  INV_X1    g705(.A(new_n841), .ZN(G390));
  NAND4_X1  g706(.A1(new_n655), .A2(new_n550), .A3(G330), .A4(new_n643), .ZN(new_n843));
  INV_X1    g707(.A(new_n843), .ZN(new_n844));
  AND3_X1   g708(.A1(new_n680), .A2(new_n691), .A3(new_n681), .ZN(new_n845));
  AOI21_X1  g709(.A(new_n689), .B1(new_n698), .B2(new_n655), .ZN(new_n846));
  NOR3_X1   g710(.A1(new_n845), .A2(new_n692), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g711(.A1(new_n846), .A2(new_n682), .ZN(new_n848));
  INV_X1    g712(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g713(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g714(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g715(.A1(new_n699), .A2(new_n690), .ZN(new_n852));
  NAND3_X1  g716(.A1(new_n693), .A2(new_n852), .A3(new_n694), .ZN(new_n853));
  NAND3_X1  g717(.A1(new_n853), .A2(new_n843), .A3(new_n848), .ZN(new_n854));
  INV_X1    g718(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g719(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g720(.A1(new_n588), .A2(G132), .B1(new_n765), .B2(G159), .ZN(new_n857));
  INV_X1    g721(.A(G128), .ZN(new_n858));
  OAI221_X1 g722(.A(new_n857), .B1(new_n137), .B2(new_n577), .C1(new_n858), .C2(new_n619), .ZN(new_n859));
  NOR2_X1   g723(.A1(new_n570), .A2(new_n620), .ZN(new_n860));
  XNOR2_X1  g724(.A(new_n860), .B(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g725(.A1(new_n582), .A2(G125), .ZN(new_n862));
  XNOR2_X1  g726(.A(KEYINPUT54), .B(G143), .ZN(new_n863));
  OR2_X1    g727(.A1(new_n574), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g728(.A1(new_n861), .A2(new_n217), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  AOI211_X1 g729(.A(new_n859), .B(new_n865), .C1(G137), .C2(new_n567), .ZN(new_n866));
  AOI22_X1  g730(.A1(G283), .A2(new_n576), .B1(new_n571), .B2(G87), .ZN(new_n867));
  OAI221_X1 g731(.A(new_n867), .B1(new_n139), .B2(new_n577), .C1(new_n176), .C2(new_n587), .ZN(new_n868));
  NOR2_X1   g732(.A1(new_n574), .A2(new_n386), .ZN(new_n869));
  NOR2_X1   g733(.A1(new_n581), .A2(new_n584), .ZN(new_n870));
  OAI211_X1 g734(.A(new_n187), .B(new_n832), .C1(new_n621), .C2(new_n157), .ZN(new_n871));
  NOR4_X1   g735(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g736(.A(new_n564), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g737(.A1(new_n845), .A2(new_n692), .A3(new_n561), .ZN(new_n874));
  AOI211_X1 g738(.A(new_n558), .B(new_n874), .C1(new_n202), .C2(new_n638), .ZN(new_n875));
  AOI22_X1  g739(.A1(new_n856), .A2(new_n556), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g740(.A(new_n482), .B1(new_n551), .B2(new_n319), .ZN(new_n877));
  NAND3_X1  g741(.A1(new_n550), .A2(G330), .A3(new_n643), .ZN(new_n878));
  AOI22_X1  g742(.A1(new_n475), .A2(new_n508), .B1(new_n298), .B2(new_n652), .ZN(new_n879));
  NAND2_X1  g743(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g744(.A1(new_n843), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g745(.A1(new_n881), .A2(new_n698), .ZN(new_n882));
  INV_X1    g746(.A(new_n698), .ZN(new_n883));
  NAND3_X1  g747(.A1(new_n843), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g748(.A(new_n877), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g749(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g750(.A(new_n886), .B1(new_n851), .B2(new_n855), .ZN(new_n887));
  NAND3_X1  g751(.A1(new_n850), .A2(new_n854), .A3(new_n885), .ZN(new_n888));
  NAND3_X1  g752(.A1(new_n887), .A2(new_n524), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g753(.A1(new_n876), .A2(new_n889), .ZN(G378));
  NAND3_X1  g754(.A1(new_n679), .A2(G330), .A3(new_n683), .ZN(new_n891));
  NAND2_X1  g755(.A1(new_n247), .A2(new_n656), .ZN(new_n892));
  XOR2_X1   g756(.A(new_n892), .B(KEYINPUT55), .Z(new_n893));
  XNOR2_X1  g757(.A(new_n893), .B(KEYINPUT56), .ZN(new_n894));
  XOR2_X1   g758(.A(new_n266), .B(new_n894), .Z(new_n895));
  NAND2_X1  g759(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g760(.A(new_n895), .ZN(new_n897));
  NAND4_X1  g761(.A1(new_n679), .A2(G330), .A3(new_n683), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g762(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g763(.A(new_n701), .ZN(new_n900));
  NAND2_X1  g764(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g765(.A1(new_n896), .A2(new_n701), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g766(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g767(.A1(new_n903), .A2(new_n556), .ZN(new_n904));
  NAND2_X1  g768(.A1(new_n895), .A2(new_n560), .ZN(new_n905));
  OAI22_X1  g769(.A1(new_n574), .A2(new_n618), .B1(new_n585), .B2(new_n620), .ZN(new_n906));
  NAND2_X1  g770(.A1(new_n588), .A2(G128), .ZN(new_n907));
  OAI221_X1 g771(.A(new_n907), .B1(new_n570), .B2(new_n863), .C1(new_n621), .C2(new_n625), .ZN(new_n908));
  AOI211_X1 g772(.A(new_n906), .B(new_n908), .C1(G125), .C2(new_n576), .ZN(new_n909));
  XNOR2_X1  g773(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  AOI211_X1 g774(.A(G33), .B(G41), .C1(new_n582), .C2(G124), .ZN(new_n911));
  OAI211_X1 g775(.A(new_n910), .B(new_n911), .C1(new_n594), .C2(new_n577), .ZN(new_n912));
  NOR2_X1   g776(.A1(new_n217), .A2(G41), .ZN(new_n913));
  OAI21_X1  g777(.A(new_n137), .B1(G33), .B2(G41), .ZN(new_n914));
  OAI21_X1  g778(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g779(.A1(G116), .A2(new_n576), .B1(new_n591), .B2(new_n424), .ZN(new_n916));
  NAND2_X1  g780(.A1(new_n578), .A2(G58), .ZN(new_n917));
  OAI211_X1 g781(.A(new_n916), .B(new_n917), .C1(new_n157), .C2(new_n587), .ZN(new_n918));
  AOI211_X1 g782(.A(new_n794), .B(new_n918), .C1(G97), .C2(new_n567), .ZN(new_n919));
  NAND2_X1  g783(.A1(new_n582), .A2(G283), .ZN(new_n920));
  NAND4_X1  g784(.A1(new_n919), .A2(new_n772), .A3(new_n913), .A4(new_n920), .ZN(new_n921));
  XOR2_X1   g785(.A(new_n921), .B(KEYINPUT58), .Z(new_n922));
  OAI21_X1  g786(.A(new_n564), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g787(.A1(new_n638), .A2(new_n137), .ZN(new_n924));
  NAND4_X1  g788(.A1(new_n905), .A2(new_n557), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g789(.A1(new_n904), .A2(new_n925), .ZN(new_n926));
  INV_X1    g790(.A(new_n877), .ZN(new_n927));
  NAND2_X1  g791(.A1(new_n888), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g792(.A1(new_n896), .A2(new_n701), .A3(new_n898), .ZN(new_n929));
  AOI21_X1  g793(.A(new_n701), .B1(new_n896), .B2(new_n898), .ZN(new_n930));
  OAI21_X1  g794(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g795(.A1(new_n931), .A2(KEYINPUT57), .ZN(new_n932));
  INV_X1    g796(.A(KEYINPUT57), .ZN(new_n933));
  OAI211_X1 g797(.A(new_n928), .B(new_n933), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g798(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g799(.A(new_n926), .B1(new_n935), .B2(new_n524), .ZN(new_n936));
  INV_X1    g800(.A(new_n936), .ZN(G375));
  NAND2_X1  g801(.A1(new_n882), .A2(new_n884), .ZN(new_n938));
  NOR2_X1   g802(.A1(new_n938), .A2(new_n927), .ZN(new_n939));
  INV_X1    g803(.A(new_n939), .ZN(new_n940));
  INV_X1    g804(.A(new_n740), .ZN(new_n941));
  NAND3_X1  g805(.A1(new_n940), .A2(new_n941), .A3(new_n886), .ZN(new_n942));
  OAI22_X1  g806(.A1(new_n619), .A2(new_n625), .B1(new_n618), .B2(new_n587), .ZN(new_n943));
  AOI21_X1  g807(.A(new_n943), .B1(G150), .B2(new_n591), .ZN(new_n944));
  OAI221_X1 g808(.A(new_n944), .B1(new_n137), .B2(new_n585), .C1(new_n858), .C2(new_n581), .ZN(new_n945));
  AOI21_X1  g809(.A(new_n187), .B1(new_n571), .B2(G159), .ZN(new_n946));
  OAI211_X1 g810(.A(new_n946), .B(new_n917), .C1(new_n621), .C2(new_n863), .ZN(new_n947));
  AOI22_X1  g811(.A1(G294), .A2(new_n576), .B1(new_n578), .B2(G77), .ZN(new_n948));
  AND2_X1   g812(.A1(new_n948), .A2(new_n792), .ZN(new_n949));
  OAI221_X1 g813(.A(new_n949), .B1(new_n632), .B2(new_n587), .C1(new_n452), .C2(new_n581), .ZN(new_n950));
  AOI21_X1  g814(.A(new_n217), .B1(new_n571), .B2(G97), .ZN(new_n951));
  OAI221_X1 g815(.A(new_n951), .B1(new_n157), .B2(new_n574), .C1(new_n176), .C2(new_n621), .ZN(new_n952));
  OAI22_X1  g816(.A1(new_n945), .A2(new_n947), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g817(.A1(new_n953), .A2(new_n564), .ZN(new_n954));
  AOI21_X1  g818(.A(new_n558), .B1(new_n139), .B2(new_n638), .ZN(new_n955));
  OAI211_X1 g819(.A(new_n954), .B(new_n955), .C1(new_n655), .C2(new_n561), .ZN(new_n956));
  INV_X1    g820(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g821(.A(new_n957), .B1(new_n938), .B2(new_n556), .ZN(new_n958));
  NAND2_X1  g822(.A1(new_n942), .A2(new_n958), .ZN(G381));
  INV_X1    g823(.A(G378), .ZN(new_n960));
  NAND2_X1  g824(.A1(new_n936), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g825(.A1(new_n961), .A2(G381), .ZN(new_n962));
  INV_X1    g826(.A(G396), .ZN(new_n963));
  INV_X1    g827(.A(G393), .ZN(new_n964));
  NAND3_X1  g828(.A1(new_n758), .A2(new_n841), .A3(new_n780), .ZN(new_n965));
  NOR2_X1   g829(.A1(new_n965), .A2(G384), .ZN(new_n966));
  NAND4_X1  g830(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n966), .ZN(G407));
  OAI211_X1 g831(.A(G407), .B(G213), .C1(G343), .C2(new_n961), .ZN(G409));
  INV_X1    g832(.A(new_n965), .ZN(new_n969));
  AOI21_X1  g833(.A(new_n841), .B1(new_n758), .B2(new_n780), .ZN(new_n970));
  NOR3_X1   g834(.A1(new_n969), .A2(new_n970), .A3(G393), .ZN(new_n971));
  NAND2_X1  g835(.A1(G387), .A2(G390), .ZN(new_n972));
  AOI21_X1  g836(.A(new_n964), .B1(new_n972), .B2(new_n965), .ZN(new_n973));
  OAI21_X1  g837(.A(G396), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g838(.A(G393), .B1(new_n969), .B2(new_n970), .ZN(new_n975));
  NAND3_X1  g839(.A1(new_n972), .A2(new_n964), .A3(new_n965), .ZN(new_n976));
  NAND3_X1  g840(.A1(new_n975), .A2(new_n976), .A3(new_n963), .ZN(new_n977));
  NAND2_X1  g841(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g842(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g843(.A1(new_n507), .A2(G213), .ZN(new_n980));
  AND2_X1   g844(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n981));
  NOR2_X1   g845(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n982));
  OAI211_X1 g846(.A(new_n524), .B(new_n886), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  AND3_X1   g847(.A1(new_n983), .A2(G384), .A3(new_n958), .ZN(new_n984));
  AOI21_X1  g848(.A(G384), .B1(new_n983), .B2(new_n958), .ZN(new_n985));
  NOR2_X1   g849(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g850(.A(new_n524), .ZN(new_n987));
  AOI21_X1  g851(.A(new_n987), .B1(new_n932), .B2(new_n934), .ZN(new_n988));
  NOR3_X1   g852(.A1(new_n988), .A2(new_n960), .A3(new_n926), .ZN(new_n989));
  INV_X1    g853(.A(new_n925), .ZN(new_n990));
  AOI21_X1  g854(.A(new_n990), .B1(new_n903), .B2(new_n556), .ZN(new_n991));
  NAND3_X1  g855(.A1(new_n903), .A2(new_n941), .A3(new_n928), .ZN(new_n992));
  AOI21_X1  g856(.A(G378), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g857(.A(new_n980), .B(new_n986), .C1(new_n989), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g858(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  INV_X1    g859(.A(new_n986), .ZN(new_n996));
  INV_X1    g860(.A(new_n980), .ZN(new_n997));
  NAND2_X1  g861(.A1(new_n997), .A2(G2897), .ZN(new_n998));
  AOI21_X1  g862(.A(new_n993), .B1(new_n936), .B2(G378), .ZN(new_n999));
  OAI211_X1 g863(.A(new_n996), .B(new_n998), .C1(new_n999), .C2(new_n997), .ZN(new_n1000));
  NOR2_X1   g864(.A1(new_n996), .A2(new_n998), .ZN(new_n1001));
  INV_X1    g865(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g866(.A1(new_n995), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g867(.A(KEYINPUT61), .ZN(new_n1004));
  OAI21_X1  g868(.A(new_n1004), .B1(new_n994), .B2(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g869(.A(new_n979), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AND3_X1   g870(.A1(new_n1000), .A2(new_n1004), .A3(new_n978), .ZN(new_n1007));
  NAND2_X1  g871(.A1(new_n994), .A2(KEYINPUT63), .ZN(new_n1008));
  NAND2_X1  g872(.A1(new_n935), .A2(new_n524), .ZN(new_n1009));
  NAND3_X1  g873(.A1(new_n1009), .A2(G378), .A3(new_n991), .ZN(new_n1010));
  INV_X1    g874(.A(new_n993), .ZN(new_n1011));
  NAND2_X1  g875(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g876(.A(KEYINPUT63), .ZN(new_n1013));
  NAND4_X1  g877(.A1(new_n1012), .A2(new_n1013), .A3(new_n980), .A4(new_n986), .ZN(new_n1014));
  AOI21_X1  g878(.A(new_n1001), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g879(.A1(new_n1007), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g880(.A1(new_n1006), .A2(new_n1016), .ZN(G405));
  NAND2_X1  g881(.A1(G375), .A2(G378), .ZN(new_n1018));
  NAND2_X1  g882(.A1(new_n1018), .A2(new_n961), .ZN(new_n1019));
  NAND2_X1  g883(.A1(new_n1019), .A2(new_n996), .ZN(new_n1020));
  NAND3_X1  g884(.A1(new_n1018), .A2(new_n961), .A3(new_n986), .ZN(new_n1021));
  AND3_X1   g885(.A1(new_n979), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g886(.A(new_n979), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1023));
  NOR2_X1   g887(.A1(new_n1022), .A2(new_n1023), .ZN(G402));
endmodule


