//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n463), .B1(new_n460), .B2(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  AOI21_X1  g050(.A(new_n468), .B1(new_n464), .B2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n472), .A2(new_n483), .A3(G138), .A4(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n468), .A2(G138), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n464), .B2(new_n466), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n468), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n476), .B2(G126), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  XNOR2_X1  g068(.A(KEYINPUT68), .B(G651), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(G543), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT69), .A2(G543), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n495), .B(KEYINPUT5), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT5), .B1(new_n496), .B2(new_n497), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT70), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(G62), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n510), .A2(new_n503), .A3(new_n500), .A4(new_n498), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n506), .A2(new_n515), .ZN(G166));
  AND2_X1   g091(.A1(G63), .A2(G651), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n503), .A2(new_n500), .A3(new_n498), .A4(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n501), .A2(KEYINPUT71), .A3(new_n503), .A4(new_n517), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT68), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n509), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(G51), .B(G543), .C1(new_n529), .C2(new_n507), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n524), .B(new_n530), .C1(new_n511), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n522), .A2(new_n532), .ZN(G168));
  NAND3_X1  g108(.A1(new_n501), .A2(G64), .A3(new_n503), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n494), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n528), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n499), .B1(new_n538), .B2(new_n508), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n511), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n536), .A2(new_n542), .ZN(G171));
  NAND4_X1  g118(.A1(new_n503), .A2(G56), .A3(new_n500), .A4(new_n498), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n537), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n501), .A2(G81), .A3(new_n503), .A4(new_n510), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT72), .B(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n539), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n550), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n494), .B1(new_n544), .B2(new_n545), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n501), .A2(new_n503), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI211_X1 g141(.A(KEYINPUT74), .B(KEYINPUT9), .C1(new_n514), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n539), .A2(G53), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n565), .A2(G651), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n511), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n501), .A2(KEYINPUT75), .A3(new_n503), .A4(new_n510), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G91), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n534), .A2(new_n535), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(new_n537), .ZN(new_n577));
  INV_X1    g152(.A(new_n511), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G90), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n577), .A2(KEYINPUT76), .A3(new_n540), .A4(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(new_n536), .B2(new_n542), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(G301));
  OAI21_X1  g158(.A(KEYINPUT77), .B1(new_n522), .B2(new_n532), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n530), .A2(new_n524), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n578), .B2(G89), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n520), .A2(new_n521), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n585), .A2(new_n591), .ZN(G286));
  INV_X1    g167(.A(G166), .ZN(G303));
  INV_X1    g168(.A(G74), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n525), .B1(new_n563), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n572), .A2(G87), .A3(new_n573), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G288));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n563), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(new_n537), .B1(G48), .B2(new_n539), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n572), .A2(G86), .A3(new_n573), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G305));
  NAND3_X1  g183(.A1(new_n501), .A2(G60), .A3(new_n503), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n494), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT79), .B(G47), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n511), .A2(new_n612), .B1(new_n514), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n611), .A2(new_n614), .ZN(G290));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(G301), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(G66), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n503), .A2(new_n500), .A3(new_n498), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT80), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G651), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n539), .A2(G54), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n572), .A2(G92), .A3(new_n573), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n573), .A4(G92), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n617), .B1(new_n631), .B2(new_n616), .ZN(G284));
  AOI21_X1  g207(.A(new_n617), .B1(new_n631), .B2(new_n616), .ZN(G321));
  NOR2_X1   g208(.A1(G286), .A2(new_n616), .ZN(new_n634));
  XNOR2_X1  g209(.A(G299), .B(KEYINPUT83), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n616), .ZN(G297));
  AOI21_X1  g211(.A(new_n634), .B1(new_n635), .B2(new_n616), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n631), .B1(new_n638), .B2(G860), .ZN(G148));
  OAI21_X1  g214(.A(KEYINPUT85), .B1(new_n556), .B2(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n631), .A2(new_n638), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT84), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n631), .A2(new_n643), .A3(new_n638), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n616), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  MUX2_X1   g220(.A(new_n640), .B(KEYINPUT85), .S(new_n645), .Z(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n472), .A2(new_n461), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  INV_X1    g226(.A(new_n469), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G135), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n476), .A2(G123), .ZN(new_n654));
  OR2_X1    g229(.A1(G99), .A2(G2105), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n655), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n658), .ZN(G156));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT87), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1341), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1348), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n673), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(G401));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n680), .B2(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2096), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NOR3_X1   g273(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(G229));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G11), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT96), .B(G28), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT30), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n710), .A2(KEYINPUT30), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n657), .B2(G29), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT97), .Z(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G21), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G168), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT95), .B(G1966), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(G5), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G171), .B2(new_n718), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n717), .B(new_n722), .C1(G1961), .C2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT98), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT26), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n729), .A2(new_n730), .B1(G105), .B2(new_n461), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n476), .A2(G129), .ZN(new_n732));
  INV_X1    g307(.A(G141), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n469), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(new_n712), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n712), .B2(G32), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT27), .B(G1996), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n712), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  INV_X1    g322(.A(G139), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n469), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n468), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n745), .B1(new_n753), .B2(new_n712), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G2072), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(G2072), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n743), .A2(new_n744), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n718), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n556), .B2(new_n718), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G1341), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(G1341), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n712), .B1(KEYINPUT24), .B2(G34), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(KEYINPUT24), .B2(G34), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2084), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n712), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n652), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n476), .A2(G128), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n712), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n712), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n779));
  INV_X1    g354(.A(G2090), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n778), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n724), .A2(G1961), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n712), .A2(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n712), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2078), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n776), .A2(new_n782), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n757), .A2(new_n760), .A3(new_n761), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n726), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G4), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n631), .B2(G16), .ZN(new_n791));
  INV_X1    g366(.A(G1348), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n718), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT23), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT100), .ZN(new_n797));
  INV_X1    g372(.A(G1956), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n789), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n718), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n718), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  AND2_X1   g380(.A1(new_n718), .A2(G6), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G305), .B2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n718), .A2(G23), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G288), .B2(G16), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT33), .B(G1976), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT91), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n807), .A2(new_n805), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n808), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT92), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G24), .B(G290), .S(G16), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1986), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n712), .A2(G25), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n652), .A2(G131), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n476), .A2(G119), .ZN(new_n826));
  OR2_X1    g401(.A1(G95), .A2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(new_n712), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G1991), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT90), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n818), .B2(new_n819), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n820), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n820), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n800), .B1(new_n838), .B2(new_n840), .ZN(G311));
  INV_X1    g416(.A(G311), .ZN(G150));
  NAND4_X1  g417(.A1(new_n501), .A2(G93), .A3(new_n503), .A4(new_n510), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT103), .B(G55), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n539), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n503), .A2(G67), .A3(new_n500), .A4(new_n498), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n537), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n631), .A2(G559), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n555), .A3(new_n551), .ZN(new_n857));
  OAI221_X1 g432(.A(new_n846), .B1(new_n553), .B2(new_n554), .C1(new_n851), .C2(new_n852), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT104), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n856), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n866), .B2(KEYINPUT39), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n855), .B1(new_n867), .B2(new_n869), .ZN(G145));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  INV_X1    g446(.A(new_n491), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n487), .A2(KEYINPUT105), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n484), .B(new_n874), .C1(new_n483), .C2(new_n486), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n738), .A2(new_n773), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n738), .A2(new_n773), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n875), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n491), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n883), .A3(new_n877), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n753), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n476), .A2(G130), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n468), .A2(KEYINPUT107), .A3(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT107), .B1(new_n468), .B2(G118), .ZN(new_n891));
  OR2_X1    g466(.A1(G106), .A2(G2105), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(G2104), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G142), .ZN(new_n894));
  OAI221_X1 g469(.A(new_n889), .B1(new_n890), .B2(new_n893), .C1(new_n894), .C2(new_n469), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n649), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n829), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n898), .A2(KEYINPUT108), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n753), .A2(new_n886), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n880), .A2(new_n884), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n888), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT108), .A3(new_n898), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n657), .B(G160), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n481), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(KEYINPUT108), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n888), .A2(new_n899), .A3(new_n906), .A4(new_n901), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n903), .B2(new_n907), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(KEYINPUT109), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(KEYINPUT109), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n871), .B(new_n908), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(G395));
  AND3_X1   g489(.A1(new_n642), .A2(new_n644), .A3(new_n863), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n863), .B1(new_n642), .B2(new_n644), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n570), .A2(new_n574), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n630), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n628), .A2(new_n629), .ZN(new_n921));
  INV_X1    g496(.A(new_n625), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(KEYINPUT111), .A3(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n630), .A2(G299), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n630), .B2(G299), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n923), .A2(new_n918), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n917), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(G288), .B(G305), .Z(new_n935));
  XNOR2_X1  g510(.A(G290), .B(G166), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n920), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n920), .B2(new_n934), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n853), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(G868), .B2(new_n942), .ZN(G295));
  OAI21_X1  g518(.A(new_n941), .B1(G868), .B2(new_n942), .ZN(G331));
  NAND3_X1  g519(.A1(new_n584), .A2(G171), .A3(new_n590), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n584), .A2(KEYINPUT112), .A3(G171), .A4(new_n590), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n580), .A2(G168), .A3(new_n582), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n857), .A2(new_n861), .A3(new_n858), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n947), .A2(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT113), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n948), .A2(new_n949), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n945), .A2(new_n946), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(new_n860), .A3(new_n862), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n863), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n924), .A2(new_n927), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n925), .A2(KEYINPUT41), .ZN(new_n963));
  OAI22_X1  g538(.A1(KEYINPUT41), .A2(new_n919), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n947), .A2(new_n950), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n951), .A2(new_n952), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n919), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n953), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n937), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n954), .A2(new_n968), .A3(new_n960), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n953), .A2(new_n957), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n933), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n974), .A3(new_n937), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(new_n871), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n871), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n937), .B1(new_n972), .B2(new_n974), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n980), .A2(KEYINPUT43), .A3(new_n981), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n970), .B2(new_n980), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n970), .A2(new_n980), .A3(new_n985), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n983), .B1(new_n989), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g565(.A(KEYINPUT115), .B(G1384), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n883), .A2(KEYINPUT116), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n876), .B2(new_n991), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G160), .A2(G40), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n829), .B(new_n832), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n999), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n738), .A2(G1996), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n738), .A2(G1996), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n773), .B(G2067), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT117), .ZN(new_n1009));
  XNOR2_X1  g584(.A(G290), .B(G1986), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n1002), .B(new_n1009), .C1(new_n999), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT62), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n994), .B1(new_n876), .B2(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(G40), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n471), .A2(new_n474), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n487), .B2(new_n491), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1015), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n721), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1017), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n883), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2084), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1023), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G168), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1013), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT120), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1020), .A3(new_n1018), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1038), .B2(new_n721), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1039), .B2(G168), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1013), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1012), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT124), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(KEYINPUT62), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n606), .A2(new_n1052), .A3(new_n607), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n606), .A2(KEYINPUT118), .A3(new_n1052), .A4(new_n607), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G86), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n606), .B1(new_n1058), .B2(new_n511), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1055), .A2(new_n1056), .B1(G1981), .B2(new_n1059), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n883), .A2(new_n1027), .A3(new_n1017), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1066), .A2(G8), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1019), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n998), .B1(new_n994), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n803), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1024), .B1(new_n883), .B2(new_n1027), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1017), .B1(new_n1070), .B2(KEYINPUT50), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1073), .B1(new_n1078), .B2(G2090), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G8), .ZN(new_n1080));
  NAND3_X1  g655(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(G166), .B2(new_n1035), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1026), .B(new_n780), .C1(new_n1028), .C2(KEYINPUT50), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1073), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(G8), .A3(new_n1084), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n600), .A2(G1976), .A3(new_n601), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1067), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1067), .A2(new_n1091), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1068), .A2(new_n1086), .A3(new_n1089), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1026), .B(new_n1098), .C1(new_n1028), .C2(KEYINPUT50), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n876), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n1100), .B2(new_n1025), .ZN(new_n1101));
  INV_X1    g676(.A(G1961), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1072), .B2(G2078), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(G2078), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1103), .B(new_n1105), .C1(new_n1038), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G301), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1097), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1047), .A2(new_n1051), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n918), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n798), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1069), .A2(new_n1071), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1116), .A2(new_n1114), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1099), .A2(new_n1101), .A3(new_n792), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1066), .A2(G2067), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1130), .A2(new_n631), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1119), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT61), .B1(new_n1125), .B2(KEYINPUT123), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1134), .A3(new_n1119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n630), .A2(KEYINPUT82), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n630), .A2(KEYINPUT82), .ZN(new_n1139));
  OR3_X1    g714(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n631), .A2(KEYINPUT60), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(new_n1129), .A3(new_n1128), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n631), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1136), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT58), .B(G1341), .Z(new_n1145));
  NAND2_X1  g720(.A1(new_n1066), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1072), .B2(G1996), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n556), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1119), .A2(KEYINPUT61), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1127), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1132), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n473), .A2(KEYINPUT125), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n473), .A2(KEYINPUT125), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(G2105), .A3(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n471), .A2(new_n1016), .A3(new_n1107), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n997), .A2(new_n1069), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1103), .A2(new_n1157), .A3(new_n1105), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G171), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT54), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1110), .B(new_n1162), .C1(new_n1109), .C2(new_n1158), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1097), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1152), .A2(new_n1049), .A3(new_n1164), .A4(new_n1050), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1067), .ZN(new_n1167));
  NOR2_X1   g742(.A1(G288), .A2(G1976), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1067), .B1(new_n1064), .B2(KEYINPUT49), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1060), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1167), .B1(new_n1171), .B2(new_n1057), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1088), .A2(G8), .A3(new_n1084), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1173), .B(new_n1096), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1166), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1057), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1068), .B2(new_n1168), .ZN(new_n1178));
  OAI211_X1 g753(.A(KEYINPUT119), .B(new_n1174), .C1(new_n1178), .C2(new_n1167), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1032), .B(G8), .C1(new_n585), .C2(new_n591), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1084), .B1(new_n1088), .B2(G8), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1184), .A2(new_n1089), .A3(new_n1068), .A4(new_n1096), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1182), .B1(new_n1097), .B2(new_n1181), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1165), .A2(new_n1180), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1011), .B1(new_n1112), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1003), .A2(G1996), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT46), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n999), .B1(new_n738), .B2(new_n1006), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1192), .B(KEYINPUT126), .Z(new_n1193));
  NOR2_X1   g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1195));
  XNOR2_X1  g770(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n830), .A2(new_n832), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1009), .A2(new_n1197), .B1(G2067), .B2(new_n773), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1003), .A2(G1986), .A3(G290), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT48), .Z(new_n1201));
  AOI22_X1  g776(.A1(new_n1198), .A2(new_n999), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1196), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1189), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g779(.A1(new_n978), .A2(new_n982), .ZN(new_n1206));
  NOR4_X1   g780(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n1206), .A2(new_n912), .A3(new_n1207), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


