//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G137), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n196), .A2(new_n197), .B1(KEYINPUT64), .B2(new_n192), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n190), .A2(KEYINPUT11), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n193), .B1(new_n189), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n206), .A3(KEYINPUT65), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(G131), .C1(new_n194), .C2(new_n198), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT0), .A3(G128), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT0), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n211), .B(new_n213), .C1(new_n216), .C2(new_n217), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(new_n209), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n211), .A2(new_n213), .A3(new_n222), .A4(G128), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n212), .B2(G146), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n225), .A2(G128), .B1(new_n211), .B2(new_n213), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n189), .B2(new_n203), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n206), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT30), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT67), .A2(G119), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT67), .A2(G119), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n239), .B2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT2), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n247), .A3(new_n245), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT67), .A2(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT67), .A2(G119), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(G116), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n236), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n245), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n246), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT30), .B1(new_n221), .B2(new_n230), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n206), .A2(new_n229), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n206), .A2(new_n262), .A3(new_n229), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n263), .A3(new_n228), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT30), .A3(new_n221), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n234), .A2(new_n256), .A3(new_n259), .A4(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT27), .Z(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n269), .B(new_n270), .Z(new_n271));
  NAND3_X1  g085(.A1(new_n264), .A2(new_n255), .A3(new_n221), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n273));
  NAND4_X1  g087(.A1(new_n266), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n231), .A2(new_n256), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n282), .B2(new_n272), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n278), .B1(new_n272), .B2(new_n279), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n285), .B2(new_n271), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n272), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT28), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n264), .A2(new_n255), .A3(new_n221), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT72), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n292), .A3(new_n280), .ZN(new_n293));
  INV_X1    g107(.A(new_n271), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(KEYINPUT73), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n286), .A2(new_n288), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n276), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n293), .B2(new_n294), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n271), .B1(new_n266), .B2(new_n272), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT74), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n292), .A2(new_n280), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n255), .B1(new_n264), .B2(new_n221), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n291), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n264), .A2(new_n221), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n256), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n272), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT28), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n304), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n294), .A2(new_n300), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n303), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n302), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT32), .B(new_n187), .C1(new_n276), .C2(new_n296), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n299), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G210), .B1(G237), .B2(G902), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT86), .Z(new_n322));
  INV_X1    g136(.A(G104), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G107), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(G107), .ZN(new_n326));
  OAI21_X1  g140(.A(G101), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(new_n323), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n329));
  INV_X1    g143(.A(G107), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G104), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n331), .A3(new_n332), .A4(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n251), .A2(KEYINPUT5), .A3(new_n252), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n239), .A2(new_n337), .A3(G116), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(G113), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n247), .B1(new_n240), .B2(new_n245), .ZN(new_n340));
  AND4_X1   g154(.A1(new_n247), .A2(new_n251), .A3(new_n252), .A4(new_n245), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n335), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n328), .A2(new_n331), .A3(new_n324), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G101), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n346), .A3(G101), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n255), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G122), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n342), .B(new_n350), .C1(new_n255), .C2(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n220), .A2(G125), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(G125), .B2(new_n227), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G224), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n354), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G902), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n360), .A2(KEYINPUT7), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT85), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(KEYINPUT85), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n358), .A2(KEYINPUT85), .A3(new_n364), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n353), .A3(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n350), .B(KEYINPUT8), .Z(new_n371));
  OAI21_X1  g185(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n334), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n373), .B2(new_n342), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n363), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n322), .B1(new_n362), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n368), .A2(new_n353), .A3(new_n369), .ZN(new_n377));
  INV_X1    g191(.A(new_n374), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n354), .A2(new_n356), .A3(new_n361), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n321), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n383), .B(KEYINPUT84), .Z(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G113), .B(G122), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT90), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT89), .B(G104), .Z(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n359), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n212), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n210), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G140), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G125), .ZN(new_n404));
  INV_X1    g218(.A(G125), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT76), .A4(KEYINPUT16), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n405), .A2(KEYINPUT16), .A3(G140), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AND4_X1   g226(.A1(G146), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n407), .B2(new_n408), .ZN(new_n414));
  AOI21_X1  g228(.A(G146), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT88), .B1(new_n396), .B2(G131), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  AOI211_X1 g232(.A(new_n418), .B(new_n205), .C1(new_n394), .C2(new_n395), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT17), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  AND4_X1   g235(.A1(G143), .A2(new_n392), .A3(new_n359), .A4(G214), .ZN(new_n422));
  AOI21_X1  g236(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n423));
  OAI21_X1  g237(.A(G131), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n418), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n394), .A2(new_n205), .A3(new_n395), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT88), .B(G131), .C1(new_n422), .C2(new_n423), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n394), .A2(new_n429), .A3(new_n205), .A4(new_n395), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT17), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n391), .B(new_n402), .C1(new_n421), .C2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n409), .A2(G146), .A3(new_n410), .A4(new_n412), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n398), .B(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n436), .B2(G146), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n417), .A2(new_n419), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n427), .A2(new_n430), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n402), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n390), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n433), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G475), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT20), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n433), .A2(new_n442), .A3(KEYINPUT91), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT91), .B1(new_n433), .B2(new_n442), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n448), .A2(new_n449), .A3(new_n445), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n210), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n434), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n425), .B2(new_n428), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n439), .A2(new_n438), .A3(new_n456), .ZN(new_n459));
  AOI211_X1 g273(.A(new_n441), .B(new_n390), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n416), .B(new_n420), .C1(KEYINPUT17), .C2(new_n431), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n391), .B1(new_n461), .B2(new_n402), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n363), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT92), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n363), .C1(new_n460), .C2(new_n462), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(G475), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(G234), .A2(G237), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(G902), .A3(G953), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n469), .B(KEYINPUT93), .Z(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(G898), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n359), .A2(G952), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(G234), .B2(G237), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G478), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G116), .ZN(new_n480));
  INV_X1    g294(.A(G116), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G122), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n330), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n212), .A2(G128), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT13), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n217), .A2(G143), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n485), .A2(new_n486), .ZN(new_n490));
  OAI21_X1  g304(.A(G134), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n485), .A2(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n188), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n188), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n483), .A2(new_n330), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n480), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G107), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT9), .B(G234), .ZN(new_n502));
  INV_X1    g316(.A(G217), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n502), .A2(new_n503), .A3(G953), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n494), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n494), .B2(new_n501), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n478), .B1(new_n507), .B2(G902), .ZN(new_n508));
  OAI221_X1 g322(.A(new_n363), .B1(KEYINPUT15), .B2(new_n477), .C1(new_n505), .C2(new_n506), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n452), .A2(new_n467), .A3(new_n476), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G221), .B1(new_n502), .B2(G902), .ZN(new_n513));
  INV_X1    g327(.A(G469), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT12), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n227), .A2(new_n334), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n333), .B(new_n327), .C1(new_n224), .C2(new_n226), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n207), .A2(new_n209), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n207), .A2(new_n209), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(KEYINPUT12), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n345), .A2(new_n220), .A3(new_n347), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT81), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n345), .A2(new_n220), .A3(KEYINPUT81), .A4(new_n347), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT82), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT10), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(KEYINPUT10), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n517), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n517), .B2(new_n531), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(new_n535), .A3(new_n519), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n524), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G140), .ZN(new_n538));
  INV_X1    g352(.A(G227), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n529), .A2(new_n535), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n521), .ZN(new_n544));
  INV_X1    g358(.A(new_n541), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n536), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n514), .B1(new_n547), .B2(new_n363), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n529), .A2(new_n535), .A3(new_n519), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n519), .B1(new_n529), .B2(new_n535), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n541), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n524), .A2(new_n536), .A3(new_n545), .ZN(new_n552));
  AOI211_X1 g366(.A(G469), .B(G902), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n513), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT83), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n545), .B1(new_n544), .B2(new_n536), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n524), .A2(new_n536), .A3(new_n545), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n514), .B(new_n363), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(G469), .A2(G902), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n559), .C1(new_n514), .C2(new_n547), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n513), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n386), .B(new_n512), .C1(new_n555), .C2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G128), .B1(new_n237), .B2(new_n238), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n235), .A2(new_n217), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT23), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n217), .B1(new_n237), .B2(new_n238), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT24), .B(G110), .Z(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(new_n565), .ZN(new_n572));
  OAI22_X1  g386(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n398), .A2(new_n210), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n573), .A2(new_n434), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT77), .B1(new_n416), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n455), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n575), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n584), .B(new_n585), .Z(new_n586));
  OAI21_X1  g400(.A(KEYINPUT78), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n573), .A2(new_n434), .A3(new_n574), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n455), .A2(new_n580), .A3(new_n581), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n580), .B1(new_n455), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(new_n586), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n588), .B(new_n586), .C1(new_n589), .C2(new_n590), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n579), .A2(new_n582), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n588), .A4(new_n586), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n587), .A2(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n503), .B1(G234), .B2(new_n363), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(G902), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT80), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n597), .A2(new_n599), .ZN(new_n605));
  AND4_X1   g419(.A1(KEYINPUT80), .A2(new_n604), .A3(new_n605), .A4(new_n602), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n605), .A3(new_n363), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT25), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT25), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n604), .A2(new_n605), .A3(new_n610), .A4(new_n363), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n611), .A3(new_n601), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n320), .A2(new_n563), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  OAI21_X1  g430(.A(new_n363), .B1(new_n276), .B2(new_n296), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(G472), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n274), .B(KEYINPUT71), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n285), .A2(new_n277), .A3(new_n271), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT73), .B1(new_n293), .B2(new_n294), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n623), .A3(new_n288), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n618), .A2(G472), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n363), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n613), .B1(new_n562), .B2(new_n555), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n379), .A2(new_n321), .A3(new_n380), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n321), .B1(new_n379), .B2(new_n380), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n384), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n476), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n477), .A2(new_n363), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n477), .B(new_n363), .C1(new_n505), .C2(new_n506), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n494), .A2(new_n501), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT33), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n505), .B2(new_n506), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n507), .A2(KEYINPUT33), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n637), .B(new_n639), .C1(new_n646), .C2(G478), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n464), .A2(G475), .A3(new_n466), .ZN(new_n648));
  INV_X1    g462(.A(new_n447), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n443), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n433), .A2(new_n442), .A3(KEYINPUT91), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n444), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n649), .B1(new_n653), .B2(KEYINPUT20), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n647), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n639), .A2(new_n637), .ZN(new_n658));
  INV_X1    g472(.A(new_n646), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(new_n477), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n452), .B2(new_n467), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT96), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n636), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n631), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NOR2_X1   g480(.A1(new_n448), .A2(new_n449), .ZN(new_n667));
  AOI22_X1  g481(.A1(KEYINPUT20), .A2(new_n653), .B1(new_n667), .B2(new_n446), .ZN(new_n668));
  OR3_X1    g482(.A1(new_n668), .A2(new_n648), .A3(new_n511), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n476), .B(KEYINPUT97), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n669), .A2(new_n384), .A3(new_n634), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n631), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  AOI21_X1  g488(.A(new_n386), .B1(new_n555), .B2(new_n562), .ZN(new_n675));
  INV_X1    g489(.A(new_n601), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n608), .B2(KEYINPUT25), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n583), .B(new_n678), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n677), .A2(new_n611), .B1(new_n602), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n512), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n619), .A2(new_n675), .A3(new_n626), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  AOI21_X1  g498(.A(new_n680), .B1(new_n562), .B2(new_n555), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n474), .B1(new_n470), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT98), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n669), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n320), .A2(new_n635), .A3(new_n685), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  AND2_X1   g505(.A1(new_n266), .A2(new_n272), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n294), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n363), .B1(new_n310), .B2(new_n271), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n299), .A2(new_n319), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT99), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n680), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n555), .A2(new_n562), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n688), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT40), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n382), .B(KEYINPUT38), .Z(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n452), .A2(new_n467), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n510), .A4(new_n385), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n698), .A2(new_n699), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  INV_X1    g526(.A(new_n688), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n647), .B(new_n713), .C1(new_n648), .C2(new_n654), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n706), .A2(KEYINPUT101), .A3(new_n647), .A4(new_n713), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n635), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT102), .A4(new_n635), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n320), .A3(new_n685), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n558), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n551), .A2(new_n552), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n514), .B1(new_n726), .B2(new_n363), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n725), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n513), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n320), .A2(new_n663), .A3(new_n614), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT104), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND4_X1  g548(.A1(new_n320), .A2(new_n671), .A3(new_n614), .A4(new_n730), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AND3_X1   g550(.A1(new_n728), .A2(new_n513), .A3(new_n635), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n320), .A2(new_n681), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  OAI21_X1  g553(.A(new_n288), .B1(new_n313), .B2(new_n271), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n288), .B(KEYINPUT105), .C1(new_n313), .C2(new_n271), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n620), .A3(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n744), .A2(new_n187), .B1(new_n617), .B2(G472), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n648), .A2(new_n654), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n747), .B2(new_n511), .ZN(new_n748));
  INV_X1    g562(.A(new_n670), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n706), .A2(KEYINPUT106), .A3(new_n510), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n751), .A3(new_n737), .A4(new_n614), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  AND2_X1   g567(.A1(new_n716), .A2(new_n717), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n745), .A2(new_n737), .A3(new_n754), .A4(new_n699), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT32), .B1(new_n624), .B2(new_n187), .ZN(new_n758));
  INV_X1    g572(.A(new_n319), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n299), .A2(KEYINPUT108), .A3(new_n319), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n318), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n513), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n560), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n382), .A2(new_n384), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n548), .A2(new_n553), .A3(new_n764), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n762), .A2(new_n614), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n320), .A2(new_n614), .A3(new_n754), .A4(new_n768), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT109), .B(G131), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G33));
  NAND4_X1  g590(.A1(new_n320), .A2(new_n614), .A3(new_n689), .A4(new_n768), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n747), .A2(new_n647), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT43), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n628), .A2(new_n680), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT44), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n514), .B1(new_n547), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n784), .B2(new_n547), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT46), .B1(new_n786), .B2(new_n559), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n553), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n559), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n763), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n701), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n782), .A2(new_n766), .A3(new_n783), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  XOR2_X1   g608(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n795));
  AOI211_X1 g609(.A(new_n763), .B(new_n795), .C1(new_n788), .C2(new_n789), .ZN(new_n796));
  NOR2_X1   g610(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n754), .A2(new_n613), .A3(new_n766), .ZN(new_n799));
  OR4_X1    g613(.A1(new_n320), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  AND2_X1   g615(.A1(new_n762), .A2(new_n614), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n730), .A2(KEYINPUT115), .A3(new_n766), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  INV_X1    g618(.A(new_n766), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n729), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n474), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n780), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT48), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n807), .A2(new_n613), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n662), .A2(new_n657), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n698), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n780), .A2(new_n475), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(new_n614), .A3(new_n745), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(KEYINPUT118), .A3(new_n737), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT118), .B1(new_n815), .B2(new_n737), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n473), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n810), .A2(new_n813), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n705), .A2(new_n729), .A3(new_n385), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n808), .A2(new_n699), .A3(new_n745), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n728), .B(KEYINPUT112), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n763), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n798), .B2(new_n796), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n766), .A3(new_n815), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n811), .A2(new_n698), .A3(new_n747), .A4(new_n660), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n819), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n833), .B2(new_n834), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT117), .B1(new_n840), .B2(KEYINPUT51), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n836), .A2(new_n842), .A3(new_n837), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n838), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n748), .A2(new_n635), .A3(new_n750), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n680), .A2(new_n765), .A3(new_n713), .A4(new_n767), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n696), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n722), .A2(new_n690), .A3(new_n755), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT52), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n467), .A2(new_n511), .A3(new_n713), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n805), .A2(new_n668), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n320), .A2(new_n685), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n745), .A2(new_n754), .A3(new_n699), .A4(new_n768), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n777), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n322), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n379), .B2(new_n380), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n385), .B(new_n749), .C1(new_n632), .C2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT113), .B1(new_n655), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n384), .B(new_n670), .C1(new_n376), .C2(new_n381), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n661), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n747), .A3(new_n510), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n629), .A3(new_n626), .A4(new_n619), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n615), .A2(new_n867), .A3(new_n682), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n857), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n735), .A2(new_n752), .A3(new_n738), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n732), .A2(new_n774), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n846), .B1(new_n852), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n774), .A2(new_n869), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n690), .A2(new_n755), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n722), .A4(new_n850), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n851), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n874), .A2(new_n879), .A3(KEYINPUT53), .A4(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n873), .A2(KEYINPUT54), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT54), .B1(new_n873), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n845), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n873), .A2(new_n883), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n873), .A2(KEYINPUT54), .A3(new_n883), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT114), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n844), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n827), .B(KEYINPUT49), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n613), .A2(new_n779), .A3(new_n763), .A4(new_n384), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT111), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n698), .A2(new_n704), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n359), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n363), .B1(new_n873), .B2(new_n883), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n354), .A2(new_n356), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n361), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n362), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n322), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT119), .Z(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n909), .B2(new_n911), .ZN(G51));
  NOR2_X1   g726(.A1(new_n884), .A2(new_n885), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n559), .B(KEYINPUT57), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n726), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n901), .B(new_n785), .C1(new_n784), .C2(new_n547), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n899), .B1(new_n916), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  INV_X1    g733(.A(new_n667), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n899), .B1(new_n919), .B2(new_n920), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G60));
  NAND2_X1  g740(.A1(new_n886), .A2(new_n891), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n637), .B(KEYINPUT59), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n659), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n646), .A2(new_n928), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n899), .B1(new_n913), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT121), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n928), .B1(new_n886), .B2(new_n891), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n932), .B(new_n935), .C1(new_n936), .C2(new_n659), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT122), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n887), .A2(new_n679), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n887), .A2(new_n941), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n900), .B(new_n942), .C1(new_n943), .C2(new_n600), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g759(.A1(G224), .A2(G953), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n471), .A2(new_n946), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n868), .B(new_n870), .C1(new_n880), .C2(new_n881), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n359), .ZN(new_n949));
  INV_X1    g763(.A(G898), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n903), .B1(new_n950), .B2(G953), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n949), .B(new_n951), .Z(G69));
  NAND2_X1  g766(.A1(new_n875), .A2(new_n722), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT124), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n711), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n234), .A2(new_n259), .A3(new_n265), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT123), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n436), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n711), .A2(new_n961), .A3(new_n954), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n661), .B1(new_n747), .B2(new_n510), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n702), .A2(new_n805), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n320), .A3(new_n614), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n793), .A2(new_n800), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n956), .A2(new_n960), .A3(new_n962), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n954), .A2(new_n793), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n802), .A2(new_n792), .A3(new_n848), .ZN(new_n971));
  AND4_X1   g785(.A1(new_n774), .A2(new_n971), .A3(new_n800), .A4(new_n777), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n968), .B1(new_n973), .B2(new_n960), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n959), .A2(G227), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n686), .B(new_n359), .C1(new_n960), .C2(new_n539), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n974), .A2(new_n359), .B1(new_n975), .B2(new_n976), .ZN(G72));
  NAND4_X1  g791(.A1(new_n956), .A2(new_n962), .A3(new_n948), .A4(new_n967), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AOI211_X1 g794(.A(new_n294), .B(new_n692), .C1(new_n978), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n692), .A2(new_n294), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n970), .A2(new_n948), .A3(new_n972), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n980), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n302), .B(KEYINPUT127), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n287), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n887), .A2(new_n980), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n900), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n981), .A2(new_n984), .A3(new_n988), .ZN(G57));
endmodule


