

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U322 ( .A(n571), .B(KEYINPUT41), .Z(n550) );
  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n425) );
  XNOR2_X1 U324 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n419) );
  XNOR2_X1 U325 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U326 ( .A(n420), .B(n419), .ZN(n421) );
  NOR2_X1 U327 ( .A1(n529), .A2(n445), .ZN(n560) );
  XNOR2_X1 U328 ( .A(n446), .B(G176GAT), .ZN(n447) );
  XNOR2_X1 U329 ( .A(n448), .B(n447), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n291) );
  XNOR2_X1 U331 ( .A(G134GAT), .B(KEYINPUT81), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U333 ( .A(n292), .B(G127GAT), .Z(n294) );
  XNOR2_X1 U334 ( .A(G113GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n327) );
  XOR2_X1 U336 ( .A(G99GAT), .B(G190GAT), .Z(n296) );
  XNOR2_X1 U337 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U339 ( .A(n327), .B(n297), .Z(n299) );
  NAND2_X1 U340 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U342 ( .A(G176GAT), .B(G183GAT), .Z(n301) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G15GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U345 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U346 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n305) );
  XNOR2_X1 U347 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(n306), .ZN(n338) );
  XOR2_X1 U350 ( .A(KEYINPUT86), .B(KEYINPUT66), .Z(n308) );
  XNOR2_X1 U351 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U353 ( .A(n338), .B(n309), .Z(n310) );
  XOR2_X1 U354 ( .A(n311), .B(n310), .Z(n493) );
  INV_X1 U355 ( .A(n493), .ZN(n529) );
  NAND2_X1 U356 ( .A1(G233GAT), .A2(G225GAT), .ZN(n317) );
  XOR2_X1 U357 ( .A(KEYINPUT1), .B(G57GAT), .Z(n313) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(G1GAT), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n315) );
  XOR2_X1 U360 ( .A(G162GAT), .B(G85GAT), .Z(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n325) );
  XOR2_X1 U363 ( .A(G148GAT), .B(KEYINPUT6), .Z(n323) );
  XOR2_X1 U364 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n319) );
  XNOR2_X1 U365 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n321) );
  XNOR2_X1 U367 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n320), .B(KEYINPUT2), .ZN(n433) );
  XNOR2_X1 U369 ( .A(n321), .B(n433), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U371 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U372 ( .A(n327), .B(n326), .Z(n514) );
  INV_X1 U373 ( .A(n514), .ZN(n487) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G204GAT), .Z(n329) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(G92GAT), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n329), .B(n328), .ZN(n342) );
  XOR2_X1 U377 ( .A(KEYINPUT90), .B(n342), .Z(n331) );
  NAND2_X1 U378 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U380 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n333) );
  XNOR2_X1 U381 ( .A(G218GAT), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U383 ( .A(G197GAT), .B(n334), .Z(n432) );
  XOR2_X1 U384 ( .A(n335), .B(n432), .Z(n337) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .Z(n358) );
  XOR2_X1 U386 ( .A(G8GAT), .B(G183GAT), .Z(n380) );
  XNOR2_X1 U387 ( .A(n358), .B(n380), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n340) );
  INV_X1 U389 ( .A(n338), .ZN(n339) );
  XOR2_X1 U390 ( .A(n340), .B(n339), .Z(n516) );
  INV_X1 U391 ( .A(n516), .ZN(n491) );
  XOR2_X1 U392 ( .A(KEYINPUT121), .B(n491), .Z(n424) );
  XOR2_X1 U393 ( .A(G99GAT), .B(G85GAT), .Z(n341) );
  XOR2_X1 U394 ( .A(KEYINPUT74), .B(n341), .Z(n371) );
  XOR2_X1 U395 ( .A(n342), .B(n371), .Z(n355) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(G78GAT), .Z(n344) );
  XNOR2_X1 U397 ( .A(G148GAT), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n438) );
  XNOR2_X1 U399 ( .A(G71GAT), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n345), .B(KEYINPUT13), .ZN(n388) );
  XNOR2_X1 U401 ( .A(n438), .B(n388), .ZN(n353) );
  XNOR2_X1 U402 ( .A(KEYINPUT72), .B(KEYINPUT75), .ZN(n347) );
  XNOR2_X1 U403 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U405 ( .A(KEYINPUT33), .B(G120GAT), .Z(n349) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n571) );
  XOR2_X1 U411 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n357) );
  XNOR2_X1 U412 ( .A(G92GAT), .B(G106GAT), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U414 ( .A(KEYINPUT65), .B(G218GAT), .Z(n360) );
  XOR2_X1 U415 ( .A(G50GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U416 ( .A(n358), .B(n436), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U418 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n366) );
  XNOR2_X1 U422 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n374) );
  XOR2_X1 U425 ( .A(G29GAT), .B(G43GAT), .Z(n370) );
  XNOR2_X1 U426 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n398) );
  INV_X1 U428 ( .A(n371), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n398), .B(n372), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n412) );
  XOR2_X1 U431 ( .A(KEYINPUT36), .B(n412), .Z(n581) );
  XOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n376) );
  XNOR2_X1 U433 ( .A(G22GAT), .B(G78GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n392) );
  XOR2_X1 U435 ( .A(G211GAT), .B(G64GAT), .Z(n378) );
  XNOR2_X1 U436 ( .A(G127GAT), .B(G155GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U438 ( .A(n380), .B(n379), .Z(n382) );
  NAND2_X1 U439 ( .A1(G231GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n384) );
  XNOR2_X1 U442 ( .A(KEYINPUT78), .B(KEYINPUT14), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n390) );
  XNOR2_X1 U445 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n387), .B(G15GAT), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n395), .B(n388), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n451) );
  NOR2_X1 U450 ( .A1(n581), .A2(n451), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT45), .B(n393), .Z(n394) );
  NOR2_X1 U452 ( .A1(n571), .A2(n394), .ZN(n411) );
  XOR2_X1 U453 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XOR2_X1 U454 ( .A(n439), .B(n395), .Z(n397) );
  XNOR2_X1 U455 ( .A(G36GAT), .B(G50GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n402) );
  XOR2_X1 U457 ( .A(n398), .B(KEYINPUT70), .Z(n400) );
  NAND2_X1 U458 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n410) );
  XOR2_X1 U461 ( .A(G8GAT), .B(G197GAT), .Z(n404) );
  XNOR2_X1 U462 ( .A(G169GAT), .B(G113GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U464 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n499) );
  NAND2_X1 U469 ( .A1(n411), .A2(n499), .ZN(n422) );
  INV_X1 U470 ( .A(n412), .ZN(n413) );
  INV_X1 U471 ( .A(n413), .ZN(n559) );
  INV_X1 U472 ( .A(n499), .ZN(n566) );
  NAND2_X1 U473 ( .A1(n566), .A2(n550), .ZN(n415) );
  INV_X1 U474 ( .A(KEYINPUT46), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  INV_X1 U476 ( .A(n451), .ZN(n575) );
  NOR2_X1 U477 ( .A1(n416), .A2(n575), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n417), .B(KEYINPUT111), .ZN(n418) );
  NOR2_X1 U479 ( .A1(n559), .A2(n418), .ZN(n420) );
  NAND2_X1 U480 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n423), .B(KEYINPUT48), .ZN(n526) );
  NAND2_X1 U482 ( .A1(n424), .A2(n526), .ZN(n426) );
  NOR2_X1 U483 ( .A1(n487), .A2(n427), .ZN(n428) );
  XOR2_X1 U484 ( .A(KEYINPUT64), .B(n428), .Z(n564) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n430) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT87), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n443) );
  XOR2_X1 U489 ( .A(n433), .B(KEYINPUT22), .Z(n435) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U492 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n462) );
  NOR2_X1 U496 ( .A1(n564), .A2(n462), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n444), .B(KEYINPUT55), .ZN(n445) );
  NAND2_X1 U498 ( .A1(n560), .A2(n550), .ZN(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n446) );
  XOR2_X1 U500 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n450) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n472) );
  NOR2_X1 U503 ( .A1(n499), .A2(n571), .ZN(n484) );
  NOR2_X1 U504 ( .A1(n559), .A2(n451), .ZN(n452) );
  XNOR2_X1 U505 ( .A(KEYINPUT16), .B(n452), .ZN(n470) );
  NOR2_X1 U506 ( .A1(n529), .A2(n516), .ZN(n453) );
  NOR2_X1 U507 ( .A1(n462), .A2(n453), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT25), .ZN(n459) );
  XOR2_X1 U509 ( .A(n491), .B(KEYINPUT91), .Z(n455) );
  XNOR2_X1 U510 ( .A(n455), .B(KEYINPUT27), .ZN(n464) );
  NAND2_X1 U511 ( .A1(n462), .A2(n529), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n456), .B(KEYINPUT26), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT94), .B(n457), .Z(n543) );
  NAND2_X1 U514 ( .A1(n464), .A2(n543), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n514), .A2(n460), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT95), .B(n461), .Z(n469) );
  XOR2_X1 U518 ( .A(n462), .B(KEYINPUT67), .Z(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT28), .B(n463), .Z(n522) );
  NAND2_X1 U520 ( .A1(n487), .A2(n464), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT92), .B(n465), .Z(n527) );
  NAND2_X1 U522 ( .A1(n522), .A2(n527), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT93), .B(n466), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n467), .A2(n529), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n482) );
  AND2_X1 U526 ( .A1(n470), .A2(n482), .ZN(n501) );
  NAND2_X1 U527 ( .A1(n484), .A2(n501), .ZN(n477) );
  NOR2_X1 U528 ( .A1(n514), .A2(n477), .ZN(n471) );
  XOR2_X1 U529 ( .A(n472), .B(n471), .Z(G1324GAT) );
  NOR2_X1 U530 ( .A1(n516), .A2(n477), .ZN(n473) );
  XOR2_X1 U531 ( .A(G8GAT), .B(n473), .Z(G1325GAT) );
  NOR2_X1 U532 ( .A1(n529), .A2(n477), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G15GAT), .B(n476), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n522), .A2(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n480), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n489) );
  NOR2_X1 U541 ( .A1(n581), .A2(n575), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n483), .ZN(n513) );
  NAND2_X1 U544 ( .A1(n513), .A2(n484), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n496) );
  NAND2_X1 U547 ( .A1(n496), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U549 ( .A(G29GAT), .B(n490), .Z(G1328GAT) );
  NAND2_X1 U550 ( .A1(n491), .A2(n496), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U552 ( .A1(n493), .A2(n496), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U555 ( .A(G50GAT), .B(KEYINPUT103), .Z(n498) );
  INV_X1 U556 ( .A(n522), .ZN(n532) );
  NAND2_X1 U557 ( .A1(n496), .A2(n532), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  NAND2_X1 U559 ( .A1(n550), .A2(n499), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n500), .Z(n512) );
  NAND2_X1 U561 ( .A1(n501), .A2(n512), .ZN(n508) );
  NOR2_X1 U562 ( .A1(n514), .A2(n508), .ZN(n503) );
  XNOR2_X1 U563 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n516), .A2(n508), .ZN(n505) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n529), .A2(n508), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(n506), .Z(n507) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n522), .A2(n508), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n512), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n514), .A2(n521), .ZN(n515) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n521), .ZN(n517) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(n517), .Z(n518) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n529), .A2(n521), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NAND2_X1 U588 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U589 ( .A(KEYINPUT113), .B(n528), .Z(n544) );
  NOR2_X1 U590 ( .A1(n529), .A2(n544), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT114), .B(n530), .Z(n531) );
  NOR2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n566), .A2(n539), .ZN(n533) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U596 ( .A1(n539), .A2(n550), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  NAND2_X1 U599 ( .A1(n539), .A2(n575), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U603 ( .A1(n539), .A2(n559), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT117), .Z(n546) );
  INV_X1 U607 ( .A(n543), .ZN(n563) );
  NOR2_X1 U608 ( .A1(n563), .A2(n544), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n555), .A2(n566), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n548) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U614 ( .A(KEYINPUT52), .B(n549), .Z(n552) );
  NAND2_X1 U615 ( .A1(n555), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n555), .A2(n575), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n559), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n566), .A2(n560), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n575), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT58), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(n562), .ZN(G1351GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT123), .B(n565), .ZN(n580) );
  INV_X1 U631 ( .A(n580), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n576), .A2(n566), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U638 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

