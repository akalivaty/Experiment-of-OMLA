//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n212));
  OR2_X1    g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT24), .A3(new_n211), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n205), .A2(new_n208), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n219), .A2(new_n212), .A3(new_n214), .A4(new_n216), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n226), .C1(new_n229), .C2(new_n225), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n231), .B(new_n227), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n227), .A2(new_n231), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n206), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n204), .A2(new_n240), .A3(new_n210), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n245));
  AOI21_X1  g044(.A(G190gat), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n243), .B1(new_n246), .B2(new_n236), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n234), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n234), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n218), .A2(new_n220), .B1(KEYINPUT64), .B2(KEYINPUT25), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n237), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n242), .B1(new_n252), .B2(KEYINPUT28), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G227gat), .ZN(new_n256));
  INV_X1    g055(.A(G233gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(KEYINPUT32), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G15gat), .B(G43gat), .Z(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n258), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n248), .B2(new_n254), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT32), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(KEYINPUT33), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT68), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272));
  INV_X1    g071(.A(new_n270), .ZN(new_n273));
  NOR4_X1   g072(.A1(new_n267), .A2(new_n272), .A3(new_n268), .A4(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n265), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT34), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n255), .B2(new_n258), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n248), .A2(new_n254), .A3(KEYINPUT34), .A4(new_n266), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n280), .B(new_n265), .C1(new_n271), .C2(new_n274), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT31), .B(G50gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(G141gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(G141gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n288), .A2(G148gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n299), .B2(new_n300), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n293), .B1(new_n296), .B2(KEYINPUT2), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n298), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT73), .B1(new_n289), .B2(new_n291), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n298), .A3(new_n305), .A4(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n297), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G197gat), .B(G204gat), .ZN(new_n312));
  INV_X1    g111(.A(G211gat), .ZN(new_n313));
  INV_X1    g112(.A(G218gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(KEYINPUT22), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT79), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n311), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n297), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n305), .A3(new_n308), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n328), .B2(new_n309), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT80), .B1(new_n332), .B2(new_n319), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n331), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n319), .B1(new_n334), .B2(new_n320), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n325), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G228gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(new_n257), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n330), .B1(new_n319), .B2(new_n320), .ZN(new_n342));
  OAI22_X1  g141(.A1(new_n342), .A2(new_n329), .B1(new_n339), .B2(new_n257), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(new_n335), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n286), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n285), .B(new_n344), .C1(new_n338), .C2(new_n340), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  INV_X1    g149(.A(G22gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT81), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n353), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n346), .B2(new_n348), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n284), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n334), .B(new_n249), .C1(new_n322), .C2(new_n329), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n329), .A2(KEYINPUT4), .A3(new_n234), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n329), .A2(new_n234), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT77), .B1(new_n329), .B2(new_n234), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n311), .A2(new_n249), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n364), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n311), .A2(new_n249), .A3(KEYINPUT77), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n379), .A3(KEYINPUT5), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n370), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n363), .B(new_n383), .C1(new_n366), .C2(new_n367), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n384), .A2(KEYINPUT5), .A3(new_n374), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n362), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n380), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n379), .B1(new_n376), .B2(KEYINPUT5), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n369), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n385), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n361), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n361), .B1(new_n389), .B2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT6), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n223), .A2(new_n247), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT71), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n250), .A2(new_n253), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT29), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n402), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n319), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n398), .A2(new_n401), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n407), .A2(new_n402), .B1(new_n397), .B2(new_n403), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(new_n319), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  INV_X1    g209(.A(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT72), .B(G64gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n406), .B(new_n414), .C1(new_n408), .C2(new_n319), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT30), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n409), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n357), .A2(KEYINPUT35), .A3(new_n396), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n393), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n386), .A2(new_n391), .A3(KEYINPUT82), .A4(new_n392), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n395), .ZN(new_n428));
  INV_X1    g227(.A(new_n279), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n275), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n275), .A2(new_n429), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n430), .A2(new_n354), .A3(new_n356), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(new_n433), .A3(new_n421), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT35), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n423), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n415), .B1(new_n409), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n437), .B2(new_n409), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n439), .A2(KEYINPUT38), .B1(new_n409), .B2(new_n415), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT38), .ZN(new_n441));
  OR3_X1    g240(.A1(new_n408), .A2(KEYINPUT83), .A3(new_n318), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n404), .A2(new_n318), .A3(new_n405), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT83), .B1(new_n408), .B2(new_n318), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n441), .B(new_n438), .C1(new_n445), .C2(new_n437), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n427), .A2(new_n395), .A3(new_n440), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n354), .A2(new_n356), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n384), .A2(new_n374), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n373), .A2(new_n375), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n449), .B(KEYINPUT39), .C1(new_n374), .C2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(new_n361), .C1(KEYINPUT39), .C2(new_n449), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n454), .A2(new_n455), .A3(new_n394), .ZN(new_n456));
  INV_X1    g255(.A(new_n421), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n396), .A2(new_n421), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n448), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n284), .A2(KEYINPUT36), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n430), .B2(new_n431), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n459), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n436), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n469));
  INV_X1    g268(.A(G15gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n351), .ZN(new_n471));
  NAND2_X1  g270(.A1(G15gat), .A2(G22gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G1gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT16), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n474), .A3(new_n472), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G8gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n477), .B2(KEYINPUT87), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n476), .B(new_n477), .C1(KEYINPUT87), .C2(new_n479), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G64gat), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT92), .B1(new_n489), .B2(G57gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491));
  INV_X1    g290(.A(G57gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(G64gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n490), .B(new_n493), .C1(new_n492), .C2(G64gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(G71gat), .B(G78gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT9), .ZN(new_n496));
  INV_X1    g295(.A(G71gat), .ZN(new_n497));
  INV_X1    g296(.A(G78gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n495), .ZN(new_n501));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n501), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n488), .B1(KEYINPUT21), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G183gat), .ZN(new_n506));
  AND2_X1   g305(.A1(G231gat), .A2(G233gat), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n469), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  INV_X1    g311(.A(new_n469), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n504), .A2(KEYINPUT21), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n313), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n515), .B(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G127gat), .B(G155gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n510), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n510), .B2(new_n514), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524));
  INV_X1    g323(.A(G43gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(G50gat), .ZN(new_n526));
  INV_X1    g325(.A(G50gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(G43gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(G43gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(G50gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT15), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT85), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n542), .A2(new_n532), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n542), .A2(new_n544), .A3(new_n529), .A4(new_n532), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n541), .A2(new_n543), .A3(new_n549), .A4(new_n545), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(KEYINPUT17), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G99gat), .B(G106gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT95), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(G99gat), .A3(G106gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT8), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n411), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n556), .B(new_n558), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n558), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  INV_X1    g369(.A(new_n556), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n547), .A2(new_n550), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G134gat), .B(G162gat), .Z(new_n581));
  AOI21_X1  g380(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n580), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n523), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n483), .B1(new_n551), .B2(new_n552), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n487), .B1(new_n547), .B2(new_n550), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n589), .B(KEYINPUT13), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n488), .A2(new_n575), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n487), .A2(new_n547), .A3(new_n550), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n592), .B2(KEYINPUT18), .ZN(new_n599));
  INV_X1    g398(.A(new_n483), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n553), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n589), .A3(new_n596), .ZN(new_n602));
  INV_X1    g401(.A(new_n593), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT90), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n594), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n606));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G113gat), .B(G141gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT91), .B1(new_n592), .B2(new_n593), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n602), .A2(new_n615), .A3(new_n603), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n614), .A2(new_n599), .A3(new_n616), .A4(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n586), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n563), .A2(new_n566), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT96), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n556), .B1(new_n625), .B2(new_n558), .ZN(new_n626));
  INV_X1    g425(.A(new_n569), .ZN(new_n627));
  OAI211_X1 g426(.A(KEYINPUT10), .B(new_n504), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n576), .A2(KEYINPUT99), .A3(KEYINPUT10), .A4(new_n504), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n500), .A2(new_n633), .A3(new_n503), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n500), .B2(new_n503), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n576), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n572), .A2(new_n633), .A3(new_n504), .A4(new_n569), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT10), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n621), .B1(new_n632), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n634), .B(new_n636), .C1(new_n572), .C2(new_n569), .ZN(new_n643));
  AND4_X1   g442(.A1(new_n633), .A2(new_n572), .A3(new_n504), .A4(new_n569), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n645), .A2(KEYINPUT100), .A3(new_n630), .A4(new_n631), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n638), .A2(new_n649), .A3(new_n639), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n648), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n632), .A2(new_n640), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n656), .B2(new_n649), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT101), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(KEYINPUT101), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n468), .A2(new_n620), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n396), .A2(KEYINPUT102), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n393), .A2(new_n666), .A3(new_n395), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n474), .ZN(G1324gat));
  NAND4_X1  g470(.A1(new_n468), .A2(new_n620), .A3(new_n457), .A4(new_n663), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT16), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n479), .ZN(new_n674));
  NOR2_X1   g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR4_X1   g477(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n674), .A4(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n672), .A2(G8gat), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT103), .B1(new_n672), .B2(G8gat), .ZN(new_n683));
  OAI22_X1  g482(.A1(new_n678), .A2(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686));
  OAI221_X1 g485(.A(new_n686), .B1(new_n682), .B2(new_n683), .C1(new_n678), .C2(new_n679), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1325gat));
  INV_X1    g487(.A(new_n430), .ZN(new_n689));
  INV_X1    g488(.A(new_n431), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n470), .B1(new_n664), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT105), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n466), .A2(KEYINPUT106), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n664), .A2(new_n470), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n699), .ZN(G1326gat));
  INV_X1    g499(.A(new_n448), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n664), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(new_n663), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(new_n523), .A3(new_n619), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n468), .A2(new_n584), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n534), .A3(new_n668), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n462), .A2(new_n465), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n701), .B1(new_n396), .B2(new_n421), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n710), .B(new_n711), .C1(new_n447), .C2(new_n458), .ZN(new_n712));
  INV_X1    g511(.A(new_n395), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n425), .B2(new_n426), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n457), .A3(new_n432), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n422), .B1(new_n715), .B2(KEYINPUT35), .ZN(new_n716));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n584), .C1(new_n712), .C2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n461), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n711), .A2(KEYINPUT107), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n459), .A2(new_n466), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n585), .B1(new_n721), .B2(new_n436), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n717), .B(new_n706), .C1(new_n722), .C2(KEYINPUT44), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n669), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n724), .ZN(G1328gat));
  OAI21_X1  g524(.A(G36gat), .B1(new_n723), .B2(new_n421), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n535), .A3(new_n457), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(G1329gat));
  OAI21_X1  g532(.A(G43gat), .B1(new_n723), .B2(new_n466), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n707), .A2(new_n525), .A3(new_n691), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G43gat), .B1(new_n723), .B2(new_n698), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n735), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g538(.A(G50gat), .B1(new_n723), .B2(new_n701), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n707), .A2(new_n527), .A3(new_n448), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g542(.A1(new_n523), .A2(new_n619), .A3(new_n585), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n663), .B(new_n744), .C1(new_n721), .C2(new_n436), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n668), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n665), .A2(KEYINPUT109), .A3(new_n667), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g551(.A1(new_n721), .A2(new_n436), .ZN(new_n753));
  INV_X1    g552(.A(new_n744), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n705), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n421), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  XNOR2_X1  g561(.A(new_n755), .B(KEYINPUT110), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n497), .B1(new_n763), .B2(new_n697), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n755), .B2(new_n692), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n745), .A2(KEYINPUT111), .A3(new_n691), .ZN(new_n767));
  AOI21_X1  g566(.A(G71gat), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n764), .A2(KEYINPUT50), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770));
  OAI21_X1  g569(.A(G71gat), .B1(new_n757), .B2(new_n698), .ZN(new_n771));
  INV_X1    g570(.A(new_n768), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n769), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n763), .A2(new_n448), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n523), .A2(new_n663), .A3(new_n618), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n717), .B(new_n777), .C1(new_n722), .C2(KEYINPUT44), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n669), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n705), .A2(new_n668), .A3(new_n565), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT112), .Z(new_n781));
  NOR2_X1   g580(.A1(new_n523), .A2(new_n618), .ZN(new_n782));
  AND4_X1   g581(.A1(KEYINPUT51), .A2(new_n753), .A3(new_n584), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n722), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n785), .ZN(G1336gat));
  NOR3_X1   g585(.A1(new_n778), .A2(new_n411), .A3(new_n421), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n753), .A2(new_n584), .A3(new_n782), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n722), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n663), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n457), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n787), .B1(new_n793), .B2(new_n411), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  AOI21_X1  g595(.A(G92gat), .B1(new_n792), .B2(new_n457), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n787), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(G1337gat));
  INV_X1    g598(.A(G99gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n778), .A2(new_n800), .A3(new_n698), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n792), .A2(new_n691), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n800), .ZN(G1338gat));
  OAI211_X1 g602(.A(new_n448), .B(new_n705), .C1(new_n783), .C2(new_n784), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n778), .B2(new_n701), .ZN(new_n806));
  INV_X1    g605(.A(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT113), .B1(new_n778), .B2(new_n701), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(G1339gat));
  INV_X1    g613(.A(new_n523), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n656), .B2(new_n649), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n648), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n816), .B(new_n647), .C1(new_n632), .C2(new_n640), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n653), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n820), .A3(KEYINPUT55), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n655), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT115), .B1(new_n824), .B2(new_n655), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n618), .B(new_n823), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n589), .B1(new_n601), .B2(new_n596), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n596), .A2(new_n597), .A3(new_n595), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n610), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n617), .B(new_n830), .C1(new_n661), .C2(new_n662), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n584), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n617), .A2(new_n830), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n822), .B2(new_n821), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n584), .B(new_n834), .C1(new_n825), .C2(new_n826), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n815), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n744), .A2(new_n705), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND4_X1   g639(.A1(KEYINPUT116), .A2(new_n840), .A3(new_n357), .A4(new_n750), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n749), .B1(new_n837), .B2(new_n839), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT116), .B1(new_n842), .B2(new_n357), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n421), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n619), .A2(G113gat), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT118), .Z(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n669), .A2(new_n457), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n840), .A2(new_n433), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n619), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(G1340gat));
  NOR2_X1   g652(.A1(new_n663), .A2(G120gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n845), .A2(new_n846), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G120gat), .B1(new_n851), .B2(new_n663), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n851), .A2(new_n858), .A3(new_n815), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n841), .A2(new_n843), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n523), .A3(new_n421), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(new_n858), .ZN(G1342gat));
  INV_X1    g661(.A(G134gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n584), .A2(new_n421), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT119), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n851), .B2(new_n585), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n860), .A2(new_n869), .A3(new_n863), .A4(new_n865), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n695), .A2(KEYINPUT122), .A3(new_n448), .A4(new_n696), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n697), .B2(new_n701), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n842), .A2(new_n421), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n288), .A3(new_n618), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n878), .B2(KEYINPUT121), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n840), .A2(new_n880), .A3(new_n448), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n850), .A2(new_n466), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n824), .A2(new_n655), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n821), .B(KEYINPUT120), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n618), .B(new_n885), .C1(new_n886), .C2(KEYINPUT55), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n584), .B1(new_n887), .B2(new_n831), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n815), .B1(new_n888), .B2(new_n836), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n701), .B1(new_n889), .B2(new_n839), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n881), .B(new_n883), .C1(new_n890), .C2(new_n880), .ZN(new_n891));
  OAI21_X1  g690(.A(G141gat), .B1(new_n891), .B2(new_n619), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n878), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n879), .B(new_n893), .ZN(G1344gat));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n290), .A3(new_n705), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n891), .B2(new_n663), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n290), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n880), .B(new_n701), .C1(new_n837), .C2(new_n839), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n705), .B(new_n883), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n895), .B1(new_n898), .B2(new_n902), .ZN(G1345gat));
  AND4_X1   g702(.A1(new_n750), .A2(new_n840), .A3(new_n875), .A4(new_n873), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n523), .A4(new_n421), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n876), .B2(new_n815), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n907), .A3(new_n294), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n523), .A2(G155gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n891), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n908), .B(KEYINPUT124), .C1(new_n891), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1346gat));
  OAI21_X1  g713(.A(G162gat), .B1(new_n891), .B2(new_n585), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n904), .A2(new_n295), .A3(new_n865), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1347gat));
  AOI21_X1  g716(.A(new_n421), .B1(new_n747), .B2(new_n748), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n618), .A2(new_n823), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n884), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n655), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n659), .A2(KEYINPUT101), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n833), .B1(new_n924), .B2(new_n660), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n585), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n523), .B1(new_n926), .B2(new_n835), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n433), .B(new_n918), .C1(new_n927), .C2(new_n838), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT125), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n840), .A2(new_n930), .A3(new_n433), .A4(new_n918), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n619), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n668), .B1(new_n837), .B2(new_n839), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(new_n457), .A3(new_n357), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n202), .A3(new_n618), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1348gat));
  NOR3_X1   g736(.A1(new_n932), .A2(new_n203), .A3(new_n663), .ZN(new_n938));
  AOI21_X1  g737(.A(G176gat), .B1(new_n935), .B2(new_n705), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(G1349gat));
  OAI21_X1  g739(.A(G183gat), .B1(new_n932), .B2(new_n815), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n523), .A3(new_n251), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n237), .A3(new_n584), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n584), .A3(new_n931), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(G190gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n946), .B2(G190gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n945), .B(KEYINPUT126), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1351gat));
  NOR3_X1   g753(.A1(new_n750), .A2(new_n697), .A3(new_n421), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n899), .B2(new_n900), .ZN(new_n956));
  OAI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n619), .ZN(new_n957));
  AND4_X1   g756(.A1(new_n457), .A2(new_n934), .A3(new_n448), .A4(new_n698), .ZN(new_n958));
  INV_X1    g757(.A(G197gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n959), .A3(new_n618), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n957), .A2(new_n960), .ZN(G1352gat));
  INV_X1    g760(.A(G204gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n958), .A2(new_n962), .A3(new_n705), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT62), .Z(new_n964));
  OAI211_X1 g763(.A(new_n705), .B(new_n955), .C1(new_n899), .C2(new_n900), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n313), .A3(new_n523), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n523), .B(new_n955), .C1(new_n899), .C2(new_n900), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n958), .A2(new_n314), .A3(new_n584), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g774(.A(KEYINPUT127), .B(new_n955), .C1(new_n899), .C2(new_n900), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n975), .A2(new_n584), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n977), .B2(new_n314), .ZN(G1355gat));
endmodule


