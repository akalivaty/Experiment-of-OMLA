//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NOR2_X1   g0048(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n214), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT68), .B1(new_n252), .B2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(new_n206), .A3(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n251), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n206), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n251), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n205), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G50), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n266), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n264), .B(new_n269), .C1(G50), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n271), .A2(new_n272), .B1(KEYINPUT71), .B2(KEYINPUT10), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n278), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n280), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(new_n285), .B2(G226), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n252), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT66), .B(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G222), .ZN(new_n292));
  XOR2_X1   g0092(.A(new_n292), .B(KEYINPUT67), .Z(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G223), .B1(G77), .B2(new_n296), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n286), .B1(new_n300), .B2(new_n280), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(new_n302), .A3(G200), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n275), .B(new_n303), .C1(new_n304), .C2(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n302), .B1(new_n301), .B2(G200), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n249), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n273), .A2(new_n274), .ZN(new_n308));
  INV_X1    g0108(.A(new_n301), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(G190), .ZN(new_n310));
  INV_X1    g0110(.A(new_n306), .ZN(new_n311));
  INV_X1    g0111(.A(new_n249), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .A4(new_n303), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n301), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT69), .B(G179), .Z(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n271), .C1(new_n301), .C2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n307), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n266), .A2(new_n218), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n267), .A2(G68), .A3(new_n268), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n256), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G50), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n262), .A2(new_n325), .B1(new_n206), .B2(G68), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n251), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT11), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n321), .B(new_n322), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n327), .A2(new_n328), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  INV_X1    g0133(.A(new_n280), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n291), .A2(G226), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G232), .A2(G1698), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n296), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n334), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n282), .B1(new_n285), .B2(G238), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT13), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n340), .B2(new_n341), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n333), .B(G169), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n344), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(new_n342), .A3(new_n341), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n333), .B1(new_n348), .B2(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n332), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(G200), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n331), .C1(new_n304), .C2(new_n348), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n288), .A2(new_n206), .A3(new_n289), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n289), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n218), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n224), .A2(new_n218), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n201), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n261), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n356), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n296), .B2(new_n206), .ZN(new_n367));
  INV_X1    g0167(.A(new_n360), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n365), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n371), .A3(new_n251), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n257), .B1(new_n205), .B2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n267), .B1(new_n257), .B2(new_n266), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(G226), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT66), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G1698), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n378), .B(new_n380), .C1(new_n294), .C2(new_n295), .ZN(new_n381));
  INV_X1    g0181(.A(G223), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n376), .B(new_n377), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n290), .A2(new_n291), .A3(G223), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n376), .A4(new_n377), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n334), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n281), .B1(new_n284), .B2(new_n225), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n314), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n280), .B1(new_n383), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n393), .B2(new_n387), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n316), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n375), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT18), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n372), .B(new_n374), .C1(new_n394), .C2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT73), .B(G190), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n398), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n372), .A2(new_n374), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n391), .A2(G200), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n403), .A4(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n372), .A2(new_n374), .B1(new_n394), .B2(new_n316), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n392), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n397), .A2(new_n405), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n355), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G244), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n281), .B1(new_n284), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n298), .A2(G238), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n416), .B1(new_n417), .B2(new_n290), .C1(new_n225), .C2(new_n381), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n418), .B2(new_n334), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n316), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT15), .B(G87), .Z(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n256), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n257), .A2(new_n262), .B1(new_n206), .B2(new_n323), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n251), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n267), .A2(G77), .A3(new_n268), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(G77), .C2(new_n270), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n419), .B2(G169), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n419), .B2(G190), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n399), .B2(new_n419), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n319), .A2(new_n413), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(G257), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G294), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n437), .C1(new_n381), .C2(new_n221), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT83), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n290), .A2(new_n291), .A3(G250), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT83), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(new_n436), .A4(new_n437), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n334), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n280), .A2(G274), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n277), .A2(G1), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  INV_X1    g0251(.A(new_n214), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n451), .A2(new_n445), .B1(new_n452), .B2(new_n279), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G264), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n399), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(G190), .B2(new_n455), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n417), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT25), .B1(new_n266), .B2(new_n417), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n252), .A2(G1), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n266), .A2(new_n251), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(G107), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n206), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n417), .A2(KEYINPUT23), .A3(G20), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n290), .A2(new_n206), .A3(G87), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT22), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n290), .A2(new_n474), .A3(new_n206), .A4(G87), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(new_n214), .B2(new_n250), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n296), .A2(G20), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n481), .B2(G87), .ZN(new_n482));
  INV_X1    g0282(.A(new_n475), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n470), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT81), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n476), .A2(new_n477), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(KEYINPUT24), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n464), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n457), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(KEYINPUT81), .A3(new_n479), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT24), .B1(new_n476), .B2(new_n477), .ZN(new_n491));
  AOI211_X1 g0291(.A(KEYINPUT81), .B(new_n471), .C1(new_n473), .C2(new_n475), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n251), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n493), .A2(new_n494), .A3(new_n463), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n493), .B2(new_n463), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n455), .A2(KEYINPUT84), .A3(G169), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n443), .A2(G179), .A3(new_n450), .A4(new_n454), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT84), .B1(new_n455), .B2(G169), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n489), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n414), .B1(new_n288), .B2(new_n289), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n291), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n291), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n280), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT76), .B1(new_n453), .B2(G257), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n448), .A2(G257), .A3(new_n280), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT76), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n450), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(G169), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n509), .A2(new_n507), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n511), .A3(new_n505), .A4(new_n504), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n334), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n453), .A2(KEYINPUT76), .A3(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n515), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n449), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n317), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n262), .A2(new_n323), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n417), .A2(KEYINPUT6), .A3(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n526), .B1(new_n532), .B2(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n417), .B1(new_n359), .B2(new_n360), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT74), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g0336(.A(KEYINPUT74), .B(new_n417), .C1(new_n359), .C2(new_n360), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n251), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n270), .A2(G97), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n462), .B2(G97), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n518), .A2(new_n525), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n538), .A2(KEYINPUT75), .A3(new_n540), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT75), .B1(new_n538), .B2(new_n540), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n521), .A2(new_n524), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n521), .A2(G190), .A3(new_n524), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n541), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n505), .B(new_n206), .C1(G33), .C2(new_n226), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n251), .C1(new_n206), .C2(G116), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT20), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n270), .A2(G116), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n462), .B2(G116), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n314), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT80), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n227), .B1(new_n288), .B2(new_n289), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n291), .ZN(new_n559));
  XOR2_X1   g0359(.A(KEYINPUT79), .B(G303), .Z(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n296), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n290), .A2(G264), .A3(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n557), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n291), .A2(new_n558), .B1(new_n560), .B2(new_n296), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(KEYINPUT80), .A3(new_n563), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n280), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n453), .A2(KEYINPUT78), .A3(G270), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n448), .A2(G270), .A3(new_n280), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n449), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n556), .B(KEYINPUT21), .C1(new_n568), .C2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT80), .B1(new_n566), .B2(new_n563), .ZN(new_n576));
  AND4_X1   g0376(.A1(KEYINPUT80), .A2(new_n559), .A3(new_n561), .A4(new_n563), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n334), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n553), .A2(new_n555), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n578), .A2(new_n573), .A3(new_n579), .A4(G179), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n573), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT21), .B1(new_n582), .B2(new_n556), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(G200), .ZN(new_n585));
  INV_X1    g0385(.A(new_n579), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n401), .C2(new_n582), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n256), .B2(new_n226), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n290), .A2(new_n206), .A3(G68), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n206), .B1(new_n338), .B2(new_n588), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n529), .A2(new_n220), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT77), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT77), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n589), .A2(new_n590), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n251), .B1(new_n266), .B2(new_n422), .ZN(new_n598));
  OAI211_X1 g0398(.A(G244), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n465), .B(new_n599), .C1(new_n381), .C2(new_n219), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n334), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n280), .B(G250), .C1(G1), .C2(new_n277), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n280), .A2(G274), .A3(new_n445), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n462), .A2(G87), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n601), .A2(G190), .A3(new_n605), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n598), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n594), .A2(new_n596), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n226), .B1(new_n253), .B2(new_n255), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n590), .B1(new_n612), .B2(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n251), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n422), .A2(new_n266), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n462), .A2(new_n421), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n601), .A2(new_n316), .A3(new_n605), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n606), .A2(new_n314), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n584), .A2(new_n587), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n503), .A2(new_n549), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n435), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n409), .A2(new_n410), .A3(new_n392), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n410), .B1(new_n409), .B2(new_n392), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n397), .A2(KEYINPUT87), .A3(new_n411), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n352), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n429), .B2(new_n354), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n405), .A2(new_n408), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n307), .A3(new_n313), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n318), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT88), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n639), .A3(new_n318), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n493), .A2(new_n463), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n500), .B2(new_n501), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n584), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n604), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n602), .A2(KEYINPUT85), .A3(new_n603), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n601), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n314), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n617), .A2(new_n649), .A3(new_n618), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n598), .A2(new_n608), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(G200), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n609), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n488), .B2(new_n457), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n644), .A2(new_n549), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n518), .A2(new_n525), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n542), .B2(new_n543), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n654), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT86), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n538), .A2(new_n540), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n658), .A2(new_n662), .A3(new_n620), .A4(new_n610), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n657), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n621), .A2(KEYINPUT86), .A3(KEYINPUT26), .A4(new_n541), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n656), .A2(new_n666), .A3(new_n650), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n641), .B1(new_n668), .B2(new_n435), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT89), .ZN(new_n672));
  INV_X1    g0472(.A(G213), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n502), .A2(new_n642), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n497), .A2(new_n502), .A3(new_n677), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n497), .A2(new_n677), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n682), .A2(new_n683), .B1(new_n503), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n584), .A2(new_n677), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n679), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT90), .B1(new_n584), .B2(new_n587), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n678), .A2(new_n586), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n584), .A2(KEYINPUT90), .A3(new_n587), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n584), .A2(new_n691), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n682), .A2(new_n683), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n503), .A2(new_n684), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n689), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(KEYINPUT92), .ZN(new_n704));
  INV_X1    g0504(.A(new_n209), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(G41), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n209), .A2(KEYINPUT92), .A3(new_n276), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n592), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n212), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT26), .B1(new_n659), .B2(new_n654), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n714));
  INV_X1    g0514(.A(new_n650), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n497), .A2(new_n502), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(new_n584), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n549), .A2(new_n655), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n713), .B(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n678), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n667), .A2(new_n678), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AND4_X1   g0525(.A1(new_n503), .A2(new_n622), .A3(new_n549), .A4(new_n678), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT93), .B1(new_n582), .B2(new_n349), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n578), .A2(new_n573), .A3(new_n728), .A4(G179), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n443), .A2(new_n454), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n545), .A2(new_n730), .A3(new_n606), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n316), .A2(new_n582), .A3(new_n545), .A4(new_n648), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n732), .A2(new_n733), .B1(new_n735), .B2(new_n455), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n737), .B2(new_n677), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n726), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n678), .B1(new_n734), .B2(new_n736), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT31), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n697), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n725), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n712), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(new_n708), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n265), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n205), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n698), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(G330), .B1(new_n694), .B2(new_n695), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT94), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n696), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n209), .A2(new_n290), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n209), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n705), .A2(new_n290), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n277), .B2(new_n213), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n244), .A2(new_n277), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n452), .B1(new_n206), .B2(G169), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT95), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT95), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n755), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n749), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT96), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n316), .A2(new_n206), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n399), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n774), .B2(new_n401), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n773), .A2(KEYINPUT96), .A3(new_n399), .A4(new_n402), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G322), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n774), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n773), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n401), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G311), .A2(new_n779), .B1(new_n781), .B2(G326), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n206), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n304), .A3(new_n399), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n290), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n206), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT98), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n790), .B1(G303), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n780), .A2(G190), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n783), .A2(new_n304), .A3(G200), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n798), .A2(new_n799), .B1(G283), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n778), .A2(new_n782), .A3(new_n797), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G50), .A2(new_n781), .B1(new_n779), .B2(G77), .ZN(new_n804));
  INV_X1    g0604(.A(new_n777), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n224), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n808), .A2(new_n218), .B1(new_n220), .B2(new_n795), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n801), .A2(G107), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n785), .A2(G159), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT32), .ZN(new_n812));
  INV_X1    g0612(.A(new_n789), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n811), .A2(KEYINPUT32), .B1(G97), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(new_n812), .A3(new_n814), .A4(new_n290), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n803), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n771), .B1(new_n817), .B2(new_n768), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n750), .A2(new_n752), .B1(new_n756), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  INV_X1    g0620(.A(new_n749), .ZN(new_n821));
  INV_X1    g0621(.A(new_n754), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n768), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n323), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n430), .A2(new_n677), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n427), .A2(new_n677), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n432), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n825), .B1(new_n827), .B2(new_n430), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G137), .A2(new_n781), .B1(new_n779), .B2(G159), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n260), .B2(new_n808), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G143), .B2(new_n777), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT34), .Z(new_n832));
  AOI21_X1  g0632(.A(new_n296), .B1(new_n785), .B2(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n224), .B2(new_n789), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n801), .A2(G68), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(G50), .C2(new_n796), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G283), .A2(new_n798), .B1(new_n781), .B2(G303), .ZN(new_n838));
  INV_X1    g0638(.A(G116), .ZN(new_n839));
  INV_X1    g0639(.A(new_n779), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  NAND2_X1  g0642(.A1(new_n796), .A2(G107), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n813), .A2(G97), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n801), .A2(G87), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n290), .B1(new_n785), .B2(G311), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G294), .B2(new_n777), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n832), .A2(new_n837), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n768), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n824), .B1(new_n828), .B2(new_n754), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n433), .A2(new_n677), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n667), .A2(KEYINPUT101), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT101), .B1(new_n667), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n828), .B1(new_n667), .B2(new_n678), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n742), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n749), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n858), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(KEYINPUT103), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n675), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n630), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n667), .A2(new_n852), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n667), .A2(KEYINPUT101), .A3(new_n852), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n825), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n332), .A2(new_n677), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n350), .A2(new_n351), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n355), .B2(KEYINPUT102), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n352), .A2(KEYINPUT102), .A3(new_n354), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT104), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n375), .A2(new_n392), .A3(new_n395), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n400), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n881), .A2(new_n403), .B1(new_n375), .B2(new_n864), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n675), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n375), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n396), .B(new_n885), .C1(new_n404), .C2(new_n400), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n412), .A2(new_n375), .A3(new_n884), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n889), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT104), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n865), .B1(new_n877), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n628), .A2(new_n633), .A3(new_n629), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n864), .A2(new_n375), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n901), .B(KEYINPUT87), .C1(new_n400), .C2(new_n404), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n882), .A2(new_n396), .B1(new_n904), .B2(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n400), .B2(new_n404), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NOR4_X1   g0707(.A1(new_n906), .A2(new_n879), .A3(KEYINPUT87), .A4(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n895), .B2(new_n896), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT105), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n908), .B(new_n905), .C1(new_n900), .C2(new_n902), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n912), .B(new_n896), .C1(new_n915), .C2(KEYINPUT38), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT39), .B1(new_n890), .B2(new_n891), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n914), .A2(new_n919), .A3(new_n631), .A4(new_n678), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n899), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n640), .A2(new_n638), .B1(new_n725), .B2(new_n434), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n921), .B(new_n922), .Z(new_n923));
  NAND3_X1  g0723(.A1(new_n873), .A2(new_n828), .A3(new_n875), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n739), .B2(new_n741), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT40), .B1(new_n925), .B2(new_n898), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n873), .A2(new_n828), .A3(new_n875), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n623), .A2(new_n677), .B1(new_n740), .B2(KEYINPUT31), .ZN(new_n928));
  INV_X1    g0728(.A(new_n741), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n910), .A2(new_n890), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n435), .B1(new_n741), .B2(new_n739), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n697), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n923), .A2(new_n937), .B1(new_n205), .B2(new_n746), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT106), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n923), .A2(new_n937), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(G116), .A3(new_n215), .A4(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n212), .A2(new_n323), .A3(new_n362), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n218), .A2(G50), .ZN(new_n949));
  OAI211_X1 g0749(.A(G1), .B(new_n265), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  OAI21_X1  g0751(.A(new_n549), .B1(new_n544), .B2(new_n678), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n659), .A2(new_n678), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n497), .A3(new_n502), .ZN(new_n955));
  INV_X1    g0755(.A(new_n541), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n677), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n685), .A2(new_n687), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n954), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n959), .B2(KEYINPUT42), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT42), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n961), .A3(new_n954), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n651), .A2(new_n677), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n715), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n654), .B2(new_n965), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n954), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n702), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n960), .A2(new_n962), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n968), .A2(new_n972), .ZN(new_n974));
  INV_X1    g0774(.A(new_n970), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n708), .B(KEYINPUT41), .ZN(new_n977));
  INV_X1    g0777(.A(new_n702), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n688), .A2(KEYINPUT44), .A3(new_n969), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT44), .B1(new_n688), .B2(new_n969), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n954), .B(new_n679), .C1(new_n685), .C2(new_n687), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT45), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n978), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n981), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n979), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n983), .B(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n989), .A3(new_n702), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n701), .A2(new_n686), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n992), .B2(new_n958), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n701), .A2(new_n686), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n685), .A2(new_n687), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(KEYINPUT107), .C2(new_n698), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n743), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n985), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n977), .B1(new_n998), .B2(new_n743), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n973), .B(new_n976), .C1(new_n999), .C2(new_n748), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n795), .A2(new_n839), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n789), .A2(new_n417), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n296), .B1(new_n784), .B2(new_n1004), .C1(new_n226), .C2(new_n800), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(new_n781), .C2(G311), .ZN(new_n1006));
  INV_X1    g0806(.A(G283), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n840), .C1(new_n787), .C2(new_n808), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1002), .B(new_n1008), .C1(new_n560), .C2(new_n777), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n777), .A2(G150), .B1(G68), .B2(new_n813), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT108), .Z(new_n1011));
  INV_X1    g0811(.A(G137), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n290), .B1(new_n784), .B2(new_n1012), .C1(new_n323), .C2(new_n800), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G50), .A2(new_n779), .B1(new_n781), .B2(G143), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n224), .B2(new_n795), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G159), .C2(new_n798), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1009), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n850), .B1(new_n1017), .B2(KEYINPUT47), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT47), .B2(new_n1017), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n770), .B1(new_n705), .B2(new_n421), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n760), .A2(new_n240), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n821), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n755), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1019), .B(new_n1022), .C1(new_n1023), .C2(new_n967), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1000), .A2(new_n1024), .ZN(G387));
  AND2_X1   g0825(.A1(new_n993), .A2(new_n996), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n685), .A2(new_n755), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n757), .A2(new_n709), .B1(G107), .B2(new_n209), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n236), .A2(G45), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n709), .B(new_n277), .C1(new_n218), .C2(new_n323), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1031));
  NOR3_X1   g0831(.A1(new_n1031), .A2(G50), .A3(new_n257), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(G50), .B2(new_n257), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n761), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1028), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n749), .B1(new_n1036), .B2(new_n770), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n795), .A2(new_n323), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n218), .A2(new_n840), .B1(new_n808), .B2(new_n257), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G97), .C2(new_n801), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n813), .A2(new_n421), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n290), .C1(new_n260), .C2(new_n784), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n781), .B2(G159), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(new_n325), .C2(new_n805), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n795), .A2(new_n787), .B1(new_n1007), .B2(new_n789), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n781), .A2(G322), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n798), .B1(new_n779), .B2(new_n560), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n805), .C2(new_n1004), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT49), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n290), .B1(new_n785), .B2(G326), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n839), .B2(new_n800), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1044), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1037), .B1(new_n1055), .B2(new_n768), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1026), .A2(new_n748), .B1(new_n1027), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n997), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n745), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1026), .A2(new_n743), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  NAND3_X1  g0861(.A1(new_n985), .A2(new_n990), .A3(new_n748), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n761), .A2(new_n247), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n769), .B1(new_n226), .B2(new_n209), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n798), .A2(new_n560), .B1(G116), .B2(new_n813), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n787), .B2(new_n840), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT111), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n290), .B1(new_n785), .B2(G322), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n810), .B(new_n1068), .C1(new_n1007), .C2(new_n795), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n777), .A2(G311), .B1(G317), .B2(new_n781), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  AOI22_X1  g0872(.A1(new_n777), .A2(G159), .B1(G150), .B2(new_n781), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n808), .A2(new_n325), .B1(new_n218), .B2(new_n795), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n840), .A2(new_n257), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n296), .B1(new_n785), .B2(G143), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n845), .B(new_n1078), .C1(new_n323), .C2(new_n789), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1070), .A2(new_n1072), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n749), .B1(new_n1063), .B2(new_n1064), .C1(new_n1081), .C2(new_n850), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT112), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1023), .B2(new_n954), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1062), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT113), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1062), .A2(KEYINPUT113), .A3(new_n1084), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n998), .A2(new_n745), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n985), .A2(new_n990), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n1058), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1089), .A2(new_n1093), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n631), .A2(new_n678), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n931), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n721), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n827), .A2(new_n430), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n825), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1095), .B(new_n1096), .C1(new_n1099), .C2(new_n876), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n914), .A2(new_n919), .ZN(new_n1101));
  OAI211_X1 g0901(.A(KEYINPUT114), .B(new_n1095), .C1(new_n870), .C2(new_n876), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n876), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n855), .B2(new_n825), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT114), .B1(new_n1105), .B2(new_n1095), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1100), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n742), .A2(new_n828), .A3(new_n1104), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1100), .B(new_n1108), .C1(new_n1103), .C2(new_n1106), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n828), .C1(new_n928), .C2(new_n929), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n876), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n855), .B2(new_n825), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1099), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n725), .A2(new_n434), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n742), .A2(new_n434), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n641), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1112), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1110), .A2(new_n1111), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n745), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1110), .A2(new_n748), .A3(new_n1111), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1101), .A2(new_n822), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n290), .B1(new_n785), .B2(G294), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n323), .B2(new_n789), .C1(new_n795), .C2(new_n220), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G97), .A2(new_n779), .B1(new_n781), .B2(G283), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n835), .C1(new_n417), .C2(new_n808), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G116), .C2(new_n777), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n795), .A2(new_n260), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1136));
  XNOR2_X1  g0936(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G137), .A2(new_n798), .B1(new_n779), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n296), .B1(new_n785), .B2(G125), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n325), .B2(new_n800), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G159), .B2(new_n813), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n781), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1140), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1137), .B(new_n1146), .C1(G132), .C2(new_n777), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n768), .B1(new_n1134), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n821), .B1(new_n257), .B2(new_n823), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT115), .Z(new_n1150));
  NAND3_X1  g0950(.A1(new_n1129), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1127), .A2(new_n1128), .A3(new_n1151), .ZN(G378));
  NOR2_X1   g0952(.A1(G33), .A2(G41), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G50), .B(new_n1153), .C1(new_n296), .C2(new_n276), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n800), .A2(new_n224), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT117), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n839), .A2(new_n1145), .B1(new_n840), .B2(new_n422), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G97), .C2(new_n798), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n276), .B(new_n296), .C1(new_n784), .C2(new_n1007), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1159), .B(new_n1038), .C1(G68), .C2(new_n813), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(new_n417), .C2(new_n805), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT58), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1154), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(G124), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(G124), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n785), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(new_n1153), .ZN(new_n1168));
  INV_X1    g0968(.A(G159), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n795), .A2(new_n1138), .B1(new_n260), .B2(new_n789), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G125), .A2(new_n781), .B1(new_n798), .B2(G132), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1012), .B2(new_n840), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G128), .C2(new_n777), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT59), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1168), .B1(new_n1169), .B2(new_n800), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1163), .B1(new_n1162), .B2(new_n1161), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n768), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n821), .B1(new_n325), .B2(new_n823), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n271), .A2(new_n884), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n319), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n307), .A2(new_n313), .A3(new_n318), .A4(new_n1180), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1178), .B(new_n1179), .C1(new_n1188), .C2(new_n754), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT119), .Z(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n934), .B2(G330), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n926), .A2(new_n933), .A3(new_n1187), .A4(new_n697), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n921), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n892), .A2(new_n897), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n932), .B1(new_n1194), .B2(new_n930), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n925), .A2(new_n1096), .A3(KEYINPUT40), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(G330), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1187), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1188), .A3(G330), .A4(new_n1196), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1198), .A2(new_n920), .A3(new_n899), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT120), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(KEYINPUT120), .B(new_n921), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1190), .B1(new_n1204), .B2(new_n748), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1121), .B(KEYINPUT121), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n1126), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1126), .A2(KEYINPUT122), .A3(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1204), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1193), .A2(new_n1200), .A3(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(KEYINPUT123), .B(new_n921), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1214), .A2(KEYINPUT57), .A3(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1126), .A2(KEYINPUT122), .A3(new_n1206), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT122), .B1(new_n1126), .B2(new_n1206), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n745), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1205), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT124), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(KEYINPUT124), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n1118), .A2(new_n748), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n290), .B1(new_n785), .B2(G303), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1041), .B(new_n1226), .C1(new_n795), .C2(new_n226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n798), .A2(G116), .B1(G77), .B2(new_n801), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n417), .B2(new_n840), .C1(new_n787), .C2(new_n1145), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(G283), .C2(new_n777), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G132), .A2(new_n781), .B1(new_n798), .B2(new_n1139), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n260), .B2(new_n840), .C1(new_n1169), .C2(new_n795), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n805), .A2(new_n1012), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n290), .B1(new_n784), .B2(new_n1144), .C1(new_n789), .C2(new_n325), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1232), .A2(new_n1156), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n768), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n821), .B1(new_n218), .B2(new_n823), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n1104), .C2(new_n754), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1225), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n977), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1116), .A2(new_n1121), .A3(new_n1117), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1123), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(G381));
  NOR4_X1   g1044(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1087), .A2(new_n1088), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1245), .A2(new_n1024), .A3(new_n1000), .A4(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(G375), .A2(G378), .A3(new_n1247), .ZN(G407));
  INV_X1    g1048(.A(G378), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n673), .A2(G343), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1205), .C1(new_n1212), .C2(new_n1220), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1241), .B(new_n1204), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1214), .A2(new_n748), .A3(new_n1215), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1189), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1249), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1253), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1242), .B1(new_n1125), .B2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1116), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n1117), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n745), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1240), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(G384), .A3(new_n1240), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1253), .A2(G2897), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT125), .Z(new_n1270));
  XNOR2_X1  g1070(.A(new_n1268), .B(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1252), .B1(new_n1259), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1268), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1259), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G390), .A2(new_n1024), .A3(new_n1000), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1246), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(new_n819), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1280), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1253), .B(new_n1268), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT63), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1273), .A2(new_n1277), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1285), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1275), .A2(new_n1289), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1272), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1282), .A2(new_n1283), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1280), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT127), .B1(new_n1298), .B2(new_n1281), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1295), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1287), .B1(new_n1293), .B2(new_n1300), .ZN(G405));
  OAI21_X1  g1101(.A(new_n1268), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1294), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1298), .A2(KEYINPUT127), .A3(new_n1281), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1274), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1221), .A2(G378), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1250), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1306), .B(new_n1308), .ZN(G402));
endmodule


