//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT2), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G155gat), .B(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n202), .A2(new_n207), .A3(new_n205), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT74), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT73), .B(G211gat), .Z(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G218gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n212), .B2(KEYINPUT74), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n214), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT72), .B(KEYINPUT22), .Z(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT73), .B(G211gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n212), .A2(KEYINPUT74), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n213), .A4(new_n218), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n220), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n211), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G228gat), .A2(G233gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n209), .A2(new_n229), .A3(new_n210), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n226), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(KEYINPUT82), .A3(new_n227), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G78gat), .B(G106gat), .Z(new_n241));
  XOR2_X1   g040(.A(KEYINPUT31), .B(G50gat), .Z(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT83), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n234), .A2(new_n237), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n231), .B1(new_n246), .B2(new_n230), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n240), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n244), .A2(KEYINPUT83), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G22gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n248), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G120gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n256), .A3(G113gat), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n253), .A2(G113gat), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT70), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(KEYINPUT70), .A3(new_n258), .ZN(new_n261));
  XOR2_X1   g060(.A(G127gat), .B(G134gat), .Z(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G120gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(KEYINPUT1), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n211), .A2(new_n264), .A3(KEYINPUT77), .A4(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT77), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n261), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(new_n259), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n209), .A2(new_n210), .A3(new_n266), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n252), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n209), .A2(new_n210), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n266), .B1(new_n269), .B2(new_n259), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n233), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n270), .A2(new_n271), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT4), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n273), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282));
  OR3_X1    g081(.A1(new_n281), .A2(KEYINPUT39), .A3(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT80), .ZN(new_n285));
  XNOR2_X1  g084(.A(G1gat), .B(G29gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n276), .A2(new_n274), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n267), .A2(new_n272), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n282), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(KEYINPUT39), .B(new_n293), .C1(new_n281), .C2(new_n282), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n283), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT40), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n291), .A2(new_n292), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT5), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n301));
  AOI211_X1 g100(.A(KEYINPUT78), .B(new_n301), .C1(new_n291), .C2(new_n292), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n267), .A2(new_n272), .A3(new_n252), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n279), .A2(KEYINPUT4), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(new_n282), .A3(new_n277), .ZN(new_n305));
  OAI22_X1  g104(.A1(new_n300), .A2(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n273), .A2(new_n280), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n307), .A2(new_n301), .A3(new_n282), .A4(new_n277), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n289), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n311));
  INV_X1    g110(.A(G226gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(KEYINPUT23), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n327));
  INV_X1    g126(.A(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n320), .A2(new_n325), .A3(new_n331), .A4(KEYINPUT25), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n331), .A2(KEYINPUT25), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n335), .A2(KEYINPUT66), .A3(new_n325), .A4(new_n320), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT23), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n331), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n334), .A2(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342));
  OR3_X1    g141(.A1(new_n341), .A2(new_n321), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n341), .B2(new_n321), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n324), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(KEYINPUT26), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT27), .B(G183gat), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT67), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n349), .A2(new_n351), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n315), .B1(new_n356), .B2(KEYINPUT29), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n237), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT76), .B(new_n315), .C1(new_n356), .C2(KEYINPUT29), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n334), .A2(new_n336), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n339), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n354), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n314), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT75), .B1(new_n356), .B2(new_n315), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n369), .A3(new_n314), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n357), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n237), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n311), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n377), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n367), .A2(new_n372), .A3(KEYINPUT30), .A4(new_n376), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n295), .B2(new_n296), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n295), .A2(new_n382), .A3(new_n296), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n310), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n386));
  INV_X1    g185(.A(new_n373), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT37), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n377), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(KEYINPUT87), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n389), .A2(KEYINPUT87), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n387), .A2(new_n391), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n386), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n388), .B1(new_n371), .B2(new_n360), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n359), .A2(new_n237), .A3(new_n361), .A4(new_n366), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n394), .A2(new_n398), .B1(new_n376), .B2(new_n387), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n306), .A2(new_n308), .ZN(new_n400));
  INV_X1    g199(.A(new_n289), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n306), .A2(new_n308), .A3(new_n289), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n309), .A2(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n251), .B(new_n385), .C1(new_n393), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT34), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n364), .A2(new_n276), .A3(new_n354), .ZN(new_n410));
  INV_X1    g209(.A(new_n276), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n340), .B2(new_n355), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n409), .A3(new_n414), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(KEYINPUT71), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n414), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420));
  XOR2_X1   g219(.A(G15gat), .B(G43gat), .Z(new_n421));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n419), .B(KEYINPUT32), .C1(new_n420), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(KEYINPUT32), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n420), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n423), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT71), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n413), .A2(new_n429), .A3(new_n409), .A4(new_n414), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n417), .A2(new_n425), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n425), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n416), .A2(KEYINPUT71), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n414), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT34), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n404), .A2(new_n403), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n309), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n406), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n251), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n441), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n438), .A2(new_n251), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT35), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n431), .A2(new_n437), .A3(new_n251), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n404), .A2(new_n403), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n406), .B1(new_n458), .B2(new_n309), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n459), .A3(new_n448), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT88), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n456), .B1(new_n405), .B2(new_n406), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n448), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n408), .A2(new_n451), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G113gat), .B(G141gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(G197gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT11), .B(G169gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT12), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474));
  INV_X1    g273(.A(G15gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(G22gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(G15gat), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(G15gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n475), .A2(G22gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT93), .ZN(new_n482));
  INV_X1    g281(.A(G1gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT16), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(G1gat), .B1(new_n479), .B2(new_n482), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n472), .B(new_n473), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n482), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT93), .B1(new_n480), .B2(new_n481), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n473), .ZN(new_n492));
  NAND2_X1  g291(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n496));
  INV_X1    g295(.A(G43gat), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT15), .B1(new_n497), .B2(G50gat), .ZN(new_n498));
  INV_X1    g297(.A(G50gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(G43gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G29gat), .A2(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n501), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT92), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n505), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT14), .B1(new_n502), .B2(new_n503), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n512), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n497), .A2(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n499), .A2(G43gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT15), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT92), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n517), .A2(new_n518), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT90), .B(KEYINPUT15), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n520), .B1(new_n500), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n499), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n496), .B(new_n513), .C1(new_n523), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n526), .B1(new_n497), .B2(G50gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n497), .A2(G50gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n524), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n501), .A2(new_n512), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n535), .A2(new_n522), .A3(new_n536), .A4(new_n517), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n496), .B1(new_n537), .B2(new_n513), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n495), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n513), .B1(new_n523), .B2(new_n529), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n487), .A2(new_n541), .A3(new_n494), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(KEYINPUT18), .A3(new_n540), .A4(new_n542), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n540), .B(KEYINPUT13), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n541), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n495), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(new_n542), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AND4_X1   g351(.A1(new_n471), .A2(new_n545), .A3(new_n546), .A4(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n543), .B2(new_n544), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n471), .B1(new_n554), .B2(new_n546), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(G85gat), .A3(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT8), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n560), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT100), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G99gat), .ZN(new_n572));
  INV_X1    g371(.A(G106gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n566), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n568), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n568), .A2(new_n577), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n531), .A2(new_n538), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n579), .A2(new_n578), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n541), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n580), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT98), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n580), .B(new_n592), .C1(new_n586), .C2(new_n587), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT102), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n594), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n602));
  OAI211_X1 g401(.A(KEYINPUT96), .B(G57gat), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(G71gat), .ZN(new_n605));
  INV_X1    g404(.A(G78gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT9), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G57gat), .ZN(new_n610));
  OR2_X1    g409(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n600), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n613));
  INV_X1    g412(.A(G64gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(G57gat), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n603), .B(new_n609), .C1(new_n612), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G57gat), .B(G64gat), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n604), .B(new_n607), .C1(new_n617), .C2(new_n608), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n495), .B1(new_n620), .B2(new_n619), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT97), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n599), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n619), .B1(new_n579), .B2(new_n578), .ZN(new_n639));
  AND2_X1   g438(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n642), .A2(new_n558), .B1(KEYINPUT8), .B2(new_n566), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n643), .A2(new_n571), .A3(new_n576), .A4(new_n565), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n568), .A2(new_n577), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n644), .A2(new_n616), .A3(new_n618), .A4(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n639), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n619), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n638), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n637), .B1(new_n639), .B2(new_n646), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n651), .B2(new_n652), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n466), .A2(new_n556), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n447), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n448), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(KEYINPUT42), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(KEYINPUT42), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n671), .B(new_n672), .C1(new_n473), .C2(new_n668), .ZN(G1325gat));
  INV_X1    g472(.A(new_n441), .ZN(new_n674));
  OAI21_X1  g473(.A(G15gat), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n663), .A2(new_n475), .A3(new_n438), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n450), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n451), .A2(new_n408), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n454), .A2(new_n465), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n556), .A2(new_n634), .A3(new_n660), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n684), .A2(new_n599), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n502), .A3(new_n664), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(new_n598), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n594), .B(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n466), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n463), .B1(new_n462), .B2(new_n448), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n463), .A2(new_n457), .A3(new_n459), .A4(new_n448), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n381), .B1(new_n446), .B2(new_n406), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n455), .B1(new_n695), .B2(new_n452), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n454), .A2(new_n465), .A3(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n697), .A2(new_n699), .B1(new_n408), .B2(new_n451), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n691), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n685), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n447), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n705), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n686), .A2(new_n503), .A3(new_n381), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT46), .Z(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n704), .B2(new_n448), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1329gat));
  NAND2_X1  g509(.A1(new_n441), .A2(G43gat), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n686), .A2(new_n438), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n704), .A2(new_n711), .B1(G43gat), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n702), .B1(new_n715), .B2(new_n682), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n684), .B2(new_n599), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n450), .B(new_n685), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n703), .A2(KEYINPUT105), .A3(new_n450), .A4(new_n685), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(G50gat), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n251), .A2(G50gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n686), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT48), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n719), .A2(G50gat), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT48), .B1(new_n729), .B2(new_n725), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n731), .A3(KEYINPUT106), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n499), .B1(new_n719), .B2(new_n720), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n726), .B1(new_n734), .B2(new_n722), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n735), .B2(new_n730), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(G1331gat));
  NAND2_X1  g536(.A1(new_n715), .A2(new_n682), .ZN(new_n738));
  INV_X1    g537(.A(new_n556), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n599), .A2(new_n739), .A3(new_n635), .A4(new_n661), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n664), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(G57gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  INV_X1    g543(.A(new_n741), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n448), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n741), .A2(new_n438), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n741), .A2(KEYINPUT108), .A3(new_n438), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n605), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n741), .A2(G71gat), .A3(new_n441), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT50), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n450), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n739), .A2(new_n634), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n703), .A2(new_n660), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n664), .ZN(new_n766));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n690), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n738), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n738), .B(new_n770), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n664), .A2(new_n558), .A3(new_n660), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n766), .A2(new_n558), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  NAND4_X1  g575(.A1(new_n703), .A2(new_n381), .A3(new_n660), .A4(new_n764), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n641), .B2(new_n640), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n448), .A2(G92gat), .A3(new_n661), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n772), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1337gat));
  AOI21_X1  g582(.A(new_n572), .B1(new_n765), .B2(new_n441), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n438), .A2(new_n572), .A3(new_n660), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n774), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT111), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n784), .B2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1338gat));
  AOI21_X1  g590(.A(new_n573), .B1(new_n765), .B2(new_n450), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n251), .A2(G106gat), .A3(new_n661), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n772), .A2(new_n773), .A3(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT53), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1339gat));
  NAND3_X1  g596(.A1(new_n636), .A2(new_n556), .A3(new_n661), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n540), .B1(new_n539), .B2(new_n542), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n550), .A2(new_n542), .A3(new_n548), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n470), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n540), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n805), .A2(new_n530), .B1(new_n487), .B2(new_n494), .ZN(new_n806));
  INV_X1    g605(.A(new_n542), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n550), .A2(new_n542), .A3(new_n548), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(KEYINPUT112), .A3(new_n470), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n554), .A2(new_n471), .A3(new_n546), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n648), .A2(new_n650), .A3(new_n638), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n816), .A2(new_n651), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n648), .A2(new_n650), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n817), .A3(new_n637), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n656), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n815), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n637), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n648), .A2(new_n650), .A3(new_n638), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n655), .B1(new_n651), .B2(new_n817), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n822), .A2(new_n658), .A3(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n690), .A2(new_n814), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT112), .B1(new_n810), .B2(new_n470), .ZN(new_n830));
  INV_X1    g629(.A(new_n470), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n802), .B(new_n831), .C1(new_n808), .C2(new_n809), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n813), .B(new_n660), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n556), .B2(new_n828), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n599), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n825), .A2(new_n826), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n657), .B1(new_n837), .B2(new_n815), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n827), .C1(new_n555), .C2(new_n553), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n829), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n798), .B1(new_n841), .B2(new_n634), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n452), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n664), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n448), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT115), .Z(new_n848));
  NOR2_X1   g647(.A1(new_n556), .A2(G113gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n664), .A3(new_n448), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n556), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1340gat));
  AND3_X1   g652(.A1(new_n660), .A2(new_n254), .A3(new_n256), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G120gat), .B1(new_n851), .B2(new_n661), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n851), .B2(new_n635), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n635), .A2(G127gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n847), .B2(new_n859), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n381), .A2(new_n690), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  INV_X1    g663(.A(new_n862), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n844), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n441), .A2(new_n447), .A3(new_n381), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n842), .A2(new_n869), .A3(new_n450), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(G141gat), .A3(new_n556), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n833), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n812), .A2(KEYINPUT118), .A3(new_n813), .A4(new_n660), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n839), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n690), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n690), .A2(new_n828), .A3(new_n814), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n634), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n798), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT57), .B(new_n450), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n829), .B1(new_n690), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n798), .B1(new_n884), .B2(new_n634), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n450), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  XNOR2_X1  g687(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n888), .B(new_n890), .C1(new_n842), .C2(new_n450), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n834), .A2(new_n835), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n690), .A3(new_n840), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n634), .B1(new_n893), .B2(new_n878), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n450), .B1(new_n894), .B2(new_n880), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT117), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n887), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n869), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n556), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(G141gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n872), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT120), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n895), .A2(new_n889), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n888), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n895), .A2(KEYINPUT117), .A3(new_n889), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n903), .B(new_n869), .C1(new_n907), .C2(new_n887), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n739), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n871), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n901), .B1(new_n910), .B2(new_n911), .ZN(G1344gat));
  NAND2_X1  g711(.A1(new_n885), .A2(new_n450), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n842), .A2(new_n450), .A3(new_n890), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n661), .A3(new_n898), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G148gat), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT59), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n660), .A3(new_n908), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  INV_X1    g724(.A(G148gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(KEYINPUT59), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n924), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n870), .A2(G148gat), .A3(new_n661), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1345gat));
  OAI21_X1  g731(.A(new_n203), .B1(new_n870), .B2(new_n635), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n902), .A2(new_n908), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n634), .A2(G155gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n934), .B2(new_n690), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n674), .A2(new_n664), .A3(new_n204), .A4(new_n862), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n895), .B2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n664), .A2(new_n448), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n843), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n328), .A3(new_n556), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n842), .A2(new_n447), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n381), .A3(new_n452), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n739), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n948), .B2(new_n328), .ZN(G1348gat));
  OAI21_X1  g748(.A(G176gat), .B1(new_n943), .B2(new_n661), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n660), .A2(new_n329), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n946), .B2(new_n951), .ZN(G1349gat));
  OAI21_X1  g751(.A(G183gat), .B1(new_n943), .B2(new_n635), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n634), .A2(new_n347), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n955), .B(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n843), .A2(new_n599), .A3(new_n942), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G190gat), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT61), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n947), .A2(new_n348), .A3(new_n599), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT125), .Z(G1351gat));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n450), .A3(new_n381), .A4(new_n674), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(G197gat), .B1(new_n966), .B2(new_n739), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n942), .A2(new_n674), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT126), .Z(new_n969));
  NOR2_X1   g768(.A1(new_n969), .A2(new_n918), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n739), .A2(G197gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT127), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n965), .A2(G204gat), .A3(new_n661), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n969), .A2(new_n918), .A3(new_n661), .ZN(new_n976));
  INV_X1    g775(.A(G204gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G1353gat));
  INV_X1    g777(.A(G211gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n968), .A2(new_n635), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n917), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT63), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n223), .A3(new_n634), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1354gat));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n222), .A3(new_n599), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n918), .A3(new_n690), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n222), .ZN(G1355gat));
endmodule


