//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n206), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n204), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n213), .B(new_n216), .C1(new_n218), .C2(new_n220), .ZN(G361));
  XNOR2_X1  g0021(.A(G238), .B(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT2), .B(G226), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n226), .B(new_n229), .Z(G358));
  XNOR2_X1  g0030(.A(G50), .B(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XOR2_X1   g0032(.A(G58), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G351));
  INV_X1    g0038(.A(KEYINPUT14), .ZN(new_n239));
  INV_X1    g0039(.A(KEYINPUT13), .ZN(new_n240));
  INV_X1    g0040(.A(KEYINPUT67), .ZN(new_n241));
  NOR2_X1   g0041(.A1(G226), .A2(G1698), .ZN(new_n242));
  AOI21_X1  g0042(.A(new_n242), .B1(new_n223), .B2(G1698), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n243), .A2(new_n248), .B1(G33), .B2(G97), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(G1), .B(G13), .C1(new_n245), .C2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n241), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n223), .A2(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n253), .B1(G226), .B2(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(KEYINPUT67), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n250), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n251), .A2(G274), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G238), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n240), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  AOI211_X1 g0070(.A(KEYINPUT13), .B(new_n268), .C1(new_n252), .C2(new_n260), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n239), .B(G169), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT67), .B1(new_n258), .B2(new_n259), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n241), .B(new_n251), .C1(new_n256), .C2(new_n257), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n261), .A2(new_n240), .A3(new_n269), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G179), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n277), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n239), .B1(new_n280), .B2(G169), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT68), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n270), .A2(new_n271), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT14), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n278), .A4(new_n272), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(new_n204), .A3(G1), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT12), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n291), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n204), .A2(G33), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n217), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(KEYINPUT11), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n290), .A2(new_n300), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n203), .A2(G20), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(G68), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT11), .B1(new_n298), .B2(new_n300), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n288), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n283), .A2(G190), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n280), .A2(G200), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(new_n307), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT16), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n246), .A2(new_n204), .A3(new_n247), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n246), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n247), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n291), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G58), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n291), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G58), .A2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n294), .A2(G159), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n314), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n300), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n317), .A2(new_n318), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n325), .B1(new_n330), .B2(G68), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  OAI211_X1 g0132(.A(KEYINPUT69), .B(new_n314), .C1(new_n319), .C2(new_n325), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n203), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n302), .B1(new_n290), .B2(new_n335), .ZN(new_n337));
  XOR2_X1   g0137(.A(new_n337), .B(KEYINPUT70), .Z(new_n338));
  NAND2_X1  g0138(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n264), .B1(new_n266), .B2(new_n223), .ZN(new_n340));
  INV_X1    g0140(.A(G226), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G223), .B2(G1698), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n254), .A2(new_n255), .ZN(new_n344));
  INV_X1    g0144(.A(G87), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n343), .A2(new_n344), .B1(new_n245), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n346), .B2(new_n259), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT66), .B(G179), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n284), .B2(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT18), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n339), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G200), .B2(new_n347), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n334), .A2(new_n358), .A3(new_n338), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT71), .A2(KEYINPUT17), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT71), .B(KEYINPUT17), .Z(new_n362));
  NAND4_X1  g0162(.A1(new_n334), .A2(new_n358), .A3(new_n338), .A4(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n353), .A2(new_n355), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n264), .B1(new_n266), .B2(new_n341), .ZN(new_n365));
  INV_X1    g0165(.A(G1698), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n344), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G223), .B1(G77), .B2(new_n344), .ZN(new_n368));
  INV_X1    g0168(.A(G222), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n248), .A2(new_n366), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n365), .B1(new_n371), .B2(new_n259), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n302), .A2(G50), .A3(new_n303), .ZN(new_n375));
  INV_X1    g0175(.A(new_n290), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(G50), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n294), .A2(G150), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n335), .B2(new_n297), .ZN(new_n379));
  INV_X1    g0179(.A(G50), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n204), .B1(new_n322), .B2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n377), .B1(new_n300), .B2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n383), .A2(KEYINPUT9), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n372), .A2(G190), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(KEYINPUT9), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n374), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT10), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n373), .B2(new_n284), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n349), .B2(new_n373), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n335), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n297), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n300), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n296), .B1(new_n203), .B2(G20), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n302), .A2(new_n397), .B1(new_n296), .B2(new_n290), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G244), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n264), .B1(new_n266), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n367), .A2(G238), .B1(G107), .B2(new_n344), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n223), .B2(new_n370), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(new_n259), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n399), .B1(new_n404), .B2(G190), .ZN(new_n405));
  INV_X1    g0205(.A(G200), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n404), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n348), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n399), .C1(G169), .C2(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR4_X1   g0210(.A1(new_n313), .A2(new_n364), .A3(new_n391), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT19), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n204), .B1(new_n257), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G97), .A2(G107), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n345), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n204), .B(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n417));
  INV_X1    g0217(.A(G97), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n412), .B1(new_n297), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n300), .B1(new_n290), .B2(new_n394), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n203), .A2(G33), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT74), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(G87), .A3(new_n302), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n203), .A2(G45), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n251), .A2(G274), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n251), .A2(G250), .A3(new_n425), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(G244), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n430));
  OAI211_X1 g0230(.A(G238), .B(new_n366), .C1(new_n254), .C2(new_n255), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G116), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n429), .B1(new_n259), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n421), .B(new_n424), .C1(new_n434), .C2(new_n406), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n259), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n427), .A2(new_n428), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(G190), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n434), .A2(KEYINPUT78), .A3(G190), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n434), .A2(new_n348), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n423), .A2(new_n302), .ZN(new_n444));
  INV_X1    g0244(.A(new_n394), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n421), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(new_n437), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n284), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT79), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n450), .ZN(new_n452));
  INV_X1    g0252(.A(new_n435), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n441), .A2(new_n440), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  AND4_X1   g0259(.A1(G274), .A2(new_n459), .A3(new_n251), .A4(new_n426), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n259), .B1(new_n426), .B2(new_n459), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(G270), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n248), .A2(G1698), .ZN(new_n463));
  INV_X1    g0263(.A(G264), .ZN(new_n464));
  INV_X1    g0264(.A(G303), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n248), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n370), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(G1698), .B1(new_n246), .B2(new_n247), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(KEYINPUT80), .A3(G257), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n462), .B1(new_n472), .B2(new_n251), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G200), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n475), .B(new_n204), .C1(G33), .C2(new_n418), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n300), .C1(new_n204), .C2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n290), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n423), .A2(new_n302), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n479), .B(new_n481), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n474), .B(new_n484), .C1(new_n356), .C2(new_n473), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  INV_X1    g0286(.A(new_n460), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n461), .A2(G270), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n469), .A2(new_n471), .ZN(new_n490));
  INV_X1    g0290(.A(new_n466), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(new_n259), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n477), .B(KEYINPUT20), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n481), .B1(new_n482), .B2(new_n480), .ZN(new_n495));
  OAI21_X1  g0295(.A(G169), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n486), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n483), .A3(G179), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n473), .A2(new_n483), .A3(KEYINPUT21), .A4(G169), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n485), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n458), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(G244), .B(new_n366), .C1(new_n254), .C2(new_n255), .ZN(new_n502));
  NOR2_X1   g0302(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n248), .A2(G244), .A3(new_n366), .A4(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G250), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n475), .A4(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(new_n259), .B1(G257), .B2(new_n461), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n284), .B1(new_n509), .B2(new_n487), .ZN(new_n510));
  INV_X1    g0310(.A(new_n504), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n475), .B(new_n507), .C1(new_n502), .C2(new_n503), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n259), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n461), .A2(G257), .ZN(new_n514));
  AND4_X1   g0314(.A1(new_n349), .A2(new_n513), .A3(new_n487), .A4(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n330), .A2(KEYINPUT73), .A3(G107), .ZN(new_n517));
  INV_X1    g0317(.A(G107), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(KEYINPUT72), .A3(KEYINPUT6), .A4(G97), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g0320(.A1(KEYINPUT6), .A2(G97), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(G107), .ZN(new_n522));
  AND2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n414), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n519), .B(new_n522), .C1(new_n524), .C2(KEYINPUT6), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT73), .B1(new_n330), .B2(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n300), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n376), .A2(G97), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n444), .B2(G97), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(KEYINPUT77), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT77), .B1(new_n529), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n516), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n531), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT75), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(KEYINPUT75), .A3(new_n531), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n509), .A2(new_n487), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n406), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n509), .A2(new_n356), .A3(new_n487), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n468), .A2(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n248), .B(new_n546), .C1(G250), .C2(G1698), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n259), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n459), .A2(new_n426), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n251), .A2(G274), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n461), .A2(G264), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n553), .A3(new_n356), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n550), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(G200), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT23), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(new_n204), .A3(G107), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT23), .B1(new_n518), .B2(G20), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(G20), .B2(new_n432), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n248), .A2(new_n204), .A3(G87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n248), .A2(new_n563), .A3(new_n204), .A4(G87), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT24), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(KEYINPUT24), .B(new_n560), .C1(new_n562), .C2(new_n564), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n300), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT25), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n376), .B2(G107), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n518), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n444), .A2(G107), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n556), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n284), .B1(new_n550), .B2(new_n553), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n550), .A2(new_n553), .ZN(new_n577));
  INV_X1    g0377(.A(G179), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n555), .A2(KEYINPUT81), .A3(G179), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(new_n569), .B2(new_n573), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT82), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n580), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n569), .A2(new_n573), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n556), .A2(new_n569), .A3(new_n573), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n411), .A2(new_n501), .A3(new_n545), .A4(new_n589), .ZN(G372));
  NAND2_X1  g0390(.A1(new_n361), .A2(new_n363), .ZN(new_n591));
  INV_X1    g0391(.A(new_n312), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n592), .A2(new_n409), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n309), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n353), .A2(new_n355), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n388), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(new_n390), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n348), .A2(new_n434), .B1(new_n446), .B2(new_n421), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT83), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT83), .B1(new_n427), .B2(new_n428), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n436), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n284), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n421), .A2(new_n424), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(G200), .B2(new_n602), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n454), .B1(new_n599), .B2(new_n603), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n587), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n499), .A2(new_n497), .A3(new_n498), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n585), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n605), .B1(new_n545), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n510), .A2(new_n515), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT77), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n536), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n532), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(KEYINPUT26), .A3(new_n457), .A4(new_n451), .ZN(new_n617));
  INV_X1    g0417(.A(new_n539), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT75), .B1(new_n529), .B2(new_n531), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n516), .B(new_n608), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n612), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n411), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n598), .A2(new_n625), .ZN(G369));
  NAND3_X1  g0426(.A1(new_n499), .A2(new_n497), .A3(new_n498), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n629), .A2(G213), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G343), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT84), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n484), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n500), .B2(new_n634), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G330), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n633), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n584), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT86), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT86), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n588), .A2(new_n582), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n585), .A2(new_n633), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n610), .A2(new_n641), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n585), .B2(new_n641), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g0452(.A(new_n652), .B(KEYINPUT87), .Z(G399));
  INV_X1    g0453(.A(new_n214), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n220), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n415), .A2(G116), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G1), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n610), .A2(new_n585), .ZN(new_n661));
  INV_X1    g0461(.A(new_n609), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n544), .A3(new_n535), .A4(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n616), .A2(new_n621), .A3(new_n457), .A4(new_n451), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n663), .A2(new_n604), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(KEYINPUT29), .A3(new_n633), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n641), .B1(new_n612), .B2(new_n623), .ZN(new_n668));
  XOR2_X1   g0468(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n667), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n513), .A2(new_n514), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n673), .A2(new_n577), .A3(new_n448), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(KEYINPUT30), .A3(G179), .A4(new_n493), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n555), .A2(new_n349), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n473), .A3(new_n540), .A4(new_n602), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n555), .A2(new_n509), .A3(new_n434), .ZN(new_n679));
  OAI211_X1 g0479(.A(G179), .B(new_n462), .C1(new_n472), .C2(new_n251), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n675), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n641), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT88), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n682), .A2(new_n688), .A3(KEYINPUT31), .A4(new_n641), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n684), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n501), .A2(new_n589), .A3(new_n545), .A4(new_n633), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n672), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n671), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n660), .B1(new_n695), .B2(G1), .ZN(G364));
  AND2_X1   g0496(.A1(new_n638), .A2(new_n639), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n289), .A2(G20), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n203), .B1(new_n698), .B2(G45), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n655), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n697), .B(new_n702), .C1(G330), .C2(new_n636), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT90), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n214), .A2(G355), .A3(new_n248), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G116), .B2(new_n214), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n248), .B(new_n654), .C1(new_n262), .C2(new_n220), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n234), .A2(G45), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n217), .B1(G20), .B2(new_n284), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n701), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n348), .A2(new_n204), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G190), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G311), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n204), .A2(G179), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(G190), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n356), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n578), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  AOI22_X1  g0527(.A1(G303), .A2(new_n724), .B1(new_n727), .B2(G294), .ZN(new_n728));
  INV_X1    g0528(.A(G283), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n722), .A2(new_n356), .A3(G200), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(new_n344), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n722), .A2(new_n718), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT91), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT91), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n721), .B(new_n731), .C1(G329), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n717), .A2(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G190), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n717), .A2(new_n725), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n739), .A2(new_n740), .B1(new_n742), .B2(G322), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n738), .A2(new_n356), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G326), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n737), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n736), .A2(G159), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT32), .ZN(new_n749));
  INV_X1    g0549(.A(new_n745), .ZN(new_n750));
  INV_X1    g0550(.A(new_n739), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n380), .A2(new_n750), .B1(new_n751), .B2(new_n291), .ZN(new_n752));
  INV_X1    g0552(.A(new_n730), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G107), .A2(new_n753), .B1(new_n727), .B2(G97), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n754), .B(new_n248), .C1(new_n345), .C2(new_n723), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n320), .A2(new_n741), .B1(new_n719), .B2(new_n296), .ZN(new_n756));
  OR3_X1    g0556(.A1(new_n752), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n747), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n716), .B1(new_n758), .B2(new_n713), .ZN(new_n759));
  INV_X1    g0559(.A(new_n712), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n636), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n703), .A2(KEYINPUT90), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n704), .A2(new_n761), .A3(new_n762), .ZN(G396));
  NOR2_X1   g0563(.A1(new_n409), .A2(new_n641), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n641), .A2(new_n399), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n407), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n764), .B1(new_n766), .B2(new_n409), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n668), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n692), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n692), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n702), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n772), .B2(KEYINPUT95), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(KEYINPUT95), .B2(new_n772), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT96), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n713), .A2(new_n710), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n719), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G143), .A2(new_n742), .B1(new_n778), .B2(G159), .ZN(new_n779));
  INV_X1    g0579(.A(G150), .ZN(new_n780));
  INV_X1    g0580(.A(G137), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n779), .B1(new_n751), .B2(new_n780), .C1(new_n781), .C2(new_n750), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT34), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n753), .A2(G68), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n380), .B2(new_n723), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT93), .Z(new_n788));
  INV_X1    g0588(.A(new_n727), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n248), .B1(new_n789), .B2(new_n320), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n736), .B2(G132), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n784), .A2(new_n785), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n735), .A2(new_n720), .B1(new_n793), .B2(new_n741), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G116), .B2(new_n778), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n745), .A2(G303), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n739), .A2(G283), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n753), .A2(G87), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n518), .B2(new_n723), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n248), .B(new_n799), .C1(G97), .C2(new_n727), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n792), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n713), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n701), .B1(G77), .B2(new_n777), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT94), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT94), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(new_n711), .C2(new_n767), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n774), .A2(new_n775), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n775), .B1(new_n774), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G384));
  NOR2_X1   g0611(.A1(new_n698), .A2(new_n203), .ZN(new_n812));
  INV_X1    g0612(.A(new_n631), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n596), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n332), .A2(new_n326), .ZN(new_n815));
  INV_X1    g0615(.A(new_n337), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n813), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n364), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n339), .A2(new_n631), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT37), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n352), .A2(new_n820), .A3(new_n821), .A4(new_n359), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n815), .A2(new_n816), .B1(new_n351), .B2(new_n631), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n823), .A2(new_n359), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n824), .B2(new_n821), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n819), .A2(KEYINPUT38), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT38), .B1(new_n819), .B2(new_n825), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n617), .A2(new_n622), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n587), .B(new_n608), .C1(new_n627), .C2(new_n581), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n535), .A2(new_n544), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n604), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n633), .B(new_n767), .C1(new_n829), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n764), .B(KEYINPUT98), .Z(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n633), .A2(new_n307), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n309), .A2(new_n312), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n308), .B(new_n641), .C1(new_n288), .C2(new_n592), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n833), .A2(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT99), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n828), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n833), .A2(new_n835), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(new_n839), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n843), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n814), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT100), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n814), .C1(new_n842), .C2(new_n845), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n309), .A2(new_n641), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n819), .A2(KEYINPUT38), .A3(new_n825), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT102), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n813), .B1(new_n334), .B2(new_n338), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n352), .A4(new_n359), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n352), .A2(new_n820), .A3(new_n359), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n856), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n364), .A2(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n855), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(KEYINPUT102), .B(KEYINPUT38), .C1(new_n863), .C2(new_n864), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT103), .B(new_n854), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n822), .A2(KEYINPUT101), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n872), .A2(new_n860), .B1(new_n364), .B2(new_n857), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT102), .B1(new_n873), .B2(KEYINPUT38), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n865), .A2(new_n855), .A3(new_n866), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT103), .B1(new_n876), .B2(new_n854), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n850), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n847), .A2(new_n849), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n411), .B(new_n667), .C1(new_n668), .C2(new_n670), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n598), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT104), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n879), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n826), .B1(new_n874), .B2(new_n875), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n687), .A2(new_n683), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n768), .B1(new_n885), .B2(new_n691), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n844), .A2(new_n886), .A3(KEYINPUT40), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n844), .A2(new_n886), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n826), .A2(new_n827), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n885), .A2(new_n691), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n411), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n895), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(G330), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n812), .B1(new_n883), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n883), .B2(new_n898), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n901), .A2(G116), .A3(new_n218), .A4(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n321), .A2(new_n219), .A3(new_n296), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n291), .A2(G50), .ZN(new_n907));
  OAI211_X1 g0707(.A(G1), .B(new_n289), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n905), .A3(new_n908), .ZN(G367));
  NAND2_X1  g0709(.A1(new_n641), .A2(new_n606), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n608), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n604), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n645), .A2(new_n646), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n697), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n538), .A2(new_n539), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n545), .B1(new_n917), .B2(new_n633), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n516), .A3(new_n641), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT106), .ZN(new_n923));
  INV_X1    g0723(.A(new_n920), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n647), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n921), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n913), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n928), .ZN(new_n930));
  INV_X1    g0730(.A(new_n913), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(new_n926), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n924), .A2(new_n649), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT42), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n616), .B1(new_n920), .B2(new_n581), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n641), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n929), .A2(new_n932), .A3(new_n938), .A4(new_n937), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n655), .B(KEYINPUT41), .Z(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT45), .B1(new_n651), .B2(new_n920), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n650), .A2(new_n944), .A3(new_n924), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n650), .A2(KEYINPUT44), .A3(new_n924), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT44), .B1(new_n650), .B2(new_n924), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n647), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n914), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n649), .B1(new_n952), .B2(new_n648), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(new_n640), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n695), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n946), .A2(new_n949), .A3(new_n647), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n951), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n942), .B1(new_n958), .B2(new_n695), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n940), .B(new_n941), .C1(new_n959), .C2(new_n700), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n654), .A2(new_n248), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n229), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n715), .B1(new_n654), .B2(new_n445), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n702), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT108), .B(G317), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n736), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n730), .A2(new_n418), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n248), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(new_n720), .C2(new_n750), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G294), .B2(new_n739), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n778), .A2(G283), .B1(G107), .B2(new_n727), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n723), .A2(new_n480), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n741), .A2(new_n465), .B1(KEYINPUT46), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(KEYINPUT46), .B2(new_n974), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n727), .A2(G68), .ZN(new_n978));
  INV_X1    g0778(.A(G143), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n780), .B2(new_n741), .C1(new_n750), .C2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT109), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n248), .B1(new_n730), .B2(new_n296), .C1(new_n320), .C2(new_n723), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n735), .A2(new_n781), .B1(new_n380), .B2(new_n719), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G159), .C2(new_n739), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n981), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n982), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT47), .Z(new_n989));
  OAI221_X1 g0789(.A(new_n964), .B1(new_n760), .B2(new_n912), .C1(new_n989), .C2(new_n803), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n960), .A2(new_n990), .ZN(G387));
  OR3_X1    g0791(.A1(new_n226), .A2(new_n262), .A3(new_n248), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT50), .B1(new_n335), .B2(G50), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n262), .C1(new_n291), .C2(new_n296), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n335), .A2(KEYINPUT50), .A3(G50), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n344), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n657), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n654), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n714), .B1(new_n214), .B2(new_n518), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n701), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n380), .A2(new_n741), .B1(new_n719), .B2(new_n291), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n736), .B2(G150), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n745), .A2(G159), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n739), .A2(new_n392), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n789), .A2(new_n394), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n723), .A2(new_n296), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1005), .A2(new_n967), .A3(new_n1006), .A4(new_n344), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n789), .A2(new_n729), .B1(new_n723), .B2(new_n793), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G303), .A2(new_n778), .B1(new_n742), .B2(new_n965), .ZN(new_n1010));
  INV_X1    g0810(.A(G322), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n751), .B2(new_n720), .C1(new_n1011), .C2(new_n750), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT48), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n736), .A2(G326), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n248), .B1(new_n753), .B2(G116), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1008), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1000), .B1(new_n1022), .B2(new_n713), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n914), .A2(new_n712), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n954), .A2(new_n700), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n955), .A2(new_n655), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n954), .A2(new_n695), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(G393));
  AND2_X1   g0828(.A1(new_n951), .A2(new_n957), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n924), .A2(new_n712), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n961), .A2(new_n237), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n714), .B1(new_n214), .B2(new_n418), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n745), .A2(G317), .B1(new_n742), .B2(G311), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT52), .Z(new_n1034));
  AOI22_X1  g0834(.A1(G283), .A2(new_n724), .B1(new_n727), .B2(G116), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n344), .C1(new_n518), .C2(new_n730), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n735), .A2(new_n1011), .B1(new_n793), .B2(new_n719), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G303), .C2(new_n739), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n745), .A2(G150), .B1(new_n742), .B2(G159), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT51), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n724), .A2(G68), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n727), .A2(G77), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n798), .A2(new_n1041), .A3(new_n1042), .A4(new_n248), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n735), .A2(new_n979), .B1(new_n335), .B2(new_n719), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G50), .C2(new_n739), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1034), .A2(new_n1038), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n701), .B1(new_n1031), .B2(new_n1032), .C1(new_n1046), .C2(new_n803), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT111), .Z(new_n1048));
  AOI22_X1  g0848(.A1(new_n1029), .A2(new_n700), .B1(new_n1030), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1029), .A2(new_n956), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n958), .A2(new_n655), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G390));
  NAND3_X1  g0852(.A1(new_n844), .A2(new_n886), .A3(G330), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n672), .B(new_n768), .C1(new_n690), .C2(new_n691), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n844), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n666), .A2(new_n633), .A3(new_n767), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n835), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n838), .A2(new_n839), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n894), .A2(G330), .A3(new_n767), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1054), .A2(new_n844), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1055), .A2(new_n843), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n411), .A2(G330), .A3(new_n894), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n880), .A2(new_n598), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1056), .A2(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n884), .A2(new_n850), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n854), .B1(new_n867), .B2(new_n868), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT103), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n870), .A3(new_n869), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT112), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n840), .B2(new_n850), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n850), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n834), .B1(new_n668), .B2(new_n767), .ZN(new_n1076));
  OAI211_X1 g0876(.A(KEYINPUT112), .B(new_n1075), .C1(new_n1076), .C2(new_n1058), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1068), .B(new_n1061), .C1(new_n1072), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n891), .A2(new_n852), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n853), .B1(new_n874), .B2(new_n875), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n1082), .B2(KEYINPUT103), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1083), .A2(new_n1071), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1053), .B1(new_n1084), .B2(new_n1068), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1066), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n884), .A2(new_n1067), .A3(new_n850), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n871), .A2(new_n877), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1079), .B(new_n1065), .C1(new_n1090), .C2(new_n1053), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n655), .A3(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n700), .B(new_n1079), .C1(new_n1090), .C2(new_n1053), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n701), .B1(new_n392), .B2(new_n777), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n745), .A2(G128), .B1(new_n742), .B2(G132), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT113), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  AOI22_X1  g0897(.A1(new_n736), .A2(G125), .B1(new_n778), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n723), .A2(new_n780), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n344), .B1(new_n727), .B2(G159), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n380), .B2(new_n730), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n739), .B2(G137), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n736), .A2(G294), .B1(G116), .B2(new_n742), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n248), .B1(new_n724), .B2(G87), .ZN(new_n1106));
  AND4_X1   g0906(.A1(new_n786), .A2(new_n1105), .A3(new_n1042), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n751), .A2(new_n518), .B1(new_n719), .B2(new_n418), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT114), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(new_n729), .C2(new_n750), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1108), .A2(KEYINPUT114), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1104), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1094), .B1(new_n1112), .B2(new_n713), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1072), .B2(new_n711), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1093), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1092), .A2(new_n1115), .ZN(G378));
  INV_X1    g0916(.A(new_n1064), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1091), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1091), .A2(KEYINPUT117), .A3(new_n1117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n878), .A2(new_n849), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n383), .A2(new_n813), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n391), .B(new_n1124), .Z(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n888), .A2(new_n1127), .A3(G330), .A4(new_n892), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n892), .B(G330), .C1(new_n884), .C2(new_n887), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1125), .B(new_n1126), .Z(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1123), .A2(new_n847), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1128), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n879), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT57), .B1(new_n1122), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT57), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1091), .A2(KEYINPUT117), .A3(new_n1117), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT117), .B1(new_n1091), .B2(new_n1117), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n655), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1130), .A2(new_n710), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n701), .B1(G50), .B2(new_n777), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n735), .A2(new_n729), .B1(new_n394), .B2(new_n719), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n248), .A2(G41), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n978), .A2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1006), .B(new_n1148), .C1(G58), .C2(new_n753), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n418), .B2(new_n751), .C1(new_n480), .C2(new_n750), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1146), .B(new_n1150), .C1(G107), .C2(new_n742), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT115), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT58), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n380), .B1(G33), .B2(G41), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n724), .A2(new_n1097), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n789), .A2(new_n780), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(G128), .C2(new_n742), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G125), .A2(new_n745), .B1(new_n739), .B2(G132), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n781), .C2(new_n719), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n736), .A2(G124), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(G41), .C1(new_n753), .C2(G159), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1153), .B1(new_n1147), .B2(new_n1154), .C1(new_n1160), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT116), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n803), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1145), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1135), .A2(new_n700), .B1(new_n1144), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1143), .A2(new_n1170), .ZN(G375));
  NAND2_X1  g0971(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n942), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1066), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1062), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1058), .A2(new_n710), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n701), .B1(G68), .B2(new_n777), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n344), .B1(new_n730), .B2(new_n296), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1178), .B(new_n1005), .C1(G97), .C2(new_n724), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n751), .B2(new_n480), .C1(new_n793), .C2(new_n750), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n736), .A2(G303), .B1(G283), .B2(new_n742), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n518), .B2(new_n719), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n736), .A2(G128), .B1(G137), .B2(new_n742), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n780), .B2(new_n719), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n739), .A2(new_n1097), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n745), .A2(G132), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n344), .B1(new_n753), .B2(G58), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G159), .A2(new_n724), .B1(new_n727), .B2(G50), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1180), .A2(new_n1182), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1177), .B1(new_n1190), .B2(new_n713), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1175), .A2(new_n700), .B1(new_n1176), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1174), .A2(new_n1192), .ZN(G381));
  INV_X1    g0993(.A(G375), .ZN(new_n1194));
  INV_X1    g0994(.A(G378), .ZN(new_n1195));
  OR3_X1    g0995(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1196), .A2(G387), .A3(G384), .A4(G381), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(G407));
  INV_X1    g0998(.A(G343), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(G213), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1194), .A2(new_n1195), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(G407), .A2(new_n1202), .A3(G213), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT118), .ZN(G409));
  INV_X1    g1004(.A(KEYINPUT124), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n655), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT60), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1055), .A2(new_n843), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1064), .A2(new_n1209), .A3(new_n1210), .A4(KEYINPUT60), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT120), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1062), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n1064), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1208), .A2(KEYINPUT121), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT121), .B1(new_n1208), .B2(new_n1215), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1192), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(G384), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n810), .B(new_n1192), .C1(new_n1217), .C2(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1201), .A2(G2897), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G378), .B(new_n1170), .C1(new_n1136), .C2(new_n1142), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n879), .A2(new_n1133), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n879), .A2(new_n1133), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1173), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1169), .A2(new_n1144), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1135), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n699), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1195), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT119), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n942), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1170), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT119), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1195), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1225), .A2(new_n1234), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1224), .B1(new_n1240), .B2(new_n1200), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1205), .B1(new_n1241), .B2(KEYINPUT61), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1238), .B1(new_n1237), .B2(new_n1195), .ZN(new_n1244));
  AOI211_X1 g1044(.A(KEYINPUT119), .B(G378), .C1(new_n1236), .C2(new_n1170), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1201), .B1(new_n1246), .B2(new_n1225), .ZN(new_n1247));
  OAI211_X1 g1047(.A(KEYINPUT124), .B(new_n1243), .C1(new_n1247), .C2(new_n1224), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1240), .A2(new_n1200), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1252), .A3(new_n1249), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1242), .A2(new_n1248), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT122), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n960), .A2(G390), .A3(new_n990), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n960), .B2(new_n990), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  XOR2_X1   g1058(.A(G393), .B(G396), .Z(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1255), .B(new_n1261), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1254), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1260), .A2(new_n1243), .A3(new_n1262), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT123), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1265), .B(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1241), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1250), .A2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1264), .A2(new_n1272), .ZN(G405));
  NAND3_X1  g1073(.A1(new_n1260), .A2(KEYINPUT125), .A3(new_n1262), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1274), .B(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G375), .A2(new_n1195), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1225), .A3(new_n1249), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1263), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1225), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1220), .A3(new_n1219), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1276), .A2(new_n1278), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1274), .B(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(G402));
endmodule


