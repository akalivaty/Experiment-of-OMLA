//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127, new_n1128, new_n1129;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT68), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n462), .B2(new_n464), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OAI211_X1 g052(.A(KEYINPUT69), .B(G125), .C1(new_n472), .C2(new_n473), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n471), .B1(new_n479), .B2(G2105), .ZN(G160));
  NAND2_X1  g055(.A1(new_n462), .A2(new_n464), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n465), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n467), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT70), .Z(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n472), .B2(new_n473), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n466), .B2(new_n489), .ZN(new_n494));
  OAI211_X1 g069(.A(KEYINPUT71), .B(new_n490), .C1(new_n472), .C2(new_n473), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n481), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G2105), .B1(G102), .B2(new_n469), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n504), .A2(new_n506), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n504), .A3(new_n506), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n503), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n512), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT72), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT7), .Z(new_n519));
  NAND2_X1  g094(.A1(new_n507), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT73), .B(G89), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n520), .B(new_n521), .C1(new_n510), .C2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(G168));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT5), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G543), .ZN(new_n528));
  AND4_X1   g103(.A1(new_n526), .A2(new_n528), .A3(new_n504), .A4(new_n506), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G90), .B1(new_n507), .B2(G52), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT74), .Z(new_n531));
  AOI22_X1  g106(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n503), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n528), .ZN(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n529), .A2(G81), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n507), .A2(G43), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n507), .A2(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n537), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n529), .B2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n529), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n507), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT78), .ZN(G288));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n503), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n529), .A2(G86), .B1(new_n507), .B2(G48), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n537), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n577), .A2(KEYINPUT79), .A3(G651), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n507), .A2(G47), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n510), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n503), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n582), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n529), .A2(G92), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT10), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n503), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n507), .A2(G54), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n586), .B1(G868), .B2(new_n593), .ZN(G284));
  OAI21_X1  g169(.A(new_n586), .B1(G868), .B2(new_n593), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n591), .A2(new_n592), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n596), .ZN(new_n604));
  INV_X1    g179(.A(new_n549), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n596), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g183(.A1(new_n472), .A2(new_n473), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n468), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT13), .B(G2100), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n482), .A2(G123), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n467), .A2(G135), .ZN(new_n616));
  OR2_X1    g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n620), .ZN(G156));
  XOR2_X1   g196(.A(KEYINPUT15), .B(G2435), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT83), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2443), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n635), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT85), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT86), .Z(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT87), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(KEYINPUT17), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n644), .A2(new_n648), .A3(new_n642), .ZN(new_n650));
  INV_X1    g225(.A(new_n645), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n651), .A2(new_n643), .A3(new_n642), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(KEYINPUT20), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(KEYINPUT20), .C2(new_n663), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  NOR2_X1   g250(.A1(G16), .A2(G19), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n549), .B2(G16), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(G1341), .Z(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n679), .A2(G26), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n482), .A2(G128), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n467), .A2(G140), .ZN(new_n682));
  NOR2_X1   g257(.A1(G104), .A2(G2105), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n680), .B1(new_n685), .B2(G29), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n680), .B(new_n686), .S(KEYINPUT28), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2067), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G4), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n593), .B2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(G1348), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n678), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(new_n619), .ZN(new_n698));
  INV_X1    g273(.A(G28), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(KEYINPUT30), .ZN(new_n700));
  AOI21_X1  g275(.A(G29), .B1(new_n699), .B2(KEYINPUT30), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n698), .A2(G29), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI22_X1  g277(.A1(G129), .A2(new_n482), .B1(new_n467), .B2(G141), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n469), .A2(G105), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n702), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n710), .B2(new_n711), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT31), .B(G11), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT99), .B(G1956), .Z(new_n715));
  INV_X1    g290(.A(G299), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT23), .B1(new_n716), .B2(new_n689), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n689), .A2(G20), .ZN(new_n718));
  MUX2_X1   g293(.A(KEYINPUT23), .B(new_n717), .S(new_n718), .Z(new_n719));
  OAI211_X1 g294(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n689), .A2(G5), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G171), .B2(new_n689), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1961), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT96), .B1(G29), .B2(G33), .ZN(new_n724));
  OR3_X1    g299(.A1(KEYINPUT96), .A2(G29), .A3(G33), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n467), .A2(G139), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n469), .A2(G103), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  INV_X1    g304(.A(new_n609), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n727), .B(new_n729), .C1(new_n465), .C2(new_n731), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n724), .B(new_n725), .C1(new_n732), .C2(new_n679), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT98), .B(G2072), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n720), .A2(new_n723), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G35), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G162), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n689), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n689), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(new_n679), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n679), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2084), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n715), .B2(new_n719), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n736), .A2(new_n741), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n696), .A2(new_n697), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n679), .A2(G27), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n679), .ZN(new_n755));
  INV_X1    g330(.A(G2078), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n679), .A2(G25), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n467), .A2(G131), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT88), .ZN(new_n761));
  OR2_X1    g336(.A1(G95), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n482), .A2(G119), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n679), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT35), .B(G1991), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n767), .B(new_n768), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n689), .A2(G24), .ZN(new_n770));
  INV_X1    g345(.A(G290), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n689), .ZN(new_n772));
  INV_X1    g347(.A(G1986), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n689), .A2(G22), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n689), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT91), .B(G1971), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n689), .A2(G23), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n569), .A2(KEYINPUT90), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n566), .A2(new_n781), .A3(new_n567), .A4(new_n568), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n779), .B1(new_n783), .B2(new_n689), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT89), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n778), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n769), .B(new_n774), .C1(new_n791), .C2(KEYINPUT34), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT92), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT93), .Z(new_n795));
  AOI21_X1  g370(.A(new_n758), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n793), .A2(new_n795), .A3(new_n758), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n753), .B(new_n757), .C1(new_n796), .C2(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  AOI22_X1  g374(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n503), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT100), .Z(new_n802));
  AOI22_X1  g377(.A1(new_n529), .A2(G93), .B1(new_n507), .B2(G55), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT101), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT102), .B(G860), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT37), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n549), .A2(new_n805), .ZN(new_n809));
  INV_X1    g384(.A(new_n805), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(new_n545), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n602), .A2(new_n600), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n812), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n808), .B1(new_n816), .B2(new_n806), .ZN(G145));
  INV_X1    g392(.A(KEYINPUT103), .ZN(new_n818));
  XNOR2_X1  g393(.A(G160), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G162), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(new_n698), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n707), .B(new_n685), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G164), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT104), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n732), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n732), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n825), .B2(new_n823), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n821), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n482), .A2(G130), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n467), .A2(G142), .ZN(new_n831));
  NOR2_X1   g406(.A1(G106), .A2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT105), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n612), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n766), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n829), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g416(.A(new_n812), .B(new_n603), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n593), .A2(G299), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n602), .A2(new_n716), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT106), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT107), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n843), .A2(new_n844), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT41), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n845), .A2(KEYINPUT107), .A3(new_n849), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(new_n842), .ZN(new_n857));
  XNOR2_X1  g432(.A(G303), .B(G290), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n783), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G305), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT42), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n848), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n848), .B2(new_n857), .ZN(new_n863));
  OAI21_X1  g438(.A(G868), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(G868), .B2(new_n810), .ZN(G295));
  OAI21_X1  g440(.A(new_n864), .B1(G868), .B2(new_n810), .ZN(G331));
  XNOR2_X1  g441(.A(G301), .B(G286), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n812), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n809), .A2(new_n811), .A3(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n855), .A3(new_n854), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n845), .A3(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n860), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT108), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n872), .A2(new_n860), .A3(new_n876), .A4(new_n873), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n879));
  INV_X1    g454(.A(new_n860), .ZN(new_n880));
  INV_X1    g455(.A(new_n873), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n869), .A2(new_n870), .B1(new_n850), .B2(new_n853), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n860), .B1(new_n872), .B2(new_n873), .ZN(new_n885));
  AOI211_X1 g460(.A(G37), .B(new_n885), .C1(new_n875), .C2(new_n877), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n878), .A2(KEYINPUT43), .A3(new_n883), .ZN(new_n890));
  INV_X1    g465(.A(new_n885), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT43), .B1(new_n878), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT44), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(G397));
  XNOR2_X1  g469(.A(KEYINPUT110), .B(G40), .ZN(new_n895));
  AOI211_X1 g470(.A(new_n471), .B(new_n895), .C1(new_n479), .C2(G2105), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT50), .ZN(new_n897));
  INV_X1    g472(.A(G1384), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n501), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT112), .ZN(new_n901));
  AND4_X1   g476(.A1(new_n901), .A2(new_n501), .A3(new_n897), .A4(new_n898), .ZN(new_n902));
  AOI21_X1  g477(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n903), .B2(new_n897), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n896), .B(new_n900), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G1961), .ZN(new_n906));
  XOR2_X1   g481(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n907));
  OR2_X1    g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(KEYINPUT45), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n908), .A2(new_n756), .A3(new_n896), .A4(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT53), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n905), .A2(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n908), .A2(KEYINPUT53), .A3(G40), .A4(new_n756), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(G160), .A3(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G171), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n501), .A2(new_n898), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n903), .A2(new_n907), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n920), .A2(new_n756), .A3(new_n896), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT122), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n911), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n912), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n917), .B(KEYINPUT54), .C1(new_n926), .C2(G171), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT123), .ZN(new_n928));
  INV_X1    g503(.A(G8), .ZN(new_n929));
  NAND2_X1  g504(.A1(G303), .A2(G8), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n479), .A2(G2105), .ZN(new_n932));
  INV_X1    g507(.A(new_n895), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n470), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n899), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n935), .B(new_n740), .C1(new_n904), .C2(new_n902), .ZN(new_n936));
  INV_X1    g511(.A(G1971), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n909), .A2(new_n896), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n903), .A2(new_n907), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g515(.A(new_n929), .B(new_n931), .C1(new_n936), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n934), .A2(new_n918), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n929), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n507), .A2(G48), .ZN(new_n944));
  INV_X1    g519(.A(G86), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n510), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n572), .A2(new_n503), .ZN(new_n947));
  OAI21_X1  g522(.A(G1981), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1981), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n573), .A2(new_n574), .A3(new_n578), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT49), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT115), .Z(new_n952));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n948), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n948), .B2(new_n950), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR4_X1   g534(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT114), .A4(KEYINPUT49), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n943), .B(new_n952), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n896), .A2(new_n903), .ZN(new_n962));
  INV_X1    g537(.A(G1976), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n783), .A2(G1976), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n962), .A2(G8), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(G8), .B(new_n965), .C1(new_n934), .C2(new_n918), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT52), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n961), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n941), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n931), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n896), .B(KEYINPUT116), .C1(new_n897), .C2(new_n903), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n899), .B2(new_n934), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n903), .A2(new_n897), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n972), .A2(new_n974), .A3(new_n740), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n940), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n971), .B1(new_n977), .B2(G8), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n928), .B1(new_n970), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n968), .A2(new_n966), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n962), .A2(G8), .ZN(new_n982));
  INV_X1    g557(.A(new_n956), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n948), .A2(new_n950), .A3(new_n954), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n958), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT114), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n957), .A2(new_n953), .A3(new_n958), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n981), .B1(new_n988), .B2(new_n952), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n936), .A2(new_n940), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(G8), .A3(new_n971), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n992), .A2(KEYINPUT123), .A3(new_n978), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n927), .B1(new_n980), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2084), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n935), .B(new_n995), .C1(new_n904), .C2(new_n902), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n920), .A2(new_n896), .A3(new_n921), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n744), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G8), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G168), .A2(new_n929), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT51), .B(G8), .C1(new_n999), .C2(G286), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n999), .A2(new_n1002), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1009));
  NAND3_X1  g584(.A1(new_n912), .A2(new_n915), .A3(G301), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G301), .B1(new_n925), .B2(new_n912), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT124), .B1(new_n994), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT117), .B(G1956), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n716), .A2(KEYINPUT57), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n559), .A2(KEYINPUT118), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n559), .A2(KEYINPUT118), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n563), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n938), .A2(new_n939), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT56), .B(G2072), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1018), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n903), .A2(new_n901), .A3(new_n897), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1348), .B1(new_n1035), .B2(new_n935), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n934), .A2(new_n918), .A3(G2067), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n905), .A2(new_n692), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1037), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(KEYINPUT120), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1031), .A2(new_n1038), .A3(new_n593), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1027), .B1(new_n1018), .B2(new_n1030), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT120), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1032), .B(new_n1037), .C1(new_n905), .C2(new_n692), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT60), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(new_n1048), .A3(new_n1041), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n593), .A3(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT60), .B(new_n602), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(KEYINPUT61), .A3(new_n1031), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1031), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1043), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1996), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1028), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT58), .B(G1341), .Z(new_n1059));
  NAND2_X1  g634(.A1(new_n962), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n605), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT59), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1042), .B(new_n1044), .C1(new_n1056), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n926), .A2(G171), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1010), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1065), .A2(new_n1009), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n970), .A2(new_n979), .A3(new_n928), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT123), .B1(new_n992), .B2(new_n978), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1066), .A2(new_n1067), .A3(new_n1070), .A4(new_n927), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1015), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1006), .A2(new_n1073), .A3(new_n1007), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(new_n1012), .C1(new_n980), .C2(new_n993), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1070), .A2(KEYINPUT125), .A3(new_n1012), .A4(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n969), .A2(new_n991), .ZN(new_n1081));
  INV_X1    g656(.A(G288), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n961), .A2(new_n963), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n982), .B1(new_n1083), .B2(new_n950), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n999), .A2(G8), .A3(G168), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n971), .B1(new_n990), .B2(G8), .ZN(new_n1087));
  OR4_X1    g662(.A1(new_n1085), .A2(new_n992), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n970), .A2(new_n979), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1089), .B2(new_n1086), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1081), .B(new_n1084), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1072), .A2(new_n1080), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n908), .A2(new_n934), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT111), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n685), .B(G2067), .Z(new_n1095));
  XNOR2_X1  g670(.A(new_n707), .B(new_n1057), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n765), .A2(new_n768), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n765), .A2(new_n768), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n771), .A2(new_n773), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G290), .A2(G1986), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1094), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1092), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1094), .A2(new_n1104), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT48), .Z(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(G2067), .B2(new_n685), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1094), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1094), .A2(new_n1057), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT46), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1113), .B(new_n1115), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1095), .A2(new_n708), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1094), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT127), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1116), .B(new_n1119), .C1(new_n1114), .C2(KEYINPUT46), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1120), .A2(KEYINPUT47), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(KEYINPUT47), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1109), .B(new_n1112), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1106), .A2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g699(.A(G319), .ZN(new_n1126));
  NOR2_X1   g700(.A1(G229), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g701(.A(new_n656), .B1(new_n638), .B2(new_n640), .ZN(new_n1128));
  AOI21_X1  g702(.A(new_n1128), .B1(new_n838), .B2(new_n839), .ZN(new_n1129));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n1127), .A3(new_n1129), .ZN(G225));
  INV_X1    g704(.A(G225), .ZN(G308));
endmodule


