//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT9), .B(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(new_n191), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  INV_X1    g009(.A(G953), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(G227), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n195), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G104), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT76), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n201), .B1(new_n206), .B2(new_n200), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n204), .A2(G104), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(KEYINPUT76), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n200), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT77), .B1(new_n211), .B2(KEYINPUT3), .ZN(new_n212));
  AOI21_X1  g026(.A(G107), .B1(new_n203), .B2(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(new_n199), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n208), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G101), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n221), .A2(KEYINPUT64), .A3(G146), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT64), .B1(new_n221), .B2(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n214), .B1(new_n213), .B2(new_n199), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT76), .B(G104), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n232), .C2(G107), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n207), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT78), .B(G101), .Z(new_n235));
  AOI21_X1  g049(.A(new_n217), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n216), .A2(G101), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT79), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT79), .B1(new_n236), .B2(new_n237), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n218), .B(new_n230), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n245), .A3(new_n249), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n200), .A2(G104), .ZN(new_n253));
  OAI21_X1  g067(.A(G101), .B1(new_n213), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT80), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(G101), .C1(new_n213), .C2(new_n253), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n234), .A2(new_n235), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n220), .A3(new_n222), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n260), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n220), .B2(new_n222), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n258), .B(new_n259), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  INV_X1    g081(.A(new_n235), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n268), .B(new_n207), .C1(new_n231), .C2(new_n233), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n255), .A2(new_n257), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n221), .A2(G146), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n219), .B2(G143), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n221), .A2(KEYINPUT64), .A3(G146), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n262), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n262), .C1(new_n276), .C2(new_n264), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n278), .A2(KEYINPUT10), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n266), .A2(new_n267), .B1(new_n271), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n240), .A2(new_n252), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n252), .B1(new_n240), .B2(new_n282), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n198), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n277), .B1(new_n258), .B2(new_n259), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n265), .A2(new_n263), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n269), .A2(new_n270), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n251), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT12), .B1(new_n251), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI221_X1 g107(.A(new_n251), .B1(new_n291), .B2(KEYINPUT12), .C1(new_n287), .C2(new_n289), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n198), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n283), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n286), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n194), .B1(new_n298), .B2(new_n193), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n283), .A2(new_n295), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n283), .A2(new_n295), .A3(KEYINPUT82), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n198), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n283), .A2(new_n296), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n283), .A2(KEYINPUT83), .A3(new_n296), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n240), .A2(new_n282), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n251), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n311), .A3(G469), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n192), .B1(new_n299), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G210), .B1(G237), .B2(G902), .ZN(new_n314));
  MUX2_X1   g128(.A(new_n277), .B(new_n230), .S(G125), .Z(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT85), .B(G224), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n316), .A2(G953), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n315), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT2), .B(G113), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G116), .B(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(G116), .B(G119), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n319), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT65), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT65), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(new_n218), .C1(new_n238), .C2(new_n239), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  INV_X1    g145(.A(G116), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G119), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n333), .B2(new_n329), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n322), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n271), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G122), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n328), .A2(new_n338), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n339), .A2(KEYINPUT84), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n340), .A2(KEYINPUT6), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  INV_X1    g158(.A(new_n342), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n344), .B(new_n345), .C1(new_n328), .C2(new_n338), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n318), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT86), .B(new_n318), .C1(new_n343), .C2(new_n346), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n336), .B1(new_n269), .B2(new_n270), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n339), .B(KEYINPUT8), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n317), .A2(KEYINPUT7), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n315), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT87), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n340), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n191), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n314), .B1(new_n351), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n314), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n367), .B(new_n364), .C1(new_n349), .C2(new_n350), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n187), .B(new_n313), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(G113), .B(G122), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(new_n202), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n196), .A3(G214), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n221), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT18), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(new_n249), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(KEYINPUT18), .A3(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n219), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n383));
  INV_X1    g197(.A(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G125), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(KEYINPUT16), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(G146), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n375), .B(G131), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(KEYINPUT17), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n375), .A2(KEYINPUT17), .A3(G131), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT88), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n372), .B(new_n382), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT88), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n390), .B(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(new_n387), .C1(KEYINPUT17), .C2(new_n388), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n397), .A2(KEYINPUT89), .A3(new_n372), .A4(new_n382), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n397), .A2(new_n382), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n372), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n191), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G475), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n386), .A2(new_n219), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n380), .B(KEYINPUT19), .Z(new_n405));
  OAI211_X1 g219(.A(new_n388), .B(new_n404), .C1(G146), .C2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n406), .A2(new_n382), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(new_n372), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n394), .B2(new_n398), .ZN(new_n409));
  NOR2_X1   g223(.A1(G475), .A2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n409), .A2(KEYINPUT20), .A3(new_n411), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(KEYINPUT90), .ZN(new_n414));
  INV_X1    g228(.A(new_n408), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n399), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n410), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT90), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n403), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(G234), .A2(G237), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(G952), .A3(new_n196), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT96), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(G902), .A3(G953), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(G898), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G478), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT15), .ZN(new_n433));
  INV_X1    g247(.A(G122), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G116), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT95), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT91), .B(G122), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n332), .A2(new_n439), .B1(new_n436), .B2(KEYINPUT14), .ZN(new_n440));
  OAI21_X1  g254(.A(G107), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n260), .A2(G143), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT93), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n221), .A2(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G134), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n242), .A3(new_n444), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n436), .B1(new_n439), .B2(new_n332), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n441), .B(new_n448), .C1(G107), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT13), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n443), .B1(KEYINPUT92), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(KEYINPUT92), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n451), .B2(new_n444), .ZN(new_n455));
  OAI21_X1  g269(.A(G134), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n449), .B(G107), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n447), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n458), .A2(KEYINPUT94), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(KEYINPUT94), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n450), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n190), .A2(G217), .A3(new_n196), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n450), .B(new_n464), .C1(new_n459), .C2(new_n460), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n433), .B1(new_n467), .B2(G902), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n466), .B(new_n191), .C1(KEYINPUT15), .C2(new_n432), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n422), .A2(new_n431), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n370), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n230), .A2(new_n251), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n325), .A2(new_n326), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n242), .A2(G137), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n244), .A2(G134), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n250), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n278), .A2(new_n280), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n230), .A2(new_n251), .A3(KEYINPUT66), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n476), .A2(new_n477), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n476), .A2(new_n482), .A3(KEYINPUT30), .A4(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n277), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n474), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n230), .A2(new_n251), .A3(KEYINPUT66), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT66), .B1(new_n230), .B2(new_n251), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n487), .A3(KEYINPUT30), .A4(new_n482), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n485), .B1(new_n497), .B2(new_n327), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n373), .A2(new_n196), .A3(G210), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n499), .B(KEYINPUT27), .Z(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT31), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n477), .B1(new_n492), .B2(new_n496), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT31), .ZN(new_n506));
  NOR4_X1   g320(.A1(new_n505), .A2(new_n506), .A3(new_n502), .A4(new_n485), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n482), .A2(new_n474), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n327), .B1(new_n510), .B2(KEYINPUT69), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n482), .A2(new_n512), .A3(new_n474), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n327), .A2(new_n489), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n515), .B1(new_n484), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n509), .B1(new_n518), .B2(new_n503), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT70), .B(new_n502), .C1(new_n514), .C2(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n473), .B1(new_n508), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n497), .A2(new_n327), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n503), .A3(new_n484), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n506), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n498), .A2(KEYINPUT31), .A3(new_n503), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n484), .A2(new_n516), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT28), .ZN(new_n529));
  INV_X1    g343(.A(new_n513), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n512), .B1(new_n482), .B2(new_n474), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n530), .A2(new_n531), .A3(new_n327), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n532), .B2(KEYINPUT28), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT70), .B1(new_n533), .B2(new_n502), .ZN(new_n534));
  INV_X1    g348(.A(new_n520), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n527), .A2(new_n536), .A3(KEYINPUT71), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n522), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n522), .A2(new_n537), .A3(KEYINPUT72), .A4(new_n538), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n522), .A2(new_n537), .A3(KEYINPUT32), .A4(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(new_n498), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n502), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT29), .B1(new_n518), .B2(new_n503), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n477), .B1(new_n495), .B2(new_n482), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n485), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n514), .B1(new_n552), .B2(KEYINPUT28), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n503), .A2(KEYINPUT29), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G472), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n545), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n544), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n386), .B(new_n219), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n561));
  INV_X1    g375(.A(G119), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n563), .B(new_n564), .C1(G119), .C2(new_n260), .ZN(new_n565));
  XNOR2_X1  g379(.A(G119), .B(G128), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT24), .B(G110), .Z(new_n567));
  AOI22_X1  g381(.A1(new_n565), .A2(G110), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n380), .A2(new_n219), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n565), .A2(G110), .B1(new_n566), .B2(new_n567), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n404), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  INV_X1    g388(.A(G234), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n188), .A2(new_n575), .A3(G953), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n574), .B(new_n576), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n572), .A3(new_n577), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n579), .A2(new_n191), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  OR3_X1    g396(.A1(new_n581), .A2(KEYINPUT74), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n582), .B1(new_n581), .B2(KEYINPUT74), .ZN(new_n584));
  OAI21_X1  g398(.A(G217), .B1(new_n575), .B2(G902), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT73), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n579), .A2(new_n580), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n586), .A2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n559), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n592), .B1(new_n544), .B2(new_n558), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n472), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n235), .ZN(G3));
  OAI211_X1 g414(.A(new_n187), .B(new_n431), .C1(new_n366), .C2(new_n368), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n432), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n463), .A2(new_n603), .A3(new_n465), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n463), .B2(new_n465), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n467), .A2(G902), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT98), .B(G478), .Z(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n421), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n522), .A2(new_n537), .A3(new_n191), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n541), .A2(new_n614), .A3(new_n543), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n313), .A2(new_n593), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n541), .A2(new_n543), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n192), .B(new_n592), .C1(new_n299), .C2(new_n312), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(KEYINPUT97), .A3(new_n614), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n601), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n418), .A2(new_n412), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n403), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n470), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g442(.A1(new_n617), .A2(new_n620), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT35), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n578), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n573), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n590), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n587), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n615), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n370), .A2(new_n471), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  AOI21_X1  g454(.A(new_n636), .B1(new_n544), .B2(new_n558), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n425), .B1(G900), .B2(new_n426), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT100), .Z(new_n643));
  NOR3_X1   g457(.A1(new_n470), .A2(new_n627), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n370), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT101), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n370), .A2(new_n641), .A3(new_n647), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT102), .B(G128), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G30));
  XOR2_X1   g465(.A(new_n643), .B(KEYINPUT39), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n313), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(KEYINPUT40), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(KEYINPUT40), .ZN(new_n655));
  INV_X1    g469(.A(new_n187), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n422), .A2(new_n470), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n654), .A2(new_n655), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n498), .A2(new_n502), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n191), .B1(new_n552), .B2(new_n503), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n545), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n635), .B1(new_n544), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n345), .B1(new_n328), .B2(new_n338), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT6), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n340), .A2(KEYINPUT6), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n665), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT86), .B1(new_n668), .B2(new_n318), .ZN(new_n669));
  INV_X1    g483(.A(new_n350), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n365), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n367), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n351), .A2(new_n314), .A3(new_n365), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT38), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n659), .A2(new_n664), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT103), .B(G143), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G45));
  NOR2_X1   g494(.A1(new_n610), .A2(new_n643), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n370), .A2(new_n641), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT104), .B(G146), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G48));
  INV_X1    g498(.A(new_n610), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n298), .A2(new_n193), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n296), .B1(new_n310), .B2(new_n283), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n283), .A2(new_n295), .A3(new_n296), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n193), .B(new_n191), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n192), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n625), .A2(new_n596), .A3(new_n685), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n625), .A2(new_n596), .A3(new_n628), .A4(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AOI21_X1  g510(.A(new_n656), .B1(new_n672), .B2(new_n673), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n691), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n471), .A3(new_n641), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  XNOR2_X1  g514(.A(new_n538), .B(KEYINPUT105), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n553), .A2(new_n503), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n701), .B1(new_n508), .B2(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n614), .A2(new_n593), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n690), .A2(new_n192), .A3(new_n430), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n697), .A2(new_n704), .A3(new_n657), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  AND3_X1   g521(.A1(new_n614), .A2(new_n635), .A3(new_n703), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n708), .A3(new_n681), .A4(new_n691), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  INV_X1    g524(.A(new_n681), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n672), .A2(new_n187), .A3(new_n673), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n304), .A2(new_n311), .A3(G469), .ZN(new_n714));
  INV_X1    g528(.A(new_n194), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n689), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n299), .A2(KEYINPUT106), .A3(new_n312), .ZN(new_n718));
  INV_X1    g532(.A(new_n192), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n711), .A2(new_n712), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n539), .A2(new_n542), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n592), .B1(new_n558), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(KEYINPUT42), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n712), .A2(new_n720), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n596), .A4(new_n681), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n721), .B2(new_n596), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(G131), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G33));
  NAND3_X1  g547(.A1(new_n725), .A2(new_n596), .A3(new_n644), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT109), .B(G134), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G36));
  NAND2_X1  g550(.A1(new_n304), .A2(new_n311), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n193), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n715), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n744), .A2(new_n745), .B1(new_n193), .B2(new_n298), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n742), .A2(new_n743), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n715), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n192), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n413), .A2(KEYINPUT90), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n418), .A2(new_n419), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n412), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n403), .A3(new_n609), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT43), .B1(new_n753), .B2(KEYINPUT111), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n421), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(KEYINPUT112), .A3(new_n403), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n609), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n759), .B1(new_n753), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n754), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n615), .A3(new_n635), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n366), .A2(new_n368), .A3(new_n656), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n615), .A4(new_n635), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n749), .A2(new_n768), .A3(new_n652), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  NOR4_X1   g584(.A1(new_n559), .A2(new_n711), .A3(new_n712), .A4(new_n593), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n746), .A2(new_n748), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n719), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n384), .ZN(G42));
  NAND3_X1  g593(.A1(new_n544), .A2(new_n593), .A3(new_n663), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n758), .A2(new_n656), .A3(new_n192), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n690), .B(KEYINPUT49), .Z(new_n783));
  NAND4_X1  g597(.A1(new_n676), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n686), .A2(new_n192), .A3(new_n689), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n776), .A2(new_n777), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n425), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n762), .A2(new_n787), .A3(new_n704), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n766), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT118), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n766), .A2(new_n691), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT119), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n425), .B1(new_n792), .B2(KEYINPUT119), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n793), .A2(new_n794), .A3(new_n781), .ZN(new_n795));
  INV_X1    g609(.A(new_n609), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n422), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n793), .A2(new_n794), .A3(new_n708), .A4(new_n762), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n676), .A2(new_n656), .A3(new_n691), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(KEYINPUT50), .A3(new_n788), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT50), .B1(new_n799), .B2(new_n788), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n797), .B(new_n798), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT120), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n802), .B1(new_n786), .B2(new_n790), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT51), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n793), .A2(new_n794), .A3(new_n723), .A4(new_n762), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT48), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n795), .A2(new_n685), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n196), .A2(G952), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n788), .B2(new_n698), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n808), .B1(new_n807), .B2(KEYINPUT117), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n717), .A2(new_n719), .A3(new_n718), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n766), .A2(new_n822), .A3(new_n681), .A4(new_n708), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n636), .A2(new_n627), .A3(new_n643), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n468), .A2(KEYINPUT113), .A3(new_n469), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT113), .B1(new_n468), .B2(new_n469), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n313), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n559), .A2(new_n766), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n559), .A2(new_n593), .A3(new_n644), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n766), .A2(new_n822), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n823), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n734), .A2(KEYINPUT114), .A3(new_n823), .A4(new_n829), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n621), .A2(new_n692), .A3(new_n638), .A4(new_n706), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n599), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n827), .A2(new_n421), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n601), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n617), .A3(new_n620), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n699), .A2(new_n695), .A3(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n731), .A2(new_n836), .A3(new_n838), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n682), .A2(new_n709), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n697), .A2(new_n657), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n720), .A2(new_n643), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n664), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n649), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n845), .B1(new_n648), .B2(new_n646), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n849), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n843), .A2(new_n844), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n844), .B1(new_n843), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n821), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n853), .B2(new_n849), .ZN(new_n860));
  AND4_X1   g674(.A1(KEYINPUT52), .A2(new_n649), .A3(new_n846), .A4(new_n849), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT115), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n836), .A2(new_n838), .A3(new_n731), .A4(new_n842), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n862), .B(new_n844), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n843), .B(new_n855), .C1(KEYINPUT115), .C2(KEYINPUT53), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n821), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT54), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n820), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n784), .B1(new_n872), .B2(new_n873), .ZN(G75));
  OAI21_X1  g688(.A(KEYINPUT53), .B1(new_n863), .B2(new_n864), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n843), .A2(new_n844), .A3(new_n855), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n191), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(G210), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT121), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n668), .B(new_n318), .Z(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n880), .A2(new_n882), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n885), .A2(new_n879), .A3(new_n883), .A4(new_n882), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n196), .A2(G952), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(G51));
  NAND3_X1  g702(.A1(new_n875), .A2(KEYINPUT54), .A3(new_n876), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n858), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n194), .B(KEYINPUT57), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n890), .A2(new_n891), .B1(new_n286), .B2(new_n297), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT122), .ZN(new_n893));
  INV_X1    g707(.A(new_n747), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n892), .A2(KEYINPUT122), .B1(new_n894), .B2(new_n878), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n887), .B1(new_n893), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  OR3_X1    g711(.A1(new_n897), .A2(KEYINPUT123), .A3(new_n409), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT123), .B1(new_n897), .B2(new_n409), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n887), .B1(new_n897), .B2(new_n409), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G60));
  OR2_X1    g715(.A1(new_n604), .A2(new_n605), .ZN(new_n902));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT59), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n890), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n887), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n871), .B(new_n904), .C1(new_n859), .C2(new_n867), .ZN(new_n908));
  INV_X1    g722(.A(new_n902), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(KEYINPUT124), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n877), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n633), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n589), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n906), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n316), .B2(new_n428), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n838), .A2(new_n842), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n928), .B2(G953), .ZN(new_n929));
  INV_X1    g743(.A(new_n668), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(G898), .B2(new_n196), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G69));
  XOR2_X1   g746(.A(new_n497), .B(new_n405), .Z(new_n933));
  INV_X1    g747(.A(new_n853), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n678), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  INV_X1    g750(.A(new_n778), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n595), .A2(new_n598), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n653), .B1(new_n839), .B2(new_n610), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n766), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n936), .A2(new_n769), .A3(new_n937), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n933), .B1(new_n941), .B2(new_n196), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n749), .A2(new_n652), .A3(new_n847), .A4(new_n723), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n731), .A3(new_n734), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n778), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n769), .A2(new_n947), .A3(new_n853), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n769), .B2(new_n853), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n778), .A2(new_n945), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(KEYINPUT127), .C1(new_n949), .C2(new_n948), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n196), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n933), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n942), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n196), .B1(G227), .B2(G900), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  AOI221_X4 g776(.A(new_n942), .B1(new_n958), .B2(new_n962), .C1(new_n954), .C2(new_n956), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(G72));
  NAND3_X1  g778(.A1(new_n951), .A2(new_n928), .A3(new_n953), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  AOI211_X1 g781(.A(new_n503), .B(new_n546), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n941), .B2(new_n927), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n660), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n547), .A2(new_n524), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n869), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n968), .A2(new_n970), .A3(new_n887), .A4(new_n972), .ZN(G57));
endmodule


