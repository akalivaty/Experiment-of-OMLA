//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT79), .B(G197gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(G204gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G197gat), .ZN(new_n212));
  INV_X1    g011(.A(G197gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(KEYINPUT79), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g014(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT29), .B1(new_n216), .B2(KEYINPUT89), .ZN(new_n217));
  INV_X1    g016(.A(new_n206), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n208), .A2(G204gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(KEYINPUT79), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(G197gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n220), .A2(new_n221), .A3(G204gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n207), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n215), .ZN(new_n225));
  INV_X1    g024(.A(new_n207), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n218), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n217), .B1(new_n228), .B2(KEYINPUT89), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g033(.A1(G141gat), .A2(G148gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G155gat), .ZN(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(KEYINPUT81), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G162gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n234), .B1(new_n246), .B2(G155gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n238), .A3(new_n240), .A4(new_n235), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(G162gat), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT2), .B1(new_n251), .B2(new_n239), .ZN(new_n252));
  AND4_X1   g051(.A1(new_n238), .A2(new_n233), .A3(new_n240), .A4(new_n235), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT82), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n242), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT84), .B(new_n242), .C1(new_n250), .C2(new_n254), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n229), .A2(new_n230), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n248), .B1(new_n247), .B2(new_n249), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT82), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n260), .A2(new_n261), .B1(new_n241), .B2(new_n236), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n230), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n228), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n205), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT3), .B1(new_n228), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n204), .B1(new_n267), .B2(new_n262), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n268), .A2(KEYINPUT90), .A3(new_n265), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n226), .B1(new_n225), .B2(new_n218), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n264), .B1(new_n271), .B2(new_n216), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n230), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n205), .B1(new_n273), .B2(new_n255), .ZN(new_n274));
  INV_X1    g073(.A(new_n228), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT29), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n266), .B1(new_n269), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(G22gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(G78gat), .B(G106gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(G50gat), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT90), .B1(new_n268), .B2(new_n265), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n274), .A2(new_n270), .A3(new_n277), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G22gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n288), .B(new_n266), .C1(KEYINPUT91), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n279), .A2(new_n289), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(G22gat), .A3(new_n266), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n285), .B(KEYINPUT88), .Z(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G134gat), .ZN(new_n303));
  INV_X1    g102(.A(G134gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G127gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT72), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G113gat), .A2(G120gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n301), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n299), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n310), .A4(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n262), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT83), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n298), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n257), .A2(new_n315), .A3(new_n258), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT4), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n318), .B1(new_n323), .B2(new_n263), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n262), .A2(new_n315), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT85), .B1(new_n326), .B2(KEYINPUT4), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n320), .B2(KEYINPUT4), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n319), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n263), .ZN(new_n330));
  INV_X1    g129(.A(new_n318), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n298), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n257), .A2(new_n334), .A3(new_n315), .A4(new_n258), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT86), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(KEYINPUT4), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n335), .B2(KEYINPUT86), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n333), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT0), .ZN(new_n343));
  XNOR2_X1  g142(.A(G57gat), .B(G85gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT95), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n341), .A2(new_n349), .A3(KEYINPUT6), .A4(new_n346), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n340), .A3(new_n345), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT6), .B1(new_n341), .B2(new_n346), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n348), .A2(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G226gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(new_n203), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT64), .B(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(G169gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  OAI22_X1  g161(.A1(new_n357), .A2(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(G183gat), .B2(G190gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n356), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(KEYINPUT65), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(G183gat), .A3(G190gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n372), .A3(new_n366), .ZN(new_n373));
  INV_X1    g172(.A(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT66), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G190gat), .ZN(new_n377));
  INV_X1    g176(.A(G183gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n364), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n362), .B1(KEYINPUT23), .B2(new_n360), .ZN(new_n381));
  INV_X1    g180(.A(G176gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n358), .A2(new_n382), .A3(KEYINPUT23), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT25), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT67), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n380), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n380), .B2(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n369), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n362), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT70), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n360), .A2(new_n390), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n358), .A2(new_n382), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n391), .A2(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT70), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n395), .A2(new_n397), .B1(G183gat), .B2(G190gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT66), .B(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT27), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(G183gat), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n400), .B2(G183gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n378), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n399), .A2(new_n401), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n399), .A2(KEYINPUT28), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n378), .A2(KEYINPUT27), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n401), .A2(new_n409), .A3(KEYINPUT69), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT69), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n378), .A2(KEYINPUT27), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n400), .A2(G183gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n398), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT29), .B(new_n355), .C1(new_n389), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT71), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(new_n408), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n419), .A2(new_n420), .B1(new_n405), .B2(new_n406), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n393), .A2(new_n394), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(KEYINPUT70), .B2(new_n396), .ZN(new_n423));
  INV_X1    g222(.A(new_n397), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n367), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n418), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT71), .B(new_n398), .C1(new_n407), .C2(new_n415), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n389), .A2(new_n426), .A3(new_n427), .A4(new_n355), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n228), .B1(new_n417), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n389), .A2(new_n426), .A3(new_n427), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n355), .A2(KEYINPUT29), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n389), .A2(new_n416), .A3(new_n355), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n275), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n431), .B1(new_n430), .B2(new_n436), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT38), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n430), .A2(new_n440), .A3(new_n436), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n275), .B1(new_n417), .B2(new_n429), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n434), .A2(new_n228), .A3(new_n435), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n440), .B(KEYINPUT80), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT38), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n437), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n444), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n297), .B1(new_n353), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n454));
  INV_X1    g253(.A(new_n449), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n434), .A2(new_n275), .A3(new_n435), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n389), .A2(new_n416), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n433), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n275), .B1(new_n458), .B2(new_n428), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n455), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n454), .B1(new_n460), .B2(new_n445), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n445), .A2(new_n454), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT93), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n456), .A2(new_n441), .A3(new_n459), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n449), .B1(new_n430), .B2(new_n436), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT30), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n445), .A2(new_n454), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n257), .A2(new_n258), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n334), .A4(new_n315), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n336), .A3(new_n338), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n331), .B1(new_n474), .B2(new_n330), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT39), .B1(new_n316), .B2(new_n318), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT94), .B(KEYINPUT39), .Z(new_n478));
  AOI21_X1  g277(.A(new_n346), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n341), .A2(new_n346), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT40), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n470), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n468), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n487), .A3(new_n351), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n488), .B2(new_n347), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n291), .A2(new_n491), .A3(new_n295), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n291), .B2(new_n295), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n453), .A2(new_n485), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n432), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT73), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n312), .A2(new_n314), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(new_n389), .A3(new_n426), .A4(new_n427), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT74), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n507));
  AOI211_X1 g306(.A(new_n507), .B(new_n504), .C1(new_n498), .C2(new_n502), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT32), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT33), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n506), .B2(new_n508), .ZN(new_n511));
  XOR2_X1   g310(.A(G15gat), .B(G43gat), .Z(new_n512));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n514), .ZN(new_n516));
  OAI221_X1 g315(.A(KEYINPUT32), .B1(new_n510), .B2(new_n516), .C1(new_n506), .C2(new_n508), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT34), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n518), .A3(new_n504), .A4(new_n502), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT34), .B1(new_n503), .B2(new_n505), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n520), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n515), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n515), .B2(new_n517), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n496), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT78), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT78), .B(new_n496), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n517), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n525), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g333(.A(KEYINPUT76), .B(new_n524), .C1(new_n515), .C2(new_n517), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT36), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n489), .B(new_n296), .C1(new_n534), .C2(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n297), .A2(KEYINPUT35), .ZN(new_n540));
  INV_X1    g339(.A(new_n353), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n527), .ZN(new_n542));
  INV_X1    g341(.A(new_n470), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n495), .A2(new_n537), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT98), .B(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G29gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(G29gat), .A2(G36gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT14), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(KEYINPUT14), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G43gat), .B(G50gat), .Z(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT99), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n551), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n554), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n558));
  INV_X1    g357(.A(new_n556), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n558), .B(new_n559), .C1(KEYINPUT99), .C2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT100), .ZN(new_n563));
  INV_X1    g362(.A(G1gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n562), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(KEYINPUT16), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G8gat), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n565), .B2(new_n569), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n557), .B(new_n561), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n561), .A2(new_n557), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n565), .A2(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G8gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n561), .B2(new_n557), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n573), .B(new_n574), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT97), .ZN(new_n589));
  XOR2_X1   g388(.A(G169gat), .B(G197gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT96), .B(KEYINPUT11), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT12), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n591), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n557), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n578), .A2(new_n600), .A3(new_n579), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n573), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n574), .B(KEYINPUT13), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(KEYINPUT17), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(new_n578), .A3(new_n579), .A4(new_n576), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n606), .A2(KEYINPUT18), .A3(new_n574), .A4(new_n573), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n582), .A2(new_n584), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(new_n604), .A3(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(new_n599), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n587), .A2(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n545), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G57gat), .B(G64gat), .Z(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  INV_X1    g415(.A(G71gat), .ZN(new_n617));
  INV_X1    g416(.A(G78gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G78gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n615), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT102), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n623), .A2(new_n615), .A3(KEYINPUT102), .A4(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n302), .ZN(new_n631));
  AOI211_X1 g430(.A(new_n572), .B(new_n571), .C1(KEYINPUT21), .C2(new_n627), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n239), .ZN(new_n635));
  XOR2_X1   g434(.A(G183gat), .B(G211gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n633), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G85gat), .A2(G92gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT7), .ZN(new_n640));
  XNOR2_X1  g439(.A(G99gat), .B(G106gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(G99gat), .A2(G106gat), .ZN(new_n642));
  INV_X1    g441(.A(G85gat), .ZN(new_n643));
  INV_X1    g442(.A(G92gat), .ZN(new_n644));
  AOI22_X1  g443(.A1(KEYINPUT8), .A2(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n641), .B1(new_n640), .B2(new_n645), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n605), .A2(new_n576), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n655));
  NAND2_X1  g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656));
  OAI22_X1  g455(.A1(new_n600), .A2(new_n649), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G190gat), .B(G218gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT105), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n656), .A2(new_n655), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT103), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n663), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n660), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n654), .A2(new_n658), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n661), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n666), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n667), .B1(new_n654), .B2(new_n658), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n657), .B(new_n660), .C1(new_n652), .C2(new_n653), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n638), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(G230gat), .A2(G233gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n627), .A2(new_n648), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n625), .B(new_n626), .C1(new_n646), .C2(new_n647), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n649), .A2(KEYINPUT106), .A3(new_n626), .A4(new_n625), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT10), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n648), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n680), .A2(G230gat), .A3(G233gat), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G120gat), .B(G148gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(G176gat), .B(G204gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n675), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n614), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n488), .A2(new_n347), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(new_n564), .ZN(G1324gat));
  NOR2_X1   g497(.A1(new_n695), .A2(new_n543), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT108), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n695), .B2(new_n543), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(G8gat), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT16), .B(G8gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT109), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n699), .A2(KEYINPUT42), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n700), .B2(new_n702), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n703), .B(new_n707), .C1(new_n708), .C2(new_n709), .ZN(G1325gat));
  INV_X1    g509(.A(G15gat), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n695), .A2(new_n711), .A3(new_n537), .ZN(new_n712));
  INV_X1    g511(.A(new_n542), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n695), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(G1326gat));
  INV_X1    g517(.A(new_n494), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n695), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT43), .B(G22gat), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  INV_X1    g521(.A(new_n638), .ZN(new_n723));
  INV_X1    g522(.A(new_n693), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n674), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT111), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n614), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(G29gat), .A3(new_n696), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT45), .Z(new_n730));
  NAND2_X1  g529(.A1(new_n495), .A2(new_n537), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n539), .A2(new_n544), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n674), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(KEYINPUT44), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n545), .B2(new_n674), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n725), .A2(new_n613), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n740), .B2(new_n696), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n730), .A2(new_n741), .ZN(G1328gat));
  OAI21_X1  g541(.A(new_n546), .B1(new_n740), .B2(new_n543), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n728), .A2(new_n543), .A3(new_n546), .ZN(new_n744));
  NAND2_X1  g543(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT112), .B(KEYINPUT46), .Z(new_n747));
  OAI211_X1 g546(.A(new_n743), .B(new_n746), .C1(new_n744), .C2(new_n747), .ZN(G1329gat));
  INV_X1    g547(.A(new_n537), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n738), .A2(new_n749), .A3(new_n739), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n611), .A2(new_n612), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n610), .A2(KEYINPUT101), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n755), .B2(new_n608), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n713), .A2(G43gat), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n727), .A2(new_n733), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n758), .B(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(G43gat), .B2(new_n750), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n763));
  OAI21_X1  g562(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(G1330gat));
  NAND3_X1  g563(.A1(new_n738), .A2(new_n297), .A3(new_n739), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G50gat), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n728), .A2(G50gat), .A3(new_n719), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(KEYINPUT48), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n735), .A2(new_n737), .A3(new_n494), .A4(new_n739), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n770), .A2(new_n771), .A3(G50gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(G50gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n772), .A2(new_n773), .A3(new_n767), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n769), .B1(new_n774), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g574(.A1(new_n675), .A2(new_n756), .A3(new_n724), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n733), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n733), .A2(KEYINPUT116), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n696), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(G57gat), .Z(G1332gat));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n470), .A3(new_n780), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  OAI21_X1  g586(.A(G71gat), .B1(new_n781), .B2(new_n537), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n779), .A2(new_n617), .A3(new_n542), .A4(new_n780), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(KEYINPUT50), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1334gat));
  NOR2_X1   g593(.A1(new_n781), .A2(new_n719), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n618), .ZN(G1335gat));
  NOR2_X1   g595(.A1(new_n545), .A2(new_n674), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n638), .A2(new_n756), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n797), .A2(KEYINPUT51), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n696), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n801), .A2(new_n643), .A3(new_n802), .A4(new_n693), .ZN(new_n803));
  INV_X1    g602(.A(new_n798), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n724), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n738), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n696), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(G1336gat));
  NOR3_X1   g607(.A1(new_n543), .A2(G92gat), .A3(new_n724), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n799), .B2(new_n800), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n735), .A2(new_n737), .A3(new_n470), .A4(new_n805), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G92gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g613(.A1(new_n713), .A2(G99gat), .A3(new_n724), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G99gat), .B1(new_n806), .B2(new_n537), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1338gat));
  NOR3_X1   g617(.A1(new_n296), .A2(G106gat), .A3(new_n724), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n799), .B2(new_n800), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n735), .A2(new_n737), .A3(new_n297), .A4(new_n805), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n738), .A2(new_n494), .A3(new_n805), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n801), .A2(new_n819), .B1(new_n825), .B2(G106gat), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G1339gat));
  OR3_X1    g627(.A1(new_n682), .A2(new_n676), .A3(new_n683), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(KEYINPUT54), .A3(new_n684), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n676), .C1(new_n682), .C2(new_n683), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n690), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT55), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n756), .A2(new_n836), .A3(new_n692), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n574), .B1(new_n606), .B2(new_n573), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n602), .A2(new_n603), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n593), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT118), .B(new_n593), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n587), .A2(new_n609), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n693), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n838), .A2(KEYINPUT119), .A3(new_n847), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n674), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n845), .A2(new_n846), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n692), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n734), .A2(new_n836), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n723), .ZN(new_n858));
  AND4_X1   g657(.A1(new_n613), .A2(new_n638), .A3(new_n674), .A4(new_n724), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n696), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n534), .A2(new_n535), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n296), .A4(new_n543), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n756), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n713), .B(new_n494), .C1(new_n858), .C2(new_n860), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n470), .A2(new_n696), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n307), .A3(new_n613), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n865), .A2(new_n869), .ZN(G1340gat));
  AOI21_X1  g669(.A(G120gat), .B1(new_n864), .B2(new_n693), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n868), .A2(new_n308), .A3(new_n724), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(G1341gat));
  NAND3_X1  g672(.A1(new_n864), .A2(new_n302), .A3(new_n638), .ZN(new_n874));
  OAI21_X1  g673(.A(G127gat), .B1(new_n868), .B2(new_n723), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1342gat));
  NAND3_X1  g675(.A1(new_n864), .A2(new_n304), .A3(new_n734), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n868), .B2(new_n674), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  NOR3_X1   g680(.A1(new_n749), .A2(new_n296), .A3(new_n470), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n861), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n231), .B1(new_n883), .B2(new_n613), .ZN(new_n884));
  OR2_X1    g683(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n638), .B1(new_n852), .B2(new_n856), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n886), .B(new_n297), .C1(new_n887), .C2(new_n859), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT120), .B1(new_n834), .B2(new_n835), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n890), .B(KEYINPUT55), .C1(new_n830), .C2(new_n833), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n613), .A2(new_n854), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n892), .A2(new_n893), .B1(new_n853), .B2(new_n693), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n856), .B1(new_n894), .B2(new_n734), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n859), .B1(new_n895), .B2(new_n723), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n896), .B2(new_n719), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n537), .A2(new_n867), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n888), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n756), .A2(G141gat), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n884), .B(new_n885), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n901), .B(new_n902), .ZN(G1344gat));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n897), .A3(new_n693), .A4(new_n898), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n232), .A2(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT122), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n895), .A2(new_n723), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n886), .B(new_n494), .C1(new_n911), .C2(new_n859), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n898), .A2(new_n693), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n296), .B1(new_n858), .B2(new_n860), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n912), .B(new_n913), .C1(new_n914), .C2(new_n886), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G148gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT123), .B1(new_n916), .B2(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n918), .B(new_n919), .C1(new_n915), .C2(G148gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n910), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n883), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n232), .A3(new_n693), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1345gat));
  NOR3_X1   g723(.A1(new_n899), .A2(new_n239), .A3(new_n723), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n883), .A2(KEYINPUT124), .A3(new_n723), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(G155gat), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT124), .B1(new_n883), .B2(new_n723), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(new_n246), .B1(new_n899), .B2(new_n674), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n734), .A2(new_n251), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n883), .B2(new_n931), .ZN(G1347gat));
  AOI21_X1  g731(.A(new_n802), .B1(new_n858), .B2(new_n860), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n862), .A2(new_n296), .A3(new_n470), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n358), .B1(new_n936), .B2(new_n613), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n543), .A2(new_n802), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n866), .A2(G169gat), .A3(new_n756), .A4(new_n938), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(new_n382), .B1(new_n936), .B2(new_n724), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n866), .A2(new_n357), .A3(new_n693), .A4(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT125), .Z(G1349gat));
  NAND3_X1  g743(.A1(new_n866), .A2(new_n638), .A3(new_n938), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G183gat), .ZN(new_n946));
  INV_X1    g745(.A(new_n936), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n419), .A3(new_n638), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n946), .A2(new_n948), .A3(new_n949), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n947), .A2(new_n399), .A3(new_n734), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n866), .A2(new_n734), .A3(new_n938), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G190gat), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n537), .A2(new_n297), .A3(new_n470), .ZN(new_n962));
  OAI221_X1 g761(.A(new_n696), .B1(new_n887), .B2(new_n859), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n756), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n914), .A2(new_n886), .ZN(new_n966));
  INV_X1    g765(.A(new_n912), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n537), .A2(new_n938), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n613), .A2(new_n213), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  NAND3_X1  g770(.A1(new_n964), .A2(new_n210), .A3(new_n693), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n964), .A2(new_n974), .A3(new_n210), .A4(new_n693), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n969), .A2(new_n693), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n973), .B(new_n975), .C1(new_n210), .C2(new_n976), .ZN(G1353gat));
  INV_X1    g776(.A(G211gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n978), .A3(new_n638), .ZN(new_n979));
  INV_X1    g778(.A(new_n966), .ZN(new_n980));
  INV_X1    g779(.A(new_n968), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n980), .A2(new_n638), .A3(new_n912), .A4(new_n981), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  INV_X1    g784(.A(G218gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n964), .A2(new_n986), .A3(new_n734), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n969), .A2(new_n734), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(new_n986), .ZN(G1355gat));
endmodule


