//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g032(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n467), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n470), .B1(new_n463), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(G112), .B2(new_n463), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n474), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n481), .A2(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n463), .A2(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n489), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n474), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n463), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .A3(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n506), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(new_n503), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(G166));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n504), .B2(new_n506), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT71), .B(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n507), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n511), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n524), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n507), .A2(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n532), .B1(new_n512), .B2(new_n533), .C1(new_n534), .C2(new_n503), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  AOI22_X1  g111(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n503), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G81), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n507), .A2(G43), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n520), .A2(G91), .ZN(new_n550));
  OAI21_X1  g125(.A(G65), .B1(new_n517), .B2(new_n518), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT74), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  AND4_X1   g132(.A1(new_n557), .A2(new_n510), .A3(G53), .A4(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n557), .B1(new_n507), .B2(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n549), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n505), .A2(KEYINPUT6), .A3(G651), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT6), .B1(new_n505), .B2(G651), .ZN(new_n563));
  OAI211_X1 g138(.A(G53), .B(G543), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n507), .A2(new_n557), .A3(G53), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OR2_X1    g144(.A1(KEYINPUT5), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(KEYINPUT5), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n552), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n574), .A2(G651), .A3(new_n553), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n567), .A2(new_n575), .A3(KEYINPUT75), .A4(new_n550), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n561), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G299));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n507), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n512), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n519), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n510), .A2(G86), .A3(new_n511), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n507), .A2(G48), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n520), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n507), .A2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n519), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT76), .Z(new_n599));
  AOI21_X1  g174(.A(KEYINPUT10), .B1(new_n520), .B2(G92), .ZN(new_n600));
  AND4_X1   g175(.A1(KEYINPUT10), .A2(new_n510), .A3(G92), .A4(new_n511), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n519), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n602), .A2(KEYINPUT77), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n600), .B2(new_n601), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n599), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n599), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n577), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n577), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n542), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(G559), .B1(new_n607), .B2(new_n610), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n474), .A2(new_n468), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n482), .A2(G135), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT79), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(new_n485), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G123), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n626), .A2(new_n627), .B1(new_n630), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n629), .B(new_n640), .C1(new_n630), .C2(new_n639), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT80), .B(KEYINPUT14), .Z(new_n642));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n644), .B2(new_n645), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n647), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n652), .B2(new_n654), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT81), .Z(new_n660));
  NOR2_X1   g235(.A1(G2072), .A2(G2078), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n444), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(KEYINPUT17), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n658), .B(new_n659), .C1(new_n444), .C2(new_n661), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n660), .A3(new_n658), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT82), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n681), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n676), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n678), .A2(new_n679), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n685), .B(new_n676), .S(new_n686), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n684), .A2(new_n687), .A3(new_n689), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n693), .B1(new_n691), .B2(new_n694), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n674), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(new_n673), .A3(new_n695), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(G229));
  INV_X1    g276(.A(KEYINPUT103), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G33), .ZN(new_n704));
  NAND2_X1  g279(.A1(G115), .A2(G2104), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n465), .ZN(new_n706));
  INV_X1    g281(.A(G127), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n710));
  NAND2_X1  g285(.A1(G103), .A2(G2104), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G2105), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n482), .A2(G139), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n709), .A2(KEYINPUT95), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n704), .B1(new_n719), .B2(G29), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(new_n442), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT96), .Z(new_n722));
  OAI211_X1 g297(.A(G129), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT97), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT97), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n474), .A2(new_n725), .A3(G129), .A4(G2105), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT26), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g307(.A(G141), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n468), .A2(G105), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT98), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n727), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n727), .B2(new_n735), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G29), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT99), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G29), .C2(G32), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n739), .A2(KEYINPUT99), .A3(G29), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G34), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n703), .B1(new_n746), .B2(G34), .ZN(new_n748));
  OAI22_X1  g323(.A1(new_n476), .A2(new_n703), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n720), .B2(new_n442), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n722), .A2(KEYINPUT100), .A3(new_n745), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT101), .B(KEYINPUT31), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G11), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT102), .B(G28), .Z(new_n761));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n703), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n760), .B1(new_n763), .B2(new_n764), .C1(new_n638), .C2(new_n703), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n703), .A2(G27), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n499), .B2(G29), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n443), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n443), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n749), .A2(new_n750), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n758), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n703), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n703), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT29), .B(G2090), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n754), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n754), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G1966), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n778), .A2(G1966), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n772), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n754), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT23), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n577), .B2(new_n754), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n753), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n722), .A2(new_n745), .A3(new_n752), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G116), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n467), .B1(new_n793), .B2(G2105), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT91), .B1(G104), .B2(G2105), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(KEYINPUT91), .A2(G104), .A3(G2105), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(G140), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n799));
  OAI211_X1 g374(.A(G128), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT92), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n703), .A2(G26), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT28), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2067), .ZN(new_n808));
  NOR2_X1   g383(.A1(G4), .A2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n611), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n542), .A2(G16), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n754), .A2(G19), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT89), .B(G1341), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n808), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT94), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n808), .A2(new_n822), .A3(new_n812), .A4(new_n819), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n789), .A2(new_n792), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(G16), .A2(G23), .ZN(new_n825));
  NAND2_X1  g400(.A1(G288), .A2(KEYINPUT87), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n520), .A2(G87), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT87), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n827), .A2(new_n828), .A3(new_n580), .A4(new_n581), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n825), .B1(new_n830), .B2(new_n754), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT33), .B(G1976), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G6), .A2(G16), .ZN(new_n835));
  INV_X1    g410(.A(G305), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(G16), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT32), .B(G1981), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n754), .A2(G22), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G166), .B2(new_n754), .ZN(new_n841));
  INV_X1    g416(.A(G1971), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n831), .A2(new_n833), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n834), .A2(new_n839), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n703), .A2(G25), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G107), .B2(new_n463), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT84), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n482), .A2(G131), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n636), .A2(G119), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n847), .B1(new_n855), .B2(new_n703), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT35), .B(G1991), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT85), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n856), .B(new_n858), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n754), .A2(G24), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT86), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(G290), .B2(G16), .ZN(new_n862));
  INV_X1    g437(.A(G1986), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT88), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n859), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n845), .A2(KEYINPUT34), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n846), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n865), .A3(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n866), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n846), .A2(new_n868), .A3(new_n872), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n702), .B1(new_n824), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n871), .A2(new_n873), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n821), .A2(new_n823), .ZN(new_n877));
  AND4_X1   g452(.A1(new_n792), .A2(new_n753), .A3(new_n788), .A4(new_n783), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT103), .A4(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n875), .A2(new_n879), .ZN(G311));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G150));
  XOR2_X1   g456(.A(KEYINPUT107), .B(G860), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G67), .ZN(new_n884));
  INV_X1    g459(.A(G80), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n519), .A2(new_n884), .B1(new_n885), .B2(new_n501), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  OAI221_X1 g463(.A(new_n888), .B1(new_n885), .B2(new_n501), .C1(new_n519), .C2(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(G651), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n510), .A2(G93), .A3(new_n511), .ZN(new_n892));
  OAI211_X1 g467(.A(G55), .B(G543), .C1(new_n562), .C2(new_n563), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n892), .A2(new_n893), .A3(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT106), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n890), .B(new_n898), .C1(new_n894), .C2(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n543), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n542), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT38), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n608), .B(KEYINPUT77), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n617), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n903), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n883), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n896), .A2(new_n883), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n910), .B(KEYINPUT37), .Z(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(G145));
  AND3_X1   g487(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n499), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n493), .A2(new_n474), .B1(new_n495), .B2(new_n497), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n801), .A2(new_n490), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n738), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n727), .A2(new_n735), .A3(new_n736), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n916), .B(new_n914), .C1(new_n737), .C2(new_n738), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n717), .A2(new_n718), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n727), .A2(new_n735), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n914), .A3(new_n916), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n715), .A3(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n923), .A2(new_n854), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n854), .B1(new_n923), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n625), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n923), .A2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n855), .ZN(new_n933));
  INV_X1    g508(.A(new_n625), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n923), .A2(new_n854), .A3(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n636), .A2(G130), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n482), .A2(G142), .ZN(new_n939));
  OR2_X1    g514(.A1(G106), .A2(G2105), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n940), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n638), .B(G160), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(G162), .Z(new_n945));
  INV_X1    g520(.A(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n931), .A2(new_n936), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n943), .A2(KEYINPUT108), .A3(new_n945), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n943), .A2(new_n947), .ZN(new_n953));
  INV_X1    g528(.A(new_n945), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n952), .A2(KEYINPUT40), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT40), .B1(new_n952), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(G395));
  INV_X1    g533(.A(G290), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n826), .A3(new_n829), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n826), .B2(new_n829), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT111), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n830), .A2(G290), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n960), .ZN(new_n966));
  NAND2_X1  g541(.A1(G303), .A2(new_n836), .ZN(new_n967));
  NAND2_X1  g542(.A1(G166), .A2(G305), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n969), .B(KEYINPUT111), .C1(new_n962), .C2(new_n961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT42), .Z(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n510), .A2(G91), .A3(new_n511), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n573), .B1(new_n511), .B2(G65), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n503), .B1(new_n977), .B2(KEYINPUT74), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n978), .B2(new_n574), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT75), .B1(new_n979), .B2(new_n567), .ZN(new_n980));
  AND4_X1   g555(.A1(KEYINPUT75), .A2(new_n567), .A3(new_n575), .A4(new_n550), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n561), .A2(KEYINPUT109), .A3(new_n576), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n608), .A3(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n577), .A2(new_n975), .A3(new_n602), .A4(new_n606), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n984), .A2(KEYINPUT41), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT41), .B1(new_n984), .B2(new_n985), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n902), .B(new_n621), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(KEYINPUT110), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n984), .A2(KEYINPUT41), .A3(new_n985), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT41), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n608), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n561), .B2(new_n576), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n985), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n989), .A2(new_n991), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n984), .A2(new_n985), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(new_n989), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n990), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT112), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n990), .B(new_n1004), .C1(new_n998), .C2(new_n1001), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n974), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1005), .A2(new_n974), .ZN(new_n1007));
  OAI21_X1  g582(.A(G868), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n896), .A2(new_n619), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(G295));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1009), .ZN(G331));
  XOR2_X1   g586(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n1012));
  NOR2_X1   g587(.A1(G171), .A2(G168), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G301), .A2(G286), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n899), .A2(new_n543), .ZN(new_n1016));
  INV_X1    g591(.A(new_n894), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n892), .A2(new_n893), .A3(new_n891), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n898), .B1(new_n1019), .B2(new_n890), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n901), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n900), .A2(new_n1024), .A3(new_n901), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n997), .A2(new_n991), .A3(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n984), .A2(new_n985), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n900), .A2(new_n1024), .A3(KEYINPUT114), .A4(new_n901), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1028), .A2(new_n1023), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n973), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1027), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1027), .A2(new_n1032), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n991), .A3(new_n997), .ZN(new_n1041));
  AND4_X1   g616(.A1(new_n985), .A2(new_n1023), .A3(new_n984), .A4(new_n1025), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n973), .A2(KEYINPUT115), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n971), .A2(new_n1046), .A3(new_n972), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G37), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1038), .A2(new_n1039), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1052));
  AOI21_X1  g627(.A(G37), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1039), .B1(new_n1038), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1012), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1038), .A2(new_n1039), .A3(new_n1053), .ZN(new_n1056));
  INV_X1    g631(.A(G37), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1042), .B1(new_n988), .B2(new_n1040), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1048), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT44), .B(new_n1056), .C1(new_n1060), .C2(new_n1039), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1061), .ZN(G397));
  INV_X1    g637(.A(G1384), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n499), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT45), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n470), .B(G40), .C1(new_n463), .C2(new_n475), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1996), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT117), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT46), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G2067), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n801), .B(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1068), .B1(new_n1076), .B2(new_n924), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT47), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1068), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n926), .A2(new_n1069), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(new_n1075), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1071), .B2(new_n739), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n858), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT127), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n801), .A2(G2067), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1068), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n854), .B(new_n858), .Z(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1068), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1068), .A2(new_n863), .A3(new_n959), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT48), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1079), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G290), .B(new_n863), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1092), .B1(new_n1080), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1067), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1384), .B1(new_n915), .B2(new_n490), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT45), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1971), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G113), .A2(G2104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n463), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n466), .A2(new_n469), .ZN(new_n1107));
  INV_X1    g682(.A(G40), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT50), .B(G1384), .C1(new_n915), .C2(new_n490), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1111), .A2(new_n1112), .A3(G2090), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(G8), .B1(new_n513), .B2(new_n515), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT55), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G305), .A2(G1981), .ZN(new_n1120));
  INV_X1    g695(.A(G1981), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n587), .A2(new_n1121), .A3(new_n588), .A4(new_n589), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(KEYINPUT49), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1120), .A2(new_n1125), .A3(KEYINPUT49), .A4(new_n1122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT49), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1128));
  INV_X1    g703(.A(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1109), .B2(new_n1101), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1109), .B1(new_n1101), .B2(KEYINPUT45), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1065), .B(G1384), .C1(new_n915), .C2(new_n490), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1064), .A2(KEYINPUT50), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1109), .A3(new_n1138), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1136), .A2(G1971), .B1(new_n1139), .B2(G2090), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(G8), .A3(new_n1117), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n826), .A2(G1976), .A3(new_n829), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1130), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1143), .A2(new_n1130), .ZN(new_n1145));
  INV_X1    g720(.A(G1976), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT52), .B1(G288), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1119), .A2(new_n1133), .A3(new_n1141), .A4(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1066), .A2(new_n1102), .A3(new_n443), .A4(new_n1109), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n757), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1102), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(G171), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1966), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1137), .A2(new_n1138), .A3(new_n750), .A4(new_n1109), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(G168), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G8), .ZN(new_n1162));
  AOI21_X1  g737(.A(G168), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT51), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT51), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1165), .A3(G8), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT62), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1164), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1157), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1129), .B(G286), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1149), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1117), .B1(new_n1140), .B2(G8), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1148), .A2(new_n1133), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1178), .A2(KEYINPUT63), .A3(new_n1179), .A4(new_n1173), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1133), .A2(new_n1182), .B1(new_n1121), .B2(new_n836), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1148), .A2(new_n1133), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1183), .A2(new_n1131), .B1(new_n1184), .B2(new_n1141), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1171), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1149), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(G301), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1156), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT54), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1188), .A2(new_n1192), .A3(new_n1167), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(KEYINPUT124), .A3(G301), .A4(new_n1152), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1191), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1155), .A2(new_n1200), .A3(G171), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n787), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1204));
  XNOR2_X1  g779(.A(KEYINPUT56), .B(G2072), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1066), .A2(new_n1102), .A3(new_n1109), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT57), .B1(new_n556), .B2(new_n560), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT57), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n979), .A2(new_n1208), .A3(new_n567), .ZN(new_n1209));
  AOI22_X1  g784(.A1(new_n1204), .A2(new_n1206), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n1211));
  OAI21_X1  g786(.A(KEYINPUT61), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1209), .A2(new_n1207), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1067), .B1(new_n1064), .B2(KEYINPUT50), .ZN(new_n1214));
  AOI21_X1  g789(.A(G1956), .B1(new_n1214), .B2(new_n1138), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1205), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1134), .A2(new_n1135), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1213), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1212), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(KEYINPUT119), .B(G1996), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1066), .A2(new_n1102), .A3(new_n1109), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1109), .A2(new_n1101), .ZN(new_n1224));
  XOR2_X1   g799(.A(KEYINPUT58), .B(G1341), .Z(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n542), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT120), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT121), .ZN(new_n1229));
  NAND4_X1  g804(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(KEYINPUT59), .ZN(new_n1230));
  OAI21_X1  g805(.A(KEYINPUT59), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1218), .A2(new_n1211), .A3(KEYINPUT61), .A4(new_n1219), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1221), .A2(new_n1230), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n811), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1109), .A2(new_n1101), .A3(new_n1074), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1236), .A2(KEYINPUT60), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1240), .ZN(new_n1241));
  OAI22_X1  g816(.A1(new_n1239), .A2(new_n611), .B1(new_n1241), .B2(KEYINPUT60), .ZN(new_n1242));
  OR2_X1    g817(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n904), .B1(new_n1238), .B2(KEYINPUT123), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g820(.A1(new_n1235), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1218), .B1(new_n904), .B2(new_n1241), .ZN(new_n1247));
  AND2_X1   g822(.A1(new_n1247), .A2(new_n1219), .ZN(new_n1248));
  OAI211_X1 g823(.A(new_n1193), .B(new_n1203), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1249));
  AOI211_X1 g824(.A(KEYINPUT126), .B(new_n1099), .C1(new_n1187), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1251));
  AOI21_X1  g826(.A(new_n1185), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1252));
  INV_X1    g827(.A(new_n1235), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1254));
  OAI221_X1 g829(.A(new_n1254), .B1(KEYINPUT60), .B2(new_n1241), .C1(new_n611), .C2(new_n1239), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1248), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g831(.A1(new_n1203), .A2(new_n1188), .A3(new_n1192), .A4(new_n1167), .ZN(new_n1257));
  OAI211_X1 g832(.A(new_n1171), .B(new_n1252), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  INV_X1    g833(.A(new_n1099), .ZN(new_n1259));
  AOI21_X1  g834(.A(new_n1251), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1097), .B1(new_n1250), .B2(new_n1260), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g836(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1263));
  AND3_X1   g837(.A1(new_n931), .A2(new_n936), .A3(new_n946), .ZN(new_n1264));
  AOI21_X1  g838(.A(new_n946), .B1(new_n931), .B2(new_n936), .ZN(new_n1265));
  NOR2_X1   g839(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g840(.A(KEYINPUT108), .B1(new_n1266), .B2(new_n945), .ZN(new_n1267));
  INV_X1    g841(.A(new_n951), .ZN(new_n1268));
  OAI21_X1  g842(.A(new_n955), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g843(.A(G319), .B(new_n671), .C1(new_n655), .C2(new_n656), .ZN(new_n1270));
  AOI21_X1  g844(.A(new_n1270), .B1(new_n698), .B2(new_n700), .ZN(new_n1271));
  NAND2_X1  g845(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g846(.A1(new_n1263), .A2(new_n1272), .ZN(G308));
  OAI211_X1 g847(.A(new_n1269), .B(new_n1271), .C1(new_n1051), .C2(new_n1054), .ZN(G225));
endmodule


